`define WIDTH  256

//`define FPGA

