// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`ifndef SYNTHESIS
  export "DPI-C" function simutil_get_scramble_key;

  function int simutil_get_scramble_key(output bit [127:0] val);
    int valid;
    valid = key_valid_i && DataKeyWidth == 128 ? 1 : 0;
    if (valid == 1) val = key_i;
    return valid;
  endfunction

  export "DPI-C" function simutil_get_scramble_nonce;

  function int simutil_get_scramble_nonce(output bit [319:0] nonce);
    int valid;
    valid = key_valid_i && NonceWidth <= 320 ? 1 : 0;
    if (valid == 1) begin
       nonce = '0;
       nonce[NonceWidth-1:0] = nonce_i;
    end
    return valid;
  endfunction
`endif


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * Memory loader for simulation
 *
 * Include this file in a memory primitive to load a memory array from
 * simulation.
 *
 * Requirements:
 * - A memory array named `mem`.
 * - A parameter `Width` giving the memory width (word size) in bit.
 * - A parameter `Depth` giving the memory depth in words.
 * - A parameter `MemInitFile` with a file path of a VMEM file to be loaded into
 *   the memory if not empty.
 *
 * Note this works with memories up to a maximum width of 312 bits. Should this maximum width be
 * increased all of the `simutil_set_mem` and `simutil_get_mem` call sites must be found (e.g. using
 * git grep) and adjusted appropriately.
 */

`ifndef SYNTHESIS
  // Task for loading 'mem' with SystemVerilog system task $readmemh()
  export "DPI-C" task simutil_memload;

  task simutil_memload;
    input string file;
    $readmemh(file, mem);
  endtask

  // Function for setting a specific element in |mem|
  // Returns 1 (true) for success, 0 (false) for errors.
  export "DPI-C" function simutil_set_mem;

  function int simutil_set_mem(input int index, input bit [311:0] val);
    int valid;
    valid = Width > 312 || index >= Depth ? 0 : 1;
    if (valid == 1) mem[index] = val[Width-1:0];
    return valid;
  endfunction

  // Function for getting a specific element in |mem|
  export "DPI-C" function simutil_get_mem;

  function int simutil_get_mem(input int index, output bit [311:0] val);
    int valid;
    valid = Width > 312 || index >= Depth ? 0 : 1;
    if (valid == 1) begin
      val = 0;
      val[Width-1:0] = mem[index];
    end
    return valid;
  endfunction
`endif

initial begin
  logic show_mem_paths;

  // Print the hierarchical path to the memory to help make formal connectivity checks easy.
  void'($value$plusargs("show_mem_paths=%0b", show_mem_paths));
  if (show_mem_paths) $display("%m");

  if (MemInitFile != "") begin : gen_meminit
      $display("Initializing memory %m from file '%s'.", MemInitFile);
      $readmemh(MemInitFile, mem);
  end
end


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Macro bodies included by prim_assert.sv for tools that don't support assertions. See
// prim_assert.sv for documentation for each of the macros.

`define ASSERT_I(__name, __prop)
`define ASSERT_INIT(__name, __prop)
`define ASSERT_INIT_NET(__name, __prop)
`define ASSERT_FINAL(__name, __prop)
`define ASSERT_AT_RESET(__name, __prop, __rst = `ASSERT_DEFAULT_RST)
`define ASSERT_AT_RESET_AND_FINAL(__name, __prop, __rst = `ASSERT_DEFAULT_RST)
`define ASSERT(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST)
`define ASSERT_NEVER(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST)
`define ASSERT_KNOWN(__name, __sig, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST)
`define COVER(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST)
`define ASSUME(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST)
`define ASSUME_I(__name, __prop)


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Macro bodies included by prim_assert.sv for tools that support full SystemVerilog and SVA syntax.
// See prim_assert.sv for documentation for each of the macros.

`define ASSERT_I(__name, __prop) \
  __name: assert (__prop)        \
    else begin                   \
      `ASSERT_ERROR(__name)      \
    end

// Formal tools will ignore the initial construct, so use static assertion as a workaround.
// This workaround terminates design elaboration if the __prop predict is false.
// It calls $fatal() with the first argument equal to 2, it outputs the statistics about the memory
// and CPU time.
`define ASSERT_INIT(__name, __prop)                                                  \
`ifdef FPV_ON                                                                        \
  if (!(__prop)) $fatal(2, "Fatal static assertion [%s]: (%s) is not true.",         \
                        (__name), (__prop));                                         \
`else                                                                                \
  initial begin                                                                      \
    __name: assert (__prop)                                                          \
      else begin                                                                     \
        `ASSERT_ERROR(__name)                                                        \
      end                                                                            \
  end                                                                                \
`endif

`define ASSERT_INIT_NET(__name, __prop)                                                   \
  initial begin                                                                      \
    // When a net is assigned with a value, the assignment is evaluated after        \
    // initial in Xcelium. Add 1ps delay to check value after the assignment is      \
    // completed.                                                                    \
    #1ps;                                                                            \
    __name: assert (__prop)                                                          \
      else begin                                                                     \
        `ASSERT_ERROR(__name)                                                        \
      end                                                                            \
  end                                                                                \

`define ASSERT_FINAL(__name, __prop)                                         \
  final begin                                                                \
    __name: assert (__prop || $test$plusargs("disable_assert_final_checks")) \
      else begin                                                             \
        `ASSERT_ERROR(__name)                                                \
      end                                                                    \
  end

`define ASSERT_AT_RESET(__name, __prop, __rst = `ASSERT_DEFAULT_RST)         \
  // `__rst` is active-high for these macros, so trigger on its posedge.     \
  // The values inside the property are sampled just before the trigger,     \
  // which is necessary to make the evaluation of `__prop` on a reset edge   \
  // meaningful.  On any reset posedge at the start of time, `__rst` itself  \
  // is unknown, and at that time `__prop` is likely not initialized either, \
  // so this assertion does not evaluate `__prop` when `__rst` is unknown.   \
  __name: assert property (@(posedge __rst) $isunknown(__rst) || (__prop))   \
    else begin                                                               \
      `ASSERT_ERROR(__name)                                                  \
    end

`define ASSERT_AT_RESET_AND_FINAL(__name, __prop, __rst = `ASSERT_DEFAULT_RST) \
    `ASSERT_AT_RESET(AtReset_``__name``, __prop, __rst)                        \
    `ASSERT_FINAL(Final_``__name``, __prop)

`define ASSERT(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  __name: assert property (@(posedge __clk) disable iff ((__rst) !== '0) (__prop))       \
    else begin                                                                           \
      `ASSERT_ERROR(__name)                                                              \
    end

`define ASSERT_NEVER(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  __name: assert property (@(posedge __clk) disable iff ((__rst) !== '0) not (__prop))         \
    else begin                                                                                 \
      `ASSERT_ERROR(__name)                                                                    \
    end

`define ASSERT_KNOWN(__name, __sig, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  `ASSERT(__name, !$isunknown(__sig), __clk, __rst)

`define COVER(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  __name: cover property (@(posedge __clk) disable iff ((__rst) !== '0) (__prop));

`define ASSUME(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  __name: assume property (@(posedge __clk) disable iff ((__rst) !== '0) (__prop))       \
    else begin                                                                           \
      `ASSERT_ERROR(__name)                                                              \
    end

`define ASSUME_I(__name, __prop) \
  __name: assume (__prop)        \
    else begin                   \
      `ASSERT_ERROR(__name)      \
    end


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Macro bodies included by prim_assert.sv for formal verification with Yosys. See prim_assert.sv
// for documentation for each of the macros.

`define ASSERT_I(__name, __prop)    \
  always_comb begin : __name        \
    assert (__prop);                \
  end

`define ASSERT_INIT(__name, __prop)    \
  initial begin : __name               \
    assert (__prop);                   \
  end

`define ASSERT_INIT_NET(__name, __prop) \
  initial begin : __name                \
    #1ps assert (__prop);               \
  end

// This doesn't make much sense for a formal tool (we never get to the final block!)
`define ASSERT_FINAL(__name, __prop)

// This needs sampling just before reset assertion and thus requires an event scheduler, which Yosys
// may or may not implement, so we leave it blank for the time being.
`define ASSERT_AT_RESET(__name, __prop, __rst = `ASSERT_DEFAULT_RST)

`define ASSERT_AT_RESET_AND_FINAL(__name, __prop, __rst = `ASSERT_DEFAULT_RST) \
  `ASSERT_AT_RESET(AtReset_``__name``, __prop, __rst)                          \
  `ASSERT_FINAL(Final_``__name``, __prop)

`define ASSERT(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  always_ff @(posedge __clk) begin                                                       \
    if (! (__rst !== '0)) __name: assert (__prop);                                       \
  end

`define ASSERT_NEVER(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  always_ff @(posedge __clk) begin                                                             \
    if (! (__rst !== '0)) __name: assert (! (__prop));                                         \
  end

// Yosys uses 2-state logic, so this doesn't make sense here
`define ASSERT_KNOWN(__name, __sig, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST)

`define COVER(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  always_ff @(posedge __clk) begin : __name                                             \
    cover ((! (__rst !== '0)) && (__prop));                                             \
  end

`define ASSUME(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  always_ff @(posedge __clk) begin                                                       \
    if (! (__rst !== '0)) __name: assume (__prop);                                       \
  end

`define ASSUME_I(__name, __prop)              \
  always_comb begin : __name                  \
    assume (__prop);                          \
  end


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// // Macros and helper code for security countermeasures.

`ifndef PRIM_ASSERT_SEC_CM_SVH
`define PRIM_ASSERT_SEC_CM_SVH

`define _SEC_CM_ALERT_MAX_CYC 30

// Helper macros
`define ASSERT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_, MAX_CYCLES_, ERR_NAME_) \
  `ASSERT(FpvSecCm``NAME_``, \
          $rose(PRIM_HIER_.ERR_NAME_) && !(GATE_) \
          |-> ##[0:MAX_CYCLES_] (ALERT_.alert_p)) \
  `ifdef INC_ASSERT \
  assign PRIM_HIER_.unused_assert_connected = 1'b1; \
  `endif \
  `ASSUME_FPV(``NAME_``TriggerAfterAlertInit_S, $stable(rst_ni) == 0 |-> \
              PRIM_HIER_.ERR_NAME_ == 0 [*10])

`define ASSERT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_, MAX_CYCLES_, ERR_NAME_, CLK_, RST_) \
  `ASSERT(FpvSecCm``NAME_``, \
          $rose(PRIM_HIER_.ERR_NAME_) && !(GATE_) \
          |-> ##[0:MAX_CYCLES_] (ERR_), CLK_, RST_) \
  `ifdef INC_ASSERT \
  assign PRIM_HIER_.unused_assert_connected = 1'b1; \
  `endif

// macros for security countermeasures that will trigger alert
`define ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC) \
  `ASSERT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_, MAX_CYCLES_, err_o)

`define ASSERT_PRIM_DOUBLE_LFSR_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC) \
  `ASSERT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_, MAX_CYCLES_, err_o)

`define ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC) \
  `ASSERT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_, MAX_CYCLES_, unused_err_o)

`define ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC) \
  `ASSERT_ERROR_TRIGGER_ALERT(NAME_, PRIM_HIER_, ALERT_, GATE_, MAX_CYCLES_, err_o)

`define ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(NAME_, REG_TOP_HIER_, ALERT_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC) \
  `ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ALERT(NAME_, \
    REG_TOP_HIER_.u_prim_reg_we_check.u_prim_onehot_check, ALERT_, GATE_, MAX_CYCLES_)

// macros for security countermeasures that will trigger other errors
`define ASSERT_PRIM_FSM_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_ = 0, MAX_CYCLES_ = 2, CLK_ = clk_i, RST_ = !rst_ni) \
  `ASSERT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_, MAX_CYCLES_, unused_err_o, CLK_, RST_)

`define ASSERT_PRIM_COUNT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_ = 0, MAX_CYCLES_ = 2, CLK_ = clk_i, RST_ = !rst_ni) \
  `ASSERT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_, MAX_CYCLES_, err_o, CLK_, RST_)

`define ASSERT_PRIM_DOUBLE_LFSR_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_ = 0, MAX_CYCLES_ = 2, CLK_ = clk_i, RST_ = !rst_ni) \
  `ASSERT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_, MAX_CYCLES_, err_o, CLK_, RST_)

`define ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC, CLK_ = clk_i, RST_ = !rst_ni) \
  `ASSERT_ERROR_TRIGGER_ERR(NAME_, PRIM_HIER_, ERR_, GATE_, MAX_CYCLES_, err_o, CLK_, RST_)

`define ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ERR(NAME_, REG_TOP_HIER_, ERR_, GATE_ = 0, MAX_CYCLES_ = `_SEC_CM_ALERT_MAX_CYC, CLK_ = clk_i, RST_ = !rst_ni) \
  `ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ERR(NAME_, \
    REG_TOP_HIER_.u_prim_reg_we_check.u_prim_onehot_check, ERR_, GATE_, MAX_CYCLES_, CLK_, RST_)

`endif // PRIM_ASSERT_SEC_CM_SVH


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`ifndef PRIM_FLOP_MACROS_SV
`define PRIM_FLOP_MACROS_SV

/////////////////////////////////////
// Default Values for Macros below //
/////////////////////////////////////

`define PRIM_FLOP_CLK clk_i
`define PRIM_FLOP_RST rst_ni
`define PRIM_FLOP_RESVAL '0

/////////////////////
// Register Macros //
/////////////////////

// TODO: define other variations of register macros so that they can be used throughout all designs
// to make the code more concise.

// Register with asynchronous reset.
`define PRIM_FLOP_A(__d, __q, __resval = `PRIM_FLOP_RESVAL, __clk = `PRIM_FLOP_CLK, __rst_n = `PRIM_FLOP_RST) \
  always_ff @(posedge __clk or negedge __rst_n) begin \
    if (!__rst_n) begin                               \
      __q <= __resval;                                \
    end else begin                                    \
      __q <= __d;                                     \
    end                                               \
  end

///////////////////////////
// Macro for Sparse FSMs //
///////////////////////////

// Simulation tools typically infer FSMs and report coverage for these separately. However, tools
// like Xcelium and VCS seem to have problems inferring FSMs if the state register is not coded in
// a behavioral always_ff block in the same hierarchy. To that end, this uses a modified variant
// with a second behavioral register definition for RTL simulations so that FSMs can be inferred.
// Note that in this variant, the __q output is disconnected from prim_sparse_fsm_flop and attached
// to the behavioral flop. An assertion is added to ensure equivalence between the
// prim_sparse_fsm_flop output and the behavioral flop output in that case.
`define PRIM_FLOP_SPARSE_FSM(__name, __d, __q, __type, __resval = `PRIM_FLOP_RESVAL, __clk = `PRIM_FLOP_CLK, __rst_n = `PRIM_FLOP_RST, __alert_trigger_sva_en = 1) \
  `ifdef SIMULATION                                   \
    prim_sparse_fsm_flop #(                           \
      .StateEnumT(__type),                            \
      .Width($bits(__type)),                          \
      .ResetValue($bits(__type)'(__resval)),          \
      .EnableAlertTriggerSVA(__alert_trigger_sva_en), \
      .CustomForceName(`PRIM_STRINGIFY(__q))          \
    ) __name (                                        \
      .clk_i   ( __clk   ),                           \
      .rst_ni  ( __rst_n ),                           \
      .state_i ( __d     ),                           \
      .state_o (         )                            \
    );                                                \
    `PRIM_FLOP_A(__d, __q, __resval, __clk, __rst_n)  \
    `ASSERT(``__name``_A, __q === ``__name``.state_o) \
  `else                                               \
    prim_sparse_fsm_flop #(                           \
      .StateEnumT(__type),                            \
      .Width($bits(__type)),                          \
      .ResetValue($bits(__type)'(__resval)),          \
      .EnableAlertTriggerSVA(__alert_trigger_sva_en)  \
    ) __name (                                        \
      .clk_i   ( __clk   ),                           \
      .rst_ni  ( __rst_n ),                           \
      .state_i ( __d     ),                           \
      .state_o ( __q     )                            \
    );                                                \
  `endif

`endif // PRIM_FLOP_MACROS_SV


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Macros and helper code for using assertions.
//  - Provides default clk and rst options to simplify code
//  - Provides boiler plate template for common assertions

`ifndef PRIM_ASSERT_SV
`define PRIM_ASSERT_SV

///////////////////
// Helper macros //
///////////////////

// Default clk and reset signals used by assertion macros below.
`define ASSERT_DEFAULT_CLK clk_i
`define ASSERT_DEFAULT_RST !rst_ni

// Converts an arbitrary block of code into a Verilog string
`define PRIM_STRINGIFY(__x) `"__x`"

// ASSERT_ERROR logs an error message with either `uvm_error or with $error.
//
// This somewhat duplicates `DV_ERROR macro defined in hw/dv/sv/dv_utils/dv_macros.svh. The reason
// for redefining it here is to avoid creating a dependency.
`define ASSERT_ERROR(__name)                                                             \
`ifdef UVM                                                                               \
  uvm_pkg::uvm_report_error("ASSERT FAILED", `PRIM_STRINGIFY(__name), uvm_pkg::UVM_NONE, \
                            `__FILE__, `__LINE__, "", 1);                                \
`else                                                                                    \
  $error("%0t: (%0s:%0d) [%m] [ASSERT FAILED] %0s", $time, `__FILE__, `__LINE__,         \
         `PRIM_STRINGIFY(__name));                                                       \
`endif

// This macro is suitable for conditionally triggering lint errors, e.g., if a Sec parameter takes
// on a non-default value. This may be required for pre-silicon/FPGA evaluation but we don't want
// to allow this for tapeout.
`define ASSERT_STATIC_LINT_ERROR(__name, __prop)     \
  localparam int __name = (__prop) ? 1 : 2;          \
  always_comb begin                                  \
    logic unused_assert_static_lint_error;           \
    unused_assert_static_lint_error = __name'(1'b1); \
  end

// Static assertions for checks inside SV packages. If the conditions is not true, this will
// trigger an error during elaboration.
`define ASSERT_STATIC_IN_PACKAGE(__name, __prop)              \
  function automatic bit assert_static_in_package_``__name(); \
    bit unused_bit [((__prop) ? 1 : -1)];                     \
    unused_bit = '{default: 1'b0};                            \
    return unused_bit[0];                                     \
  endfunction

// The basic helper macros are actually defined in "implementation headers". The macros should do
// the same thing in each case (except for the dummy flavour), but in a way that the respective
// tools support.
//
// If the tool supports assertions in some form, we also define INC_ASSERT (which can be used to
// hide signal definitions that are only used for assertions).
//
// The list of basic macros supported is:
//
//  ASSERT_I:     Immediate assertion. Note that immediate assertions are sensitive to simulation
//                glitches.
//
//  ASSERT_INIT:  Assertion in initial block. Can be used for things like parameter checking.
//
//  ASSERT_INIT_NET: Assertion in initial block. Can be used for initial value of a net.
//
//  ASSERT_FINAL: Assertion in final block. Can be used for things like queues being empty at end of
//                sim, all credits returned at end of sim, state machines in idle at end of sim.
//
//  ASSERT_AT_RESET: Assertion just before reset. Can be used to check sum-like properties that get
//                   cleared at reset.
//                   Note that unless your simulation ends with a reset, the property does not get
//                   checked at end of simulation; use ASSERT_AT_RESET_AND_FINAL if the property
//                   should also get checked at end of simulation.
//
//  ASSERT_AT_RESET_AND_FINAL: Assertion just before reset and in final block. Can be used to check
//                             sum-like properties before every reset and at the end of simulation.
//
//  ASSERT:       Assert a concurrent property directly. It can be called as a module (or
//                interface) body item.
//
//                Note: We use (__rst !== '0) in the disable iff statements instead of (__rst ==
//                '1). This properly disables the assertion in cases when reset is X at the
//                beginning of a simulation. For that case, (reset == '1) does not disable the
//                assertion.
//
//  ASSERT_NEVER: Assert a concurrent property NEVER happens
//
//  ASSERT_KNOWN: Assert that signal has a known value (each bit is either '0' or '1') after reset.
//                It can be called as a module (or interface) body item.
//
//  COVER:        Cover a concurrent property
//
//  ASSUME:       Assume a concurrent property
//
//  ASSUME_I:     Assume an immediate property

`ifdef VERILATOR
 `include "prim_assert_dummy_macros.svh"
`elsif SYNTHESIS
 `include "prim_assert_dummy_macros.svh"
`elsif YOSYS
 `include "prim_assert_yosys_macros.svh"
 `define INC_ASSERT
`else
 `include "prim_assert_dummy_macros.svh"
//  `define INC_ASSERT
`endif

//////////////////////////////
// Complex assertion macros //
//////////////////////////////

// Assert that signal is an active-high pulse with pulse length of 1 clock cycle
`define ASSERT_PULSE(__name, __sig, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  `ASSERT(__name, $rose(__sig) |=> !(__sig), __clk, __rst)

// Assert that a property is true only when an enable signal is set.  It can be called as a module
// (or interface) body item.
`define ASSERT_IF(__name, __prop, __enable, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  `ASSERT(__name, (__enable) |-> (__prop), __clk, __rst)

// Assert that signal has a known value (each bit is either '0' or '1') after reset if enable is
// set.  It can be called as a module (or interface) body item.
`define ASSERT_KNOWN_IF(__name, __sig, __enable, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  `ASSERT_KNOWN(__name``KnownEnable, __enable, __clk, __rst)                                               \
  `ASSERT_IF(__name, !$isunknown(__sig), __enable, __clk, __rst)

//////////////////////////////////
// For formal verification only //
//////////////////////////////////

// Note that the existing set of ASSERT macros specified above shall be used for FPV,
// thereby ensuring that the assertions are evaluated during DV simulations as well.

// ASSUME_FPV
// Assume a concurrent property during formal verification only.
`define ASSUME_FPV(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
`ifdef FPV_ON                                                                                \
   `ASSUME(__name, __prop, __clk, __rst)                                                     \
`endif

// ASSUME_I_FPV
// Assume a concurrent property during formal verification only.
`define ASSUME_I_FPV(__name, __prop) \
`ifdef FPV_ON                        \
   `ASSUME_I(__name, __prop)         \
`endif

// COVER_FPV
// Cover a concurrent property during formal verification
`define COVER_FPV(__name, __prop, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
`ifdef FPV_ON                                                                               \
   `COVER(__name, __prop, __clk, __rst)                                                     \
`endif

// FPV assertion that proves that the FSM control flow is linear (no loops)
// The sequence triggers whenever the state changes and stores the current state as "initial_state".
// Then thereafter we must never see that state again until reset.
// It is possible for the reset to release ahead of the clock.
// Create a small "gray" window beyond the usual rst time to avoid
// checking.
`define ASSERT_FPV_LINEAR_FSM(__name, __state, __type, __clk = `ASSERT_DEFAULT_CLK, __rst = `ASSERT_DEFAULT_RST) \
  `ifdef INC_ASSERT                                                                                              \
     bit __name``_cond;                                                                                          \
     always_ff @(posedge __clk or posedge __rst) begin                                                           \
       if (__rst) begin                                                                                          \
         __name``_cond <= 0;                                                                                     \
       end else begin                                                                                            \
         __name``_cond <= 1;                                                                                     \
       end                                                                                                       \
     end                                                                                                         \
     property __name``_p;                                                                                        \
       __type initial_state;                                                                                     \
       (!$stable(__state) & __name``_cond, initial_state = $past(__state)) |->                                   \
           (__state != initial_state) until (__rst == 1'b1);                                                     \
     endproperty                                                                                                 \
   `ASSERT(__name, __name``_p, __clk, __rst)                                                                     \
  `endif

`include "prim_assert_sec_cm.svh"
`include "prim_flop_macros.sv"

`endif // PRIM_ASSERT_SV


// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/19 
// Design Name: sm3
// Module Name: sm3_cfg
// Description:
//      SM3 模块配置信息
// Dependencies: 
//      
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
//定义设计阶段-----------------------------
//`define DESIGN_SIM
// `define DESIGN_SYNT

//模块调试开关-----------------------------
`ifdef  DESIGN_SIM
    //`define SM3_PAD_SIM_DBG
    // `define SM3_EXPND_SIM_DBG
    `define SM3_CMPRS_SIM_DBG
    // `define SM3_CMPRS_SIM_FILE_LOG
`endif

//C模型相关设置----------------------------
// `define C_MODEL_SELF_TEST

//定义 SM3 输入位宽------------------------
`define SM3_INPT_DW_32
`ifndef  SM3_INPT_DW_32
    `define SM3_INPT_DW_64
`endif

`ifdef SM3_INPT_DW_32
    `define     INPT_DW    32
`elsif SM3_INPT_DW_64
    `define     INPT_DW    64
`endif

// `define INPT_DW1        (INPT_DW - 1)
`define INPT_DW1        (`INPT_DW - 1)
`define INPT_BYTE_DW1   (`INPT_DW/8 - 1)
`define INPT_BYTE_DW    (`INPT_BYTE_DW1 + 1)

//定义 SM3 输出位宽-------------------------
// `define SM3_OTPT_DW_32
//`define SM3_OTPT_DW_64
// `define SM3_OTPT_DW_128
`define SM3_OTPT_DW_256

`ifdef SM3_OTPT_DW_32
    `define     OTPT_DW    32
`elsif SM3_OTPT_DW_64
    `define     OTPT_DW    64
`elsif SM3_OTPT_DW_128
    `define     OTPT_DW    128
`elsif SM3_OTPT_DW_256
    `define     OTPT_DW    256
`endif

`define OTPT_DW1 (OTPT_DW - 1)

//定义 SM3 字扩展模式-----------------------
`define SM3_EXPND_PRE_LOAD_REG

//定义 SM3 迭代压缩中的加法方式-----------------------
//直接使用加法符，使工具推断
//`define SM3_CMPRSS_DIRECT_ADD
//显式例化 CSA 加法器 在 SM3_CMPRSS_DIRECT_ADD 未定义时有效
`ifndef  SM3_CMPRSS_DIRECT_ADD
    `define SM3_CMPRSS_CSA_ADD
`endif

//定义仿真器 define simulator
// Modelsim_10_5(windows), default 
// EpicSim (Linux)
//`define EPICSIM
`ifndef EPICSIM
    `define MODELSIM_10_5
`endif

//定义是否使用 C 语言参考模型(DPI)
//define using C reference model or not
//`define C_MODEL_ENABLE

//定义是否 dump 波形
//define dump wave in VCD or not
//`define VCD_DUMP_ENABLE

`define WIDTH  256

//`define FPGA



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Some generally useful macros for RTL.

// Determine if __actual equals __expected with a margin of __allowed_less and __allowed_more, i.e.,
// if __actual is in the interval [__expected - __allowed_less, __expected + __allowed_more], where
// lower and upper bounds are inclusive.
//
// The caller is responsible for ensuring that the data types are such that
// (1) __actual + __allowed_less
// (2) __expected + __allowed_more
// are well defined and do not overflow and
// (3) (1) >= __expected
// (4) __actual <= (2)
// are well defined and meaningful.  Subtractions are deliberately not used, in order to prevent
// underflows.
`define WITHIN_MARGIN(__actual, __expected, __allowed_less, __allowed_more) \
  (((__actual) + (__allowed_less) >= (__expected)) &&                       \
   ((__actual) <= (__expected) + (__allowed_more)))

// Coverage pragmas, used around code for which we want to disable coverage collection.
// Don't forget to add a closing ON pragma after the code to be skipped.
//
// Some notes:
// - The first line is for VCS, the second for xcelium. It is okay to issue both regardless of
//   the tool used.
// - For xcelium it is possible to discriminate between metrics to be disabled as follows
//   //pragma coverage <metric> = on/off
//   where metric can be block | expr | toggle | fsm.

// TODO(https://github.com/chipsalliance/verible/issues/1498) Verible seems to get confused
// by these macros, so the code will inline these directives until this is fixed.
/*
`ifndef PRAGMA_COVERAGE_OFF
`define PRAGMA_COVERAGE_OFF \
/``/VCS coverage off \
/``/ pragma coverage off
`endif

`ifndef PRAGMA_COVERAGE_ON
`define PRAGMA_COVERAGE_ON \
/``/VCS coverage on \
/``/ pragma coverage on
`endif
*/


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package flash_ctrl_reg_pkg;

  // Param list
  parameter int RegNumBanks = 2;
  parameter int RegPagesPerBank = 256;
  parameter int RegBusPgmResBytes = 64;
  parameter int RegPageWidth = 8;
  parameter int RegBankWidth = 1;
  parameter int NumRegions = 8;
  parameter int NumInfoTypes = 3;
  parameter int NumInfos0 = 10;
  parameter int NumInfos1 = 1;
  parameter int NumInfos2 = 2;
  parameter int WordsPerPage = 256;
  parameter int BytesPerWord = 8;
  parameter int BytesPerPage = 2048;
  parameter int BytesPerBank = 524288;
  parameter int unsigned ExecEn = 32'ha26a38f7;
  parameter int MaxFifoDepth = 16;
  parameter int MaxFifoWidth = 5;
  parameter int NumAlerts = 5;

  // Address widths within the block
  parameter int CoreAw = 9;
  parameter int PrimAw = 7;
  parameter int MemAw = 1;

  ///////////////////////////////////////////////
  // Typedefs for registers for core interface //
  ///////////////////////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } prog_empty;
    struct packed {
      logic        q;
    } prog_lvl;
    struct packed {
      logic        q;
    } rd_full;
    struct packed {
      logic        q;
    } rd_lvl;
    struct packed {
      logic        q;
    } op_done;
    struct packed {
      logic        q;
    } corr_err;
  } flash_ctrl_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } prog_empty;
    struct packed {
      logic        q;
    } prog_lvl;
    struct packed {
      logic        q;
    } rd_full;
    struct packed {
      logic        q;
    } rd_lvl;
    struct packed {
      logic        q;
    } op_done;
    struct packed {
      logic        q;
    } corr_err;
  } flash_ctrl_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } prog_empty;
    struct packed {
      logic        q;
      logic        qe;
    } prog_lvl;
    struct packed {
      logic        q;
      logic        qe;
    } rd_full;
    struct packed {
      logic        q;
      logic        qe;
    } rd_lvl;
    struct packed {
      logic        q;
      logic        qe;
    } op_done;
    struct packed {
      logic        q;
      logic        qe;
    } corr_err;
  } flash_ctrl_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_err;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_std_err;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_err;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_prim_flash_alert;
    struct packed {
      logic        q;
      logic        qe;
    } recov_prim_flash_alert;
  } flash_ctrl_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic [3:0]  q;
  } flash_ctrl_reg2hw_dis_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } flash_ctrl_reg2hw_exec_reg_t;

  typedef struct packed {
    logic        q;
  } flash_ctrl_reg2hw_init_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } start;
    struct packed {
      logic [1:0]  q;
    } op;
    struct packed {
      logic        q;
    } prog_sel;
    struct packed {
      logic        q;
    } erase_sel;
    struct packed {
      logic        q;
    } partition_sel;
    struct packed {
      logic [1:0]  q;
    } info_sel;
    struct packed {
      logic [11:0] q;
    } num;
  } flash_ctrl_reg2hw_control_reg_t;

  typedef struct packed {
    logic [19:0] q;
  } flash_ctrl_reg2hw_addr_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } normal;
    struct packed {
      logic        q;
    } repair;
  } flash_ctrl_reg2hw_prog_type_en_reg_t;

  typedef struct packed {
    logic        q;
  } flash_ctrl_reg2hw_erase_suspend_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_mp_region_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [8:0]  q;
    } base;
    struct packed {
      logic [9:0] q;
    } size;
  } flash_ctrl_reg2hw_mp_region_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_default_region_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_bank0_info0_page_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_bank0_info1_page_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_bank0_info2_page_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_bank1_info0_page_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_bank1_info1_page_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } en;
    struct packed {
      logic [3:0]  q;
    } rd_en;
    struct packed {
      logic [3:0]  q;
    } prog_en;
    struct packed {
      logic [3:0]  q;
    } erase_en;
    struct packed {
      logic [3:0]  q;
    } scramble_en;
    struct packed {
      logic [3:0]  q;
    } ecc_en;
    struct packed {
      logic [3:0]  q;
    } he_en;
  } flash_ctrl_reg2hw_bank1_info2_page_cfg_mreg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } scramble_dis;
    struct packed {
      logic [3:0]  q;
    } ecc_dis;
  } flash_ctrl_reg2hw_hw_info_cfg_override_reg_t;

  typedef struct packed {
    logic        q;
  } flash_ctrl_reg2hw_mp_bank_cfg_shadowed_mreg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } reg_intg_err;
    struct packed {
      logic        q;
    } prog_intg_err;
    struct packed {
      logic        q;
    } lcmgr_err;
    struct packed {
      logic        q;
    } lcmgr_intg_err;
    struct packed {
      logic        q;
    } arb_fsm_err;
    struct packed {
      logic        q;
    } storage_err;
    struct packed {
      logic        q;
    } phy_fsm_err;
    struct packed {
      logic        q;
    } ctrl_cnt_err;
    struct packed {
      logic        q;
    } fifo_err;
  } flash_ctrl_reg2hw_std_fault_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } op_err;
    struct packed {
      logic        q;
    } mp_err;
    struct packed {
      logic        q;
    } rd_err;
    struct packed {
      logic        q;
    } prog_err;
    struct packed {
      logic        q;
    } prog_win_err;
    struct packed {
      logic        q;
    } prog_type_err;
    struct packed {
      logic        q;
    } seed_err;
    struct packed {
      logic        q;
    } phy_relbl_err;
    struct packed {
      logic        q;
    } phy_storage_err;
    struct packed {
      logic        q;
    } spurious_ack;
    struct packed {
      logic        q;
    } arb_err;
    struct packed {
      logic        q;
    } host_gnt_err;
  } flash_ctrl_reg2hw_fault_status_reg_t;

  typedef struct packed {
    logic [7:0]  q;
  } flash_ctrl_reg2hw_ecc_single_err_cnt_mreg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } alert_ack;
    struct packed {
      logic        q;
    } alert_trig;
  } flash_ctrl_reg2hw_phy_alert_cfg_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } flash_ctrl_reg2hw_scratch_reg_t;

  typedef struct packed {
    struct packed {
      logic [4:0]  q;
    } prog;
    struct packed {
      logic [4:0]  q;
    } rd;
  } flash_ctrl_reg2hw_fifo_lvl_reg_t;

  typedef struct packed {
    logic        q;
  } flash_ctrl_reg2hw_fifo_rst_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } prog_empty;
    struct packed {
      logic        d;
      logic        de;
    } prog_lvl;
    struct packed {
      logic        d;
      logic        de;
    } rd_full;
    struct packed {
      logic        d;
      logic        de;
    } rd_lvl;
    struct packed {
      logic        d;
      logic        de;
    } op_done;
    struct packed {
      logic        d;
      logic        de;
    } corr_err;
  } flash_ctrl_hw2reg_intr_state_reg_t;

  typedef struct packed {
    logic        d;
  } flash_ctrl_hw2reg_ctrl_regwen_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } start;
  } flash_ctrl_hw2reg_control_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } flash_ctrl_hw2reg_erase_suspend_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } done;
    struct packed {
      logic        d;
      logic        de;
    } err;
  } flash_ctrl_hw2reg_op_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } rd_full;
    struct packed {
      logic        d;
      logic        de;
    } rd_empty;
    struct packed {
      logic        d;
      logic        de;
    } prog_full;
    struct packed {
      logic        d;
      logic        de;
    } prog_empty;
    struct packed {
      logic        d;
      logic        de;
    } init_wip;
    struct packed {
      logic        d;
      logic        de;
    } initialized;
  } flash_ctrl_hw2reg_status_reg_t;

  typedef struct packed {
    logic [10:0] d;
  } flash_ctrl_hw2reg_debug_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } op_err;
    struct packed {
      logic        d;
      logic        de;
    } mp_err;
    struct packed {
      logic        d;
      logic        de;
    } rd_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_win_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_type_err;
    struct packed {
      logic        d;
      logic        de;
    } update_err;
    struct packed {
      logic        d;
      logic        de;
    } macro_err;
  } flash_ctrl_hw2reg_err_code_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } reg_intg_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_intg_err;
    struct packed {
      logic        d;
      logic        de;
    } lcmgr_err;
    struct packed {
      logic        d;
      logic        de;
    } lcmgr_intg_err;
    struct packed {
      logic        d;
      logic        de;
    } arb_fsm_err;
    struct packed {
      logic        d;
      logic        de;
    } storage_err;
    struct packed {
      logic        d;
      logic        de;
    } phy_fsm_err;
    struct packed {
      logic        d;
      logic        de;
    } ctrl_cnt_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_err;
  } flash_ctrl_hw2reg_std_fault_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } op_err;
    struct packed {
      logic        d;
      logic        de;
    } mp_err;
    struct packed {
      logic        d;
      logic        de;
    } rd_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_win_err;
    struct packed {
      logic        d;
      logic        de;
    } prog_type_err;
    struct packed {
      logic        d;
      logic        de;
    } seed_err;
    struct packed {
      logic        d;
      logic        de;
    } phy_relbl_err;
    struct packed {
      logic        d;
      logic        de;
    } phy_storage_err;
    struct packed {
      logic        d;
      logic        de;
    } spurious_ack;
    struct packed {
      logic        d;
      logic        de;
    } arb_err;
    struct packed {
      logic        d;
      logic        de;
    } host_gnt_err;
  } flash_ctrl_hw2reg_fault_status_reg_t;

  typedef struct packed {
    logic [19:0] d;
    logic        de;
  } flash_ctrl_hw2reg_err_addr_reg_t;

  typedef struct packed {
    logic [7:0]  d;
    logic        de;
  } flash_ctrl_hw2reg_ecc_single_err_cnt_mreg_t;

  typedef struct packed {
    logic [19:0] d;
    logic        de;
  } flash_ctrl_hw2reg_ecc_single_err_addr_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } init_wip;
    struct packed {
      logic        d;
      logic        de;
    } prog_normal_avail;
    struct packed {
      logic        d;
      logic        de;
    } prog_repair_avail;
  } flash_ctrl_hw2reg_phy_status_reg_t;

  typedef struct packed {
    struct packed {
      logic [4:0]  d;
    } prog;
    struct packed {
      logic [4:0]  d;
    } rd;
  } flash_ctrl_hw2reg_curr_fifo_lvl_reg_t;

  // Register -> HW type for core interface
  typedef struct packed {
    flash_ctrl_reg2hw_intr_state_reg_t intr_state; // [1333:1328]
    flash_ctrl_reg2hw_intr_enable_reg_t intr_enable; // [1327:1322]
    flash_ctrl_reg2hw_intr_test_reg_t intr_test; // [1321:1310]
    flash_ctrl_reg2hw_alert_test_reg_t alert_test; // [1309:1300]
    flash_ctrl_reg2hw_dis_reg_t dis; // [1299:1296]
    flash_ctrl_reg2hw_exec_reg_t exec; // [1295:1264]
    flash_ctrl_reg2hw_init_reg_t init; // [1263:1263]
    flash_ctrl_reg2hw_control_reg_t control; // [1262:1243]
    flash_ctrl_reg2hw_addr_reg_t addr; // [1242:1223]
    flash_ctrl_reg2hw_prog_type_en_reg_t prog_type_en; // [1222:1221]
    flash_ctrl_reg2hw_erase_suspend_reg_t erase_suspend; // [1220:1220]
    flash_ctrl_reg2hw_mp_region_cfg_mreg_t [7:0] mp_region_cfg; // [1219:996]
    flash_ctrl_reg2hw_mp_region_mreg_t [7:0] mp_region; // [995:844]
    flash_ctrl_reg2hw_default_region_reg_t default_region; // [843:820]
    flash_ctrl_reg2hw_bank0_info0_page_cfg_mreg_t [9:0] bank0_info0_page_cfg; // [819:540]
    flash_ctrl_reg2hw_bank0_info1_page_cfg_mreg_t [0:0] bank0_info1_page_cfg; // [539:512]
    flash_ctrl_reg2hw_bank0_info2_page_cfg_mreg_t [1:0] bank0_info2_page_cfg; // [511:456]
    flash_ctrl_reg2hw_bank1_info0_page_cfg_mreg_t [9:0] bank1_info0_page_cfg; // [455:176]
    flash_ctrl_reg2hw_bank1_info1_page_cfg_mreg_t [0:0] bank1_info1_page_cfg; // [175:148]
    flash_ctrl_reg2hw_bank1_info2_page_cfg_mreg_t [1:0] bank1_info2_page_cfg; // [147:92]
    flash_ctrl_reg2hw_hw_info_cfg_override_reg_t hw_info_cfg_override; // [91:84]
    flash_ctrl_reg2hw_mp_bank_cfg_shadowed_mreg_t [1:0] mp_bank_cfg_shadowed; // [83:82]
    flash_ctrl_reg2hw_std_fault_status_reg_t std_fault_status; // [81:73]
    flash_ctrl_reg2hw_fault_status_reg_t fault_status; // [72:61]
    flash_ctrl_reg2hw_ecc_single_err_cnt_mreg_t [1:0] ecc_single_err_cnt; // [60:45]
    flash_ctrl_reg2hw_phy_alert_cfg_reg_t phy_alert_cfg; // [44:43]
    flash_ctrl_reg2hw_scratch_reg_t scratch; // [42:11]
    flash_ctrl_reg2hw_fifo_lvl_reg_t fifo_lvl; // [10:1]
    flash_ctrl_reg2hw_fifo_rst_reg_t fifo_rst; // [0:0]
  } flash_ctrl_core_reg2hw_t;

  // HW -> register type for core interface
  typedef struct packed {
    flash_ctrl_hw2reg_intr_state_reg_t intr_state; // [198:187]
    flash_ctrl_hw2reg_ctrl_regwen_reg_t ctrl_regwen; // [186:186]
    flash_ctrl_hw2reg_control_reg_t control; // [185:184]
    flash_ctrl_hw2reg_erase_suspend_reg_t erase_suspend; // [183:182]
    flash_ctrl_hw2reg_op_status_reg_t op_status; // [181:178]
    flash_ctrl_hw2reg_status_reg_t status; // [177:166]
    flash_ctrl_hw2reg_debug_state_reg_t debug_state; // [165:155]
    flash_ctrl_hw2reg_err_code_reg_t err_code; // [154:139]
    flash_ctrl_hw2reg_std_fault_status_reg_t std_fault_status; // [138:121]
    flash_ctrl_hw2reg_fault_status_reg_t fault_status; // [120:97]
    flash_ctrl_hw2reg_err_addr_reg_t err_addr; // [96:76]
    flash_ctrl_hw2reg_ecc_single_err_cnt_mreg_t [1:0] ecc_single_err_cnt; // [75:58]
    flash_ctrl_hw2reg_ecc_single_err_addr_mreg_t [1:0] ecc_single_err_addr; // [57:16]
    flash_ctrl_hw2reg_phy_status_reg_t phy_status; // [15:10]
    flash_ctrl_hw2reg_curr_fifo_lvl_reg_t curr_fifo_lvl; // [9:0]
  } flash_ctrl_core_hw2reg_t;

  // Register offsets for core interface
  parameter logic [CoreAw-1:0] FLASH_CTRL_INTR_STATE_OFFSET = 9'h 0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_INTR_ENABLE_OFFSET = 9'h 4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_INTR_TEST_OFFSET = 9'h 8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ALERT_TEST_OFFSET = 9'h c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_DIS_OFFSET = 9'h 10;
  parameter logic [CoreAw-1:0] FLASH_CTRL_EXEC_OFFSET = 9'h 14;
  parameter logic [CoreAw-1:0] FLASH_CTRL_INIT_OFFSET = 9'h 18;
  parameter logic [CoreAw-1:0] FLASH_CTRL_CTRL_REGWEN_OFFSET = 9'h 1c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_CONTROL_OFFSET = 9'h 20;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ADDR_OFFSET = 9'h 24;
  parameter logic [CoreAw-1:0] FLASH_CTRL_PROG_TYPE_EN_OFFSET = 9'h 28;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ERASE_SUSPEND_OFFSET = 9'h 2c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_0_OFFSET = 9'h 30;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_1_OFFSET = 9'h 34;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_2_OFFSET = 9'h 38;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_3_OFFSET = 9'h 3c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_4_OFFSET = 9'h 40;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_5_OFFSET = 9'h 44;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_6_OFFSET = 9'h 48;
  parameter logic [CoreAw-1:0] FLASH_CTRL_REGION_CFG_REGWEN_7_OFFSET = 9'h 4c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_0_OFFSET = 9'h 50;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_1_OFFSET = 9'h 54;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_2_OFFSET = 9'h 58;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_3_OFFSET = 9'h 5c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_4_OFFSET = 9'h 60;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_5_OFFSET = 9'h 64;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_6_OFFSET = 9'h 68;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_CFG_7_OFFSET = 9'h 6c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_0_OFFSET = 9'h 70;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_1_OFFSET = 9'h 74;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_2_OFFSET = 9'h 78;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_3_OFFSET = 9'h 7c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_4_OFFSET = 9'h 80;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_5_OFFSET = 9'h 84;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_6_OFFSET = 9'h 88;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_REGION_7_OFFSET = 9'h 8c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_DEFAULT_REGION_OFFSET = 9'h 90;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_0_OFFSET = 9'h 94;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_1_OFFSET = 9'h 98;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_2_OFFSET = 9'h 9c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_3_OFFSET = 9'h a0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_4_OFFSET = 9'h a4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_5_OFFSET = 9'h a8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_6_OFFSET = 9'h ac;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_7_OFFSET = 9'h b0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_8_OFFSET = 9'h b4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_REGWEN_9_OFFSET = 9'h b8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_0_OFFSET = 9'h bc;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_1_OFFSET = 9'h c0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_2_OFFSET = 9'h c4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_3_OFFSET = 9'h c8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_4_OFFSET = 9'h cc;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_5_OFFSET = 9'h d0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_6_OFFSET = 9'h d4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_7_OFFSET = 9'h d8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_8_OFFSET = 9'h dc;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_9_OFFSET = 9'h e0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO1_REGWEN_OFFSET = 9'h e4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO1_PAGE_CFG_OFFSET = 9'h e8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO2_REGWEN_0_OFFSET = 9'h ec;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO2_REGWEN_1_OFFSET = 9'h f0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO2_PAGE_CFG_0_OFFSET = 9'h f4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK0_INFO2_PAGE_CFG_1_OFFSET = 9'h f8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_0_OFFSET = 9'h fc;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_1_OFFSET = 9'h 100;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_2_OFFSET = 9'h 104;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_3_OFFSET = 9'h 108;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_4_OFFSET = 9'h 10c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_5_OFFSET = 9'h 110;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_6_OFFSET = 9'h 114;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_7_OFFSET = 9'h 118;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_8_OFFSET = 9'h 11c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_REGWEN_9_OFFSET = 9'h 120;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_0_OFFSET = 9'h 124;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_1_OFFSET = 9'h 128;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_2_OFFSET = 9'h 12c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_3_OFFSET = 9'h 130;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_4_OFFSET = 9'h 134;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_5_OFFSET = 9'h 138;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_6_OFFSET = 9'h 13c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_7_OFFSET = 9'h 140;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_8_OFFSET = 9'h 144;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_9_OFFSET = 9'h 148;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO1_REGWEN_OFFSET = 9'h 14c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO1_PAGE_CFG_OFFSET = 9'h 150;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO2_REGWEN_0_OFFSET = 9'h 154;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO2_REGWEN_1_OFFSET = 9'h 158;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO2_PAGE_CFG_0_OFFSET = 9'h 15c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK1_INFO2_PAGE_CFG_1_OFFSET = 9'h 160;
  parameter logic [CoreAw-1:0] FLASH_CTRL_HW_INFO_CFG_OVERRIDE_OFFSET = 9'h 164;
  parameter logic [CoreAw-1:0] FLASH_CTRL_BANK_CFG_REGWEN_OFFSET = 9'h 168;
  parameter logic [CoreAw-1:0] FLASH_CTRL_MP_BANK_CFG_SHADOWED_OFFSET = 9'h 16c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_OP_STATUS_OFFSET = 9'h 170;
  parameter logic [CoreAw-1:0] FLASH_CTRL_STATUS_OFFSET = 9'h 174;
  parameter logic [CoreAw-1:0] FLASH_CTRL_DEBUG_STATE_OFFSET = 9'h 178;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ERR_CODE_OFFSET = 9'h 17c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_STD_FAULT_STATUS_OFFSET = 9'h 180;
  parameter logic [CoreAw-1:0] FLASH_CTRL_FAULT_STATUS_OFFSET = 9'h 184;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ERR_ADDR_OFFSET = 9'h 188;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ECC_SINGLE_ERR_CNT_OFFSET = 9'h 18c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ECC_SINGLE_ERR_ADDR_0_OFFSET = 9'h 190;
  parameter logic [CoreAw-1:0] FLASH_CTRL_ECC_SINGLE_ERR_ADDR_1_OFFSET = 9'h 194;
  parameter logic [CoreAw-1:0] FLASH_CTRL_PHY_ALERT_CFG_OFFSET = 9'h 198;
  parameter logic [CoreAw-1:0] FLASH_CTRL_PHY_STATUS_OFFSET = 9'h 19c;
  parameter logic [CoreAw-1:0] FLASH_CTRL_SCRATCH_OFFSET = 9'h 1a0;
  parameter logic [CoreAw-1:0] FLASH_CTRL_FIFO_LVL_OFFSET = 9'h 1a4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_FIFO_RST_OFFSET = 9'h 1a8;
  parameter logic [CoreAw-1:0] FLASH_CTRL_CURR_FIFO_LVL_OFFSET = 9'h 1ac;

  // Reset values for hwext registers and their fields for core interface
  parameter logic [5:0] FLASH_CTRL_INTR_TEST_RESVAL = 6'h 0;
  parameter logic [0:0] FLASH_CTRL_INTR_TEST_PROG_EMPTY_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_INTR_TEST_PROG_LVL_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_INTR_TEST_RD_FULL_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_INTR_TEST_RD_LVL_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_INTR_TEST_OP_DONE_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_INTR_TEST_CORR_ERR_RESVAL = 1'h 0;
  parameter logic [4:0] FLASH_CTRL_ALERT_TEST_RESVAL = 5'h 0;
  parameter logic [0:0] FLASH_CTRL_ALERT_TEST_RECOV_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_ALERT_TEST_FATAL_STD_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_ALERT_TEST_FATAL_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_ALERT_TEST_FATAL_PRIM_FLASH_ALERT_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_ALERT_TEST_RECOV_PRIM_FLASH_ALERT_RESVAL = 1'h 0;
  parameter logic [0:0] FLASH_CTRL_CTRL_REGWEN_RESVAL = 1'h 1;
  parameter logic [0:0] FLASH_CTRL_CTRL_REGWEN_EN_RESVAL = 1'h 1;
  parameter logic [10:0] FLASH_CTRL_DEBUG_STATE_RESVAL = 11'h 0;
  parameter logic [12:0] FLASH_CTRL_CURR_FIFO_LVL_RESVAL = 13'h 0;
  parameter logic [4:0] FLASH_CTRL_CURR_FIFO_LVL_PROG_RESVAL = 5'h 0;
  parameter logic [4:0] FLASH_CTRL_CURR_FIFO_LVL_RD_RESVAL = 5'h 0;

  // Window parameters for core interface
  parameter logic [CoreAw-1:0] FLASH_CTRL_PROG_FIFO_OFFSET = 9'h 1b0;
  parameter int unsigned       FLASH_CTRL_PROG_FIFO_SIZE   = 'h 4;
  parameter logic [CoreAw-1:0] FLASH_CTRL_RD_FIFO_OFFSET = 9'h 1b4;
  parameter int unsigned       FLASH_CTRL_RD_FIFO_SIZE   = 'h 4;

  // Register index for core interface
  typedef enum int {
    FLASH_CTRL_INTR_STATE,
    FLASH_CTRL_INTR_ENABLE,
    FLASH_CTRL_INTR_TEST,
    FLASH_CTRL_ALERT_TEST,
    FLASH_CTRL_DIS,
    FLASH_CTRL_EXEC,
    FLASH_CTRL_INIT,
    FLASH_CTRL_CTRL_REGWEN,
    FLASH_CTRL_CONTROL,
    FLASH_CTRL_ADDR,
    FLASH_CTRL_PROG_TYPE_EN,
    FLASH_CTRL_ERASE_SUSPEND,
    FLASH_CTRL_REGION_CFG_REGWEN_0,
    FLASH_CTRL_REGION_CFG_REGWEN_1,
    FLASH_CTRL_REGION_CFG_REGWEN_2,
    FLASH_CTRL_REGION_CFG_REGWEN_3,
    FLASH_CTRL_REGION_CFG_REGWEN_4,
    FLASH_CTRL_REGION_CFG_REGWEN_5,
    FLASH_CTRL_REGION_CFG_REGWEN_6,
    FLASH_CTRL_REGION_CFG_REGWEN_7,
    FLASH_CTRL_MP_REGION_CFG_0,
    FLASH_CTRL_MP_REGION_CFG_1,
    FLASH_CTRL_MP_REGION_CFG_2,
    FLASH_CTRL_MP_REGION_CFG_3,
    FLASH_CTRL_MP_REGION_CFG_4,
    FLASH_CTRL_MP_REGION_CFG_5,
    FLASH_CTRL_MP_REGION_CFG_6,
    FLASH_CTRL_MP_REGION_CFG_7,
    FLASH_CTRL_MP_REGION_0,
    FLASH_CTRL_MP_REGION_1,
    FLASH_CTRL_MP_REGION_2,
    FLASH_CTRL_MP_REGION_3,
    FLASH_CTRL_MP_REGION_4,
    FLASH_CTRL_MP_REGION_5,
    FLASH_CTRL_MP_REGION_6,
    FLASH_CTRL_MP_REGION_7,
    FLASH_CTRL_DEFAULT_REGION,
    FLASH_CTRL_BANK0_INFO0_REGWEN_0,
    FLASH_CTRL_BANK0_INFO0_REGWEN_1,
    FLASH_CTRL_BANK0_INFO0_REGWEN_2,
    FLASH_CTRL_BANK0_INFO0_REGWEN_3,
    FLASH_CTRL_BANK0_INFO0_REGWEN_4,
    FLASH_CTRL_BANK0_INFO0_REGWEN_5,
    FLASH_CTRL_BANK0_INFO0_REGWEN_6,
    FLASH_CTRL_BANK0_INFO0_REGWEN_7,
    FLASH_CTRL_BANK0_INFO0_REGWEN_8,
    FLASH_CTRL_BANK0_INFO0_REGWEN_9,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_0,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_1,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_2,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_3,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_4,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_5,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_6,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_7,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_8,
    FLASH_CTRL_BANK0_INFO0_PAGE_CFG_9,
    FLASH_CTRL_BANK0_INFO1_REGWEN,
    FLASH_CTRL_BANK0_INFO1_PAGE_CFG,
    FLASH_CTRL_BANK0_INFO2_REGWEN_0,
    FLASH_CTRL_BANK0_INFO2_REGWEN_1,
    FLASH_CTRL_BANK0_INFO2_PAGE_CFG_0,
    FLASH_CTRL_BANK0_INFO2_PAGE_CFG_1,
    FLASH_CTRL_BANK1_INFO0_REGWEN_0,
    FLASH_CTRL_BANK1_INFO0_REGWEN_1,
    FLASH_CTRL_BANK1_INFO0_REGWEN_2,
    FLASH_CTRL_BANK1_INFO0_REGWEN_3,
    FLASH_CTRL_BANK1_INFO0_REGWEN_4,
    FLASH_CTRL_BANK1_INFO0_REGWEN_5,
    FLASH_CTRL_BANK1_INFO0_REGWEN_6,
    FLASH_CTRL_BANK1_INFO0_REGWEN_7,
    FLASH_CTRL_BANK1_INFO0_REGWEN_8,
    FLASH_CTRL_BANK1_INFO0_REGWEN_9,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_0,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_1,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_2,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_3,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_4,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_5,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_6,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_7,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_8,
    FLASH_CTRL_BANK1_INFO0_PAGE_CFG_9,
    FLASH_CTRL_BANK1_INFO1_REGWEN,
    FLASH_CTRL_BANK1_INFO1_PAGE_CFG,
    FLASH_CTRL_BANK1_INFO2_REGWEN_0,
    FLASH_CTRL_BANK1_INFO2_REGWEN_1,
    FLASH_CTRL_BANK1_INFO2_PAGE_CFG_0,
    FLASH_CTRL_BANK1_INFO2_PAGE_CFG_1,
    FLASH_CTRL_HW_INFO_CFG_OVERRIDE,
    FLASH_CTRL_BANK_CFG_REGWEN,
    FLASH_CTRL_MP_BANK_CFG_SHADOWED,
    FLASH_CTRL_OP_STATUS,
    FLASH_CTRL_STATUS,
    FLASH_CTRL_DEBUG_STATE,
    FLASH_CTRL_ERR_CODE,
    FLASH_CTRL_STD_FAULT_STATUS,
    FLASH_CTRL_FAULT_STATUS,
    FLASH_CTRL_ERR_ADDR,
    FLASH_CTRL_ECC_SINGLE_ERR_CNT,
    FLASH_CTRL_ECC_SINGLE_ERR_ADDR_0,
    FLASH_CTRL_ECC_SINGLE_ERR_ADDR_1,
    FLASH_CTRL_PHY_ALERT_CFG,
    FLASH_CTRL_PHY_STATUS,
    FLASH_CTRL_SCRATCH,
    FLASH_CTRL_FIFO_LVL,
    FLASH_CTRL_FIFO_RST,
    FLASH_CTRL_CURR_FIFO_LVL
  } flash_ctrl_core_id_e;

  // Register width information to check illegal writes for core interface
  parameter logic [3:0] FLASH_CTRL_CORE_PERMIT [108] = '{
    4'b 0001, // index[  0] FLASH_CTRL_INTR_STATE
    4'b 0001, // index[  1] FLASH_CTRL_INTR_ENABLE
    4'b 0001, // index[  2] FLASH_CTRL_INTR_TEST
    4'b 0001, // index[  3] FLASH_CTRL_ALERT_TEST
    4'b 0001, // index[  4] FLASH_CTRL_DIS
    4'b 1111, // index[  5] FLASH_CTRL_EXEC
    4'b 0001, // index[  6] FLASH_CTRL_INIT
    4'b 0001, // index[  7] FLASH_CTRL_CTRL_REGWEN
    4'b 1111, // index[  8] FLASH_CTRL_CONTROL
    4'b 0111, // index[  9] FLASH_CTRL_ADDR
    4'b 0001, // index[ 10] FLASH_CTRL_PROG_TYPE_EN
    4'b 0001, // index[ 11] FLASH_CTRL_ERASE_SUSPEND
    4'b 0001, // index[ 12] FLASH_CTRL_REGION_CFG_REGWEN_0
    4'b 0001, // index[ 13] FLASH_CTRL_REGION_CFG_REGWEN_1
    4'b 0001, // index[ 14] FLASH_CTRL_REGION_CFG_REGWEN_2
    4'b 0001, // index[ 15] FLASH_CTRL_REGION_CFG_REGWEN_3
    4'b 0001, // index[ 16] FLASH_CTRL_REGION_CFG_REGWEN_4
    4'b 0001, // index[ 17] FLASH_CTRL_REGION_CFG_REGWEN_5
    4'b 0001, // index[ 18] FLASH_CTRL_REGION_CFG_REGWEN_6
    4'b 0001, // index[ 19] FLASH_CTRL_REGION_CFG_REGWEN_7
    4'b 1111, // index[ 20] FLASH_CTRL_MP_REGION_CFG_0
    4'b 1111, // index[ 21] FLASH_CTRL_MP_REGION_CFG_1
    4'b 1111, // index[ 22] FLASH_CTRL_MP_REGION_CFG_2
    4'b 1111, // index[ 23] FLASH_CTRL_MP_REGION_CFG_3
    4'b 1111, // index[ 24] FLASH_CTRL_MP_REGION_CFG_4
    4'b 1111, // index[ 25] FLASH_CTRL_MP_REGION_CFG_5
    4'b 1111, // index[ 26] FLASH_CTRL_MP_REGION_CFG_6
    4'b 1111, // index[ 27] FLASH_CTRL_MP_REGION_CFG_7
    4'b 0111, // index[ 28] FLASH_CTRL_MP_REGION_0
    4'b 0111, // index[ 29] FLASH_CTRL_MP_REGION_1
    4'b 0111, // index[ 30] FLASH_CTRL_MP_REGION_2
    4'b 0111, // index[ 31] FLASH_CTRL_MP_REGION_3
    4'b 0111, // index[ 32] FLASH_CTRL_MP_REGION_4
    4'b 0111, // index[ 33] FLASH_CTRL_MP_REGION_5
    4'b 0111, // index[ 34] FLASH_CTRL_MP_REGION_6
    4'b 0111, // index[ 35] FLASH_CTRL_MP_REGION_7
    4'b 0111, // index[ 36] FLASH_CTRL_DEFAULT_REGION
    4'b 0001, // index[ 37] FLASH_CTRL_BANK0_INFO0_REGWEN_0
    4'b 0001, // index[ 38] FLASH_CTRL_BANK0_INFO0_REGWEN_1
    4'b 0001, // index[ 39] FLASH_CTRL_BANK0_INFO0_REGWEN_2
    4'b 0001, // index[ 40] FLASH_CTRL_BANK0_INFO0_REGWEN_3
    4'b 0001, // index[ 41] FLASH_CTRL_BANK0_INFO0_REGWEN_4
    4'b 0001, // index[ 42] FLASH_CTRL_BANK0_INFO0_REGWEN_5
    4'b 0001, // index[ 43] FLASH_CTRL_BANK0_INFO0_REGWEN_6
    4'b 0001, // index[ 44] FLASH_CTRL_BANK0_INFO0_REGWEN_7
    4'b 0001, // index[ 45] FLASH_CTRL_BANK0_INFO0_REGWEN_8
    4'b 0001, // index[ 46] FLASH_CTRL_BANK0_INFO0_REGWEN_9
    4'b 1111, // index[ 47] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_0
    4'b 1111, // index[ 48] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_1
    4'b 1111, // index[ 49] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_2
    4'b 1111, // index[ 50] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_3
    4'b 1111, // index[ 51] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_4
    4'b 1111, // index[ 52] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_5
    4'b 1111, // index[ 53] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_6
    4'b 1111, // index[ 54] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_7
    4'b 1111, // index[ 55] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_8
    4'b 1111, // index[ 56] FLASH_CTRL_BANK0_INFO0_PAGE_CFG_9
    4'b 0001, // index[ 57] FLASH_CTRL_BANK0_INFO1_REGWEN
    4'b 1111, // index[ 58] FLASH_CTRL_BANK0_INFO1_PAGE_CFG
    4'b 0001, // index[ 59] FLASH_CTRL_BANK0_INFO2_REGWEN_0
    4'b 0001, // index[ 60] FLASH_CTRL_BANK0_INFO2_REGWEN_1
    4'b 1111, // index[ 61] FLASH_CTRL_BANK0_INFO2_PAGE_CFG_0
    4'b 1111, // index[ 62] FLASH_CTRL_BANK0_INFO2_PAGE_CFG_1
    4'b 0001, // index[ 63] FLASH_CTRL_BANK1_INFO0_REGWEN_0
    4'b 0001, // index[ 64] FLASH_CTRL_BANK1_INFO0_REGWEN_1
    4'b 0001, // index[ 65] FLASH_CTRL_BANK1_INFO0_REGWEN_2
    4'b 0001, // index[ 66] FLASH_CTRL_BANK1_INFO0_REGWEN_3
    4'b 0001, // index[ 67] FLASH_CTRL_BANK1_INFO0_REGWEN_4
    4'b 0001, // index[ 68] FLASH_CTRL_BANK1_INFO0_REGWEN_5
    4'b 0001, // index[ 69] FLASH_CTRL_BANK1_INFO0_REGWEN_6
    4'b 0001, // index[ 70] FLASH_CTRL_BANK1_INFO0_REGWEN_7
    4'b 0001, // index[ 71] FLASH_CTRL_BANK1_INFO0_REGWEN_8
    4'b 0001, // index[ 72] FLASH_CTRL_BANK1_INFO0_REGWEN_9
    4'b 1111, // index[ 73] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_0
    4'b 1111, // index[ 74] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_1
    4'b 1111, // index[ 75] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_2
    4'b 1111, // index[ 76] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_3
    4'b 1111, // index[ 77] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_4
    4'b 1111, // index[ 78] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_5
    4'b 1111, // index[ 79] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_6
    4'b 1111, // index[ 80] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_7
    4'b 1111, // index[ 81] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_8
    4'b 1111, // index[ 82] FLASH_CTRL_BANK1_INFO0_PAGE_CFG_9
    4'b 0001, // index[ 83] FLASH_CTRL_BANK1_INFO1_REGWEN
    4'b 1111, // index[ 84] FLASH_CTRL_BANK1_INFO1_PAGE_CFG
    4'b 0001, // index[ 85] FLASH_CTRL_BANK1_INFO2_REGWEN_0
    4'b 0001, // index[ 86] FLASH_CTRL_BANK1_INFO2_REGWEN_1
    4'b 1111, // index[ 87] FLASH_CTRL_BANK1_INFO2_PAGE_CFG_0
    4'b 1111, // index[ 88] FLASH_CTRL_BANK1_INFO2_PAGE_CFG_1
    4'b 0001, // index[ 89] FLASH_CTRL_HW_INFO_CFG_OVERRIDE
    4'b 0001, // index[ 90] FLASH_CTRL_BANK_CFG_REGWEN
    4'b 0001, // index[ 91] FLASH_CTRL_MP_BANK_CFG_SHADOWED
    4'b 0001, // index[ 92] FLASH_CTRL_OP_STATUS
    4'b 0001, // index[ 93] FLASH_CTRL_STATUS
    4'b 0011, // index[ 94] FLASH_CTRL_DEBUG_STATE
    4'b 0001, // index[ 95] FLASH_CTRL_ERR_CODE
    4'b 0011, // index[ 96] FLASH_CTRL_STD_FAULT_STATUS
    4'b 0011, // index[ 97] FLASH_CTRL_FAULT_STATUS
    4'b 0111, // index[ 98] FLASH_CTRL_ERR_ADDR
    4'b 0011, // index[ 99] FLASH_CTRL_ECC_SINGLE_ERR_CNT
    4'b 0111, // index[100] FLASH_CTRL_ECC_SINGLE_ERR_ADDR_0
    4'b 0111, // index[101] FLASH_CTRL_ECC_SINGLE_ERR_ADDR_1
    4'b 0001, // index[102] FLASH_CTRL_PHY_ALERT_CFG
    4'b 0001, // index[103] FLASH_CTRL_PHY_STATUS
    4'b 1111, // index[104] FLASH_CTRL_SCRATCH
    4'b 0011, // index[105] FLASH_CTRL_FIFO_LVL
    4'b 0001, // index[106] FLASH_CTRL_FIFO_RST
    4'b 0011  // index[107] FLASH_CTRL_CURR_FIFO_LVL
  };

  ///////////////////////////////////////////////
  // Typedefs for registers for prim interface //
  ///////////////////////////////////////////////

  typedef struct packed {
    struct packed {
      logic [7:0]  q;
    } field0;
    struct packed {
      logic [4:0]  q;
    } field1;
  } flash_ctrl_reg2hw_csr1_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } field0;
    struct packed {
      logic        q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic        q;
    } field3;
    struct packed {
      logic        q;
    } field4;
    struct packed {
      logic        q;
    } field5;
    struct packed {
      logic        q;
    } field6;
    struct packed {
      logic        q;
    } field7;
  } flash_ctrl_reg2hw_csr2_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } field0;
    struct packed {
      logic [3:0]  q;
    } field1;
    struct packed {
      logic [2:0]  q;
    } field2;
    struct packed {
      logic [2:0]  q;
    } field3;
    struct packed {
      logic [2:0]  q;
    } field4;
    struct packed {
      logic [2:0]  q;
    } field5;
    struct packed {
      logic        q;
    } field6;
    struct packed {
      logic [2:0]  q;
    } field7;
    struct packed {
      logic [1:0]  q;
    } field8;
    struct packed {
      logic [1:0]  q;
    } field9;
  } flash_ctrl_reg2hw_csr3_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  q;
    } field0;
    struct packed {
      logic [2:0]  q;
    } field1;
    struct packed {
      logic [2:0]  q;
    } field2;
    struct packed {
      logic [2:0]  q;
    } field3;
  } flash_ctrl_reg2hw_csr4_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  q;
    } field0;
    struct packed {
      logic [1:0]  q;
    } field1;
    struct packed {
      logic [8:0]  q;
    } field2;
    struct packed {
      logic [4:0]  q;
    } field3;
    struct packed {
      logic [3:0]  q;
    } field4;
  } flash_ctrl_reg2hw_csr5_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  q;
    } field0;
    struct packed {
      logic [2:0]  q;
    } field1;
    struct packed {
      logic [7:0]  q;
    } field2;
    struct packed {
      logic [2:0]  q;
    } field3;
    struct packed {
      logic [1:0]  q;
    } field4;
    struct packed {
      logic [1:0]  q;
    } field5;
    struct packed {
      logic [1:0]  q;
    } field6;
    struct packed {
      logic        q;
    } field7;
    struct packed {
      logic        q;
    } field8;
  } flash_ctrl_reg2hw_csr6_reg_t;

  typedef struct packed {
    struct packed {
      logic [7:0]  q;
    } field0;
    struct packed {
      logic [8:0]  q;
    } field1;
  } flash_ctrl_reg2hw_csr7_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } flash_ctrl_reg2hw_csr8_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } flash_ctrl_reg2hw_csr9_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } flash_ctrl_reg2hw_csr10_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } flash_ctrl_reg2hw_csr11_reg_t;

  typedef struct packed {
    logic [9:0] q;
  } flash_ctrl_reg2hw_csr12_reg_t;

  typedef struct packed {
    struct packed {
      logic [19:0] q;
    } field0;
    struct packed {
      logic        q;
    } field1;
  } flash_ctrl_reg2hw_csr13_reg_t;

  typedef struct packed {
    struct packed {
      logic [7:0]  q;
    } field0;
    struct packed {
      logic        q;
    } field1;
  } flash_ctrl_reg2hw_csr14_reg_t;

  typedef struct packed {
    struct packed {
      logic [7:0]  q;
    } field0;
    struct packed {
      logic        q;
    } field1;
  } flash_ctrl_reg2hw_csr15_reg_t;

  typedef struct packed {
    struct packed {
      logic [7:0]  q;
    } field0;
    struct packed {
      logic        q;
    } field1;
  } flash_ctrl_reg2hw_csr16_reg_t;

  typedef struct packed {
    struct packed {
      logic [7:0]  q;
    } field0;
    struct packed {
      logic        q;
    } field1;
  } flash_ctrl_reg2hw_csr17_reg_t;

  typedef struct packed {
    logic        q;
  } flash_ctrl_reg2hw_csr18_reg_t;

  typedef struct packed {
    logic        q;
  } flash_ctrl_reg2hw_csr19_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } field0;
    struct packed {
      logic        q;
    } field1;
    struct packed {
      logic        q;
    } field2;
  } flash_ctrl_reg2hw_csr20_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } field0;
    struct packed {
      logic        d;
      logic        de;
    } field1;
    struct packed {
      logic        d;
      logic        de;
    } field2;
    struct packed {
      logic        d;
      logic        de;
    } field3;
    struct packed {
      logic        d;
      logic        de;
    } field4;
    struct packed {
      logic        d;
      logic        de;
    } field5;
    struct packed {
      logic        d;
      logic        de;
    } field6;
    struct packed {
      logic        d;
      logic        de;
    } field7;
  } flash_ctrl_hw2reg_csr2_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } field0;
    struct packed {
      logic        d;
      logic        de;
    } field1;
    struct packed {
      logic        d;
      logic        de;
    } field2;
  } flash_ctrl_hw2reg_csr20_reg_t;

  // Register -> HW type for prim interface
  typedef struct packed {
    flash_ctrl_reg2hw_csr1_reg_t csr1; // [325:313]
    flash_ctrl_reg2hw_csr2_reg_t csr2; // [312:305]
    flash_ctrl_reg2hw_csr3_reg_t csr3; // [304:277]
    flash_ctrl_reg2hw_csr4_reg_t csr4; // [276:265]
    flash_ctrl_reg2hw_csr5_reg_t csr5; // [264:242]
    flash_ctrl_reg2hw_csr6_reg_t csr6; // [241:217]
    flash_ctrl_reg2hw_csr7_reg_t csr7; // [216:200]
    flash_ctrl_reg2hw_csr8_reg_t csr8; // [199:168]
    flash_ctrl_reg2hw_csr9_reg_t csr9; // [167:136]
    flash_ctrl_reg2hw_csr10_reg_t csr10; // [135:104]
    flash_ctrl_reg2hw_csr11_reg_t csr11; // [103:72]
    flash_ctrl_reg2hw_csr12_reg_t csr12; // [71:62]
    flash_ctrl_reg2hw_csr13_reg_t csr13; // [61:41]
    flash_ctrl_reg2hw_csr14_reg_t csr14; // [40:32]
    flash_ctrl_reg2hw_csr15_reg_t csr15; // [31:23]
    flash_ctrl_reg2hw_csr16_reg_t csr16; // [22:14]
    flash_ctrl_reg2hw_csr17_reg_t csr17; // [13:5]
    flash_ctrl_reg2hw_csr18_reg_t csr18; // [4:4]
    flash_ctrl_reg2hw_csr19_reg_t csr19; // [3:3]
    flash_ctrl_reg2hw_csr20_reg_t csr20; // [2:0]
  } flash_ctrl_prim_reg2hw_t;

  // HW -> register type for prim interface
  typedef struct packed {
    flash_ctrl_hw2reg_csr2_reg_t csr2; // [21:6]
    flash_ctrl_hw2reg_csr20_reg_t csr20; // [5:0]
  } flash_ctrl_prim_hw2reg_t;

  // Register offsets for prim interface
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR0_REGWEN_OFFSET = 7'h 0;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR1_OFFSET = 7'h 4;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR2_OFFSET = 7'h 8;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR3_OFFSET = 7'h c;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR4_OFFSET = 7'h 10;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR5_OFFSET = 7'h 14;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR6_OFFSET = 7'h 18;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR7_OFFSET = 7'h 1c;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR8_OFFSET = 7'h 20;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR9_OFFSET = 7'h 24;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR10_OFFSET = 7'h 28;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR11_OFFSET = 7'h 2c;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR12_OFFSET = 7'h 30;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR13_OFFSET = 7'h 34;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR14_OFFSET = 7'h 38;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR15_OFFSET = 7'h 3c;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR16_OFFSET = 7'h 40;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR17_OFFSET = 7'h 44;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR18_OFFSET = 7'h 48;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR19_OFFSET = 7'h 4c;
  parameter logic [PrimAw-1:0] FLASH_CTRL_CSR20_OFFSET = 7'h 50;

  // Register index for prim interface
  typedef enum int {
    FLASH_CTRL_CSR0_REGWEN,
    FLASH_CTRL_CSR1,
    FLASH_CTRL_CSR2,
    FLASH_CTRL_CSR3,
    FLASH_CTRL_CSR4,
    FLASH_CTRL_CSR5,
    FLASH_CTRL_CSR6,
    FLASH_CTRL_CSR7,
    FLASH_CTRL_CSR8,
    FLASH_CTRL_CSR9,
    FLASH_CTRL_CSR10,
    FLASH_CTRL_CSR11,
    FLASH_CTRL_CSR12,
    FLASH_CTRL_CSR13,
    FLASH_CTRL_CSR14,
    FLASH_CTRL_CSR15,
    FLASH_CTRL_CSR16,
    FLASH_CTRL_CSR17,
    FLASH_CTRL_CSR18,
    FLASH_CTRL_CSR19,
    FLASH_CTRL_CSR20
  } flash_ctrl_prim_id_e;

  // Register width information to check illegal writes for prim interface
  parameter logic [3:0] FLASH_CTRL_PRIM_PERMIT [21] = '{
    4'b 0001, // index[ 0] FLASH_CTRL_CSR0_REGWEN
    4'b 0011, // index[ 1] FLASH_CTRL_CSR1
    4'b 0001, // index[ 2] FLASH_CTRL_CSR2
    4'b 1111, // index[ 3] FLASH_CTRL_CSR3
    4'b 0011, // index[ 4] FLASH_CTRL_CSR4
    4'b 0111, // index[ 5] FLASH_CTRL_CSR5
    4'b 1111, // index[ 6] FLASH_CTRL_CSR6
    4'b 0111, // index[ 7] FLASH_CTRL_CSR7
    4'b 1111, // index[ 8] FLASH_CTRL_CSR8
    4'b 1111, // index[ 9] FLASH_CTRL_CSR9
    4'b 1111, // index[10] FLASH_CTRL_CSR10
    4'b 1111, // index[11] FLASH_CTRL_CSR11
    4'b 0011, // index[12] FLASH_CTRL_CSR12
    4'b 0111, // index[13] FLASH_CTRL_CSR13
    4'b 0011, // index[14] FLASH_CTRL_CSR14
    4'b 0011, // index[15] FLASH_CTRL_CSR15
    4'b 0011, // index[16] FLASH_CTRL_CSR16
    4'b 0011, // index[17] FLASH_CTRL_CSR17
    4'b 0001, // index[18] FLASH_CTRL_CSR18
    4'b 0001, // index[19] FLASH_CTRL_CSR19
    4'b 0001  // index[20] FLASH_CTRL_CSR20
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package jtag_pkg;

  typedef struct packed {
    logic tck;
    logic tms;
    logic trst_n;
    logic tdi;
  } jtag_req_t;

  parameter jtag_req_t JTAG_REQ_DEFAULT = '0;

  typedef struct packed {
    logic tdo;
    logic tdo_oe;
  } jtag_rsp_t;

  parameter jtag_rsp_t JTAG_RSP_DEFAULT = '0;

endpackage : jtag_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package otp_ctrl_reg_pkg;

  // Param list
  parameter int NumSramKeyReqSlots = 3;
  parameter int OtpByteAddrWidth = 11;
  parameter int NumErrorEntries = 10;
  parameter int NumDaiWords = 2;
  parameter int NumDigestWords = 2;
  parameter int NumSwCfgWindowWords = 512;
  parameter int NumPart = 8;
  parameter int VendorTestOffset = 0;
  parameter int VendorTestSize = 64;
  parameter int ScratchOffset = 0;
  parameter int ScratchSize = 56;
  parameter int VendorTestDigestOffset = 56;
  parameter int VendorTestDigestSize = 8;
  parameter int CreatorSwCfgOffset = 64;
  parameter int CreatorSwCfgSize = 800;
  parameter int CreatorSwCfgAstCfgOffset = 64;
  parameter int CreatorSwCfgAstCfgSize = 156;
  parameter int CreatorSwCfgAstInitEnOffset = 220;
  parameter int CreatorSwCfgAstInitEnSize = 4;
  parameter int CreatorSwCfgRomExtSkuOffset = 224;
  parameter int CreatorSwCfgRomExtSkuSize = 4;
  parameter int CreatorSwCfgSigverifyRsaModExpIbexEnOffset = 228;
  parameter int CreatorSwCfgSigverifyRsaModExpIbexEnSize = 4;
  parameter int CreatorSwCfgSigverifyRsaKeyEnOffset = 232;
  parameter int CreatorSwCfgSigverifyRsaKeyEnSize = 8;
  parameter int CreatorSwCfgSigverifySpxEnOffset = 240;
  parameter int CreatorSwCfgSigverifySpxEnSize = 4;
  parameter int CreatorSwCfgSigverifySpxKeyEnOffset = 244;
  parameter int CreatorSwCfgSigverifySpxKeyEnSize = 8;
  parameter int CreatorSwCfgFlashDataDefaultCfgOffset = 252;
  parameter int CreatorSwCfgFlashDataDefaultCfgSize = 4;
  parameter int CreatorSwCfgFlashInfoBootDataCfgOffset = 256;
  parameter int CreatorSwCfgFlashInfoBootDataCfgSize = 4;
  parameter int CreatorSwCfgFlashHwInfoCfgOverrideOffset = 260;
  parameter int CreatorSwCfgFlashHwInfoCfgOverrideSize = 4;
  parameter int CreatorSwCfgRngEnOffset = 264;
  parameter int CreatorSwCfgRngEnSize = 4;
  parameter int CreatorSwCfgJitterEnOffset = 268;
  parameter int CreatorSwCfgJitterEnSize = 4;
  parameter int CreatorSwCfgRetRamResetMaskOffset = 272;
  parameter int CreatorSwCfgRetRamResetMaskSize = 4;
  parameter int CreatorSwCfgManufStateOffset = 276;
  parameter int CreatorSwCfgManufStateSize = 4;
  parameter int CreatorSwCfgRomExecEnOffset = 280;
  parameter int CreatorSwCfgRomExecEnSize = 4;
  parameter int CreatorSwCfgCpuctrlOffset = 284;
  parameter int CreatorSwCfgCpuctrlSize = 4;
  parameter int CreatorSwCfgMinSecVerRomExtOffset = 288;
  parameter int CreatorSwCfgMinSecVerRomExtSize = 4;
  parameter int CreatorSwCfgMinSecVerBl0Offset = 292;
  parameter int CreatorSwCfgMinSecVerBl0Size = 4;
  parameter int CreatorSwCfgDefaultBootDataInProdEnOffset = 296;
  parameter int CreatorSwCfgDefaultBootDataInProdEnSize = 4;
  parameter int CreatorSwCfgRmaSpinEnOffset = 300;
  parameter int CreatorSwCfgRmaSpinEnSize = 4;
  parameter int CreatorSwCfgRmaSpinCyclesOffset = 304;
  parameter int CreatorSwCfgRmaSpinCyclesSize = 4;
  parameter int CreatorSwCfgRngRepcntThresholdsOffset = 308;
  parameter int CreatorSwCfgRngRepcntThresholdsSize = 4;
  parameter int CreatorSwCfgRngRepcntsThresholdsOffset = 312;
  parameter int CreatorSwCfgRngRepcntsThresholdsSize = 4;
  parameter int CreatorSwCfgRngAdaptpHiThresholdsOffset = 316;
  parameter int CreatorSwCfgRngAdaptpHiThresholdsSize = 4;
  parameter int CreatorSwCfgRngAdaptpLoThresholdsOffset = 320;
  parameter int CreatorSwCfgRngAdaptpLoThresholdsSize = 4;
  parameter int CreatorSwCfgRngBucketThresholdsOffset = 324;
  parameter int CreatorSwCfgRngBucketThresholdsSize = 4;
  parameter int CreatorSwCfgRngMarkovHiThresholdsOffset = 328;
  parameter int CreatorSwCfgRngMarkovHiThresholdsSize = 4;
  parameter int CreatorSwCfgRngMarkovLoThresholdsOffset = 332;
  parameter int CreatorSwCfgRngMarkovLoThresholdsSize = 4;
  parameter int CreatorSwCfgRngExthtHiThresholdsOffset = 336;
  parameter int CreatorSwCfgRngExthtHiThresholdsSize = 4;
  parameter int CreatorSwCfgRngExthtLoThresholdsOffset = 340;
  parameter int CreatorSwCfgRngExthtLoThresholdsSize = 4;
  parameter int CreatorSwCfgRngAlertThresholdOffset = 344;
  parameter int CreatorSwCfgRngAlertThresholdSize = 4;
  parameter int CreatorSwCfgRngHealthConfigDigestOffset = 348;
  parameter int CreatorSwCfgRngHealthConfigDigestSize = 4;
  parameter int CreatorSwCfgDigestOffset = 856;
  parameter int CreatorSwCfgDigestSize = 8;
  parameter int OwnerSwCfgOffset = 864;
  parameter int OwnerSwCfgSize = 800;
  parameter int OwnerSwCfgRomErrorReportingOffset = 864;
  parameter int OwnerSwCfgRomErrorReportingSize = 4;
  parameter int OwnerSwCfgRomBootstrapDisOffset = 868;
  parameter int OwnerSwCfgRomBootstrapDisSize = 4;
  parameter int OwnerSwCfgRomAlertClassEnOffset = 872;
  parameter int OwnerSwCfgRomAlertClassEnSize = 4;
  parameter int OwnerSwCfgRomAlertEscalationOffset = 876;
  parameter int OwnerSwCfgRomAlertEscalationSize = 4;
  parameter int OwnerSwCfgRomAlertClassificationOffset = 880;
  parameter int OwnerSwCfgRomAlertClassificationSize = 320;
  parameter int OwnerSwCfgRomLocalAlertClassificationOffset = 1200;
  parameter int OwnerSwCfgRomLocalAlertClassificationSize = 64;
  parameter int OwnerSwCfgRomAlertAccumThreshOffset = 1264;
  parameter int OwnerSwCfgRomAlertAccumThreshSize = 16;
  parameter int OwnerSwCfgRomAlertTimeoutCyclesOffset = 1280;
  parameter int OwnerSwCfgRomAlertTimeoutCyclesSize = 16;
  parameter int OwnerSwCfgRomAlertPhaseCyclesOffset = 1296;
  parameter int OwnerSwCfgRomAlertPhaseCyclesSize = 64;
  parameter int OwnerSwCfgRomAlertDigestProdOffset = 1360;
  parameter int OwnerSwCfgRomAlertDigestProdSize = 4;
  parameter int OwnerSwCfgRomAlertDigestProdEndOffset = 1364;
  parameter int OwnerSwCfgRomAlertDigestProdEndSize = 4;
  parameter int OwnerSwCfgRomAlertDigestDevOffset = 1368;
  parameter int OwnerSwCfgRomAlertDigestDevSize = 4;
  parameter int OwnerSwCfgRomAlertDigestRmaOffset = 1372;
  parameter int OwnerSwCfgRomAlertDigestRmaSize = 4;
  parameter int OwnerSwCfgRomWatchdogBiteThresholdCyclesOffset = 1376;
  parameter int OwnerSwCfgRomWatchdogBiteThresholdCyclesSize = 4;
  parameter int OwnerSwCfgRomKeymgrRomExtMeasEnOffset = 1380;
  parameter int OwnerSwCfgRomKeymgrRomExtMeasEnSize = 4;
  parameter int OwnerSwCfgManufStateOffset = 1384;
  parameter int OwnerSwCfgManufStateSize = 4;
  parameter int OwnerSwCfgDigestOffset = 1656;
  parameter int OwnerSwCfgDigestSize = 8;
  parameter int HwCfgOffset = 1664;
  parameter int HwCfgSize = 80;
  parameter int DeviceIdOffset = 1664;
  parameter int DeviceIdSize = 32;
  parameter int ManufStateOffset = 1696;
  parameter int ManufStateSize = 32;
  parameter int EnSramIfetchOffset = 1728;
  parameter int EnSramIfetchSize = 1;
  parameter int EnCsrngSwAppReadOffset = 1729;
  parameter int EnCsrngSwAppReadSize = 1;
  parameter int EnEntropySrcFwReadOffset = 1730;
  parameter int EnEntropySrcFwReadSize = 1;
  parameter int EnEntropySrcFwOverOffset = 1731;
  parameter int EnEntropySrcFwOverSize = 1;
  parameter int HwCfgDigestOffset = 1736;
  parameter int HwCfgDigestSize = 8;
  parameter int Secret0Offset = 1744;
  parameter int Secret0Size = 40;
  parameter int TestUnlockTokenOffset = 1744;
  parameter int TestUnlockTokenSize = 16;
  parameter int TestExitTokenOffset = 1760;
  parameter int TestExitTokenSize = 16;
  parameter int Secret0DigestOffset = 1776;
  parameter int Secret0DigestSize = 8;
  parameter int Secret1Offset = 1784;
  parameter int Secret1Size = 88;
  parameter int FlashAddrKeySeedOffset = 1784;
  parameter int FlashAddrKeySeedSize = 32;
  parameter int FlashDataKeySeedOffset = 1816;
  parameter int FlashDataKeySeedSize = 32;
  parameter int SramDataKeySeedOffset = 1848;
  parameter int SramDataKeySeedSize = 16;
  parameter int Secret1DigestOffset = 1864;
  parameter int Secret1DigestSize = 8;
  parameter int Secret2Offset = 1872;
  parameter int Secret2Size = 88;
  parameter int RmaTokenOffset = 1872;
  parameter int RmaTokenSize = 16;
  parameter int CreatorRootKeyShare0Offset = 1888;
  parameter int CreatorRootKeyShare0Size = 32;
  parameter int CreatorRootKeyShare1Offset = 1920;
  parameter int CreatorRootKeyShare1Size = 32;
  parameter int Secret2DigestOffset = 1952;
  parameter int Secret2DigestSize = 8;
  parameter int LifeCycleOffset = 1960;
  parameter int LifeCycleSize = 88;
  parameter int LcTransitionCntOffset = 1960;
  parameter int LcTransitionCntSize = 48;
  parameter int LcStateOffset = 2008;
  parameter int LcStateSize = 40;
  parameter int NumAlerts = 5;

  // Address widths within the block
  parameter int CoreAw = 13;
  parameter int PrimAw = 5;

  ///////////////////////////////////////////////
  // Typedefs for registers for core interface //
  ///////////////////////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } otp_operation_done;
    struct packed {
      logic        q;
    } otp_error;
  } otp_ctrl_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } otp_operation_done;
    struct packed {
      logic        q;
    } otp_error;
  } otp_ctrl_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } otp_operation_done;
    struct packed {
      logic        q;
      logic        qe;
    } otp_error;
  } otp_ctrl_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } fatal_macro_error;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_check_error;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_bus_integ_error;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_prim_otp_alert;
    struct packed {
      logic        q;
      logic        qe;
    } recov_prim_otp_alert;
  } otp_ctrl_reg2hw_alert_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } rd;
    struct packed {
      logic        q;
      logic        qe;
    } wr;
    struct packed {
      logic        q;
      logic        qe;
    } digest;
  } otp_ctrl_reg2hw_direct_access_cmd_reg_t;

  typedef struct packed {
    logic [10:0] q;
  } otp_ctrl_reg2hw_direct_access_address_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } otp_ctrl_reg2hw_direct_access_wdata_mreg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } integrity;
    struct packed {
      logic        q;
      logic        qe;
    } consistency;
  } otp_ctrl_reg2hw_check_trigger_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } otp_ctrl_reg2hw_check_timeout_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } otp_ctrl_reg2hw_integrity_check_period_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } otp_ctrl_reg2hw_consistency_check_period_reg_t;

  typedef struct packed {
    logic        q;
  } otp_ctrl_reg2hw_vendor_test_read_lock_reg_t;

  typedef struct packed {
    logic        q;
  } otp_ctrl_reg2hw_creator_sw_cfg_read_lock_reg_t;

  typedef struct packed {
    logic        q;
  } otp_ctrl_reg2hw_owner_sw_cfg_read_lock_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } otp_operation_done;
    struct packed {
      logic        d;
      logic        de;
    } otp_error;
  } otp_ctrl_hw2reg_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } vendor_test_error;
    struct packed {
      logic        d;
    } creator_sw_cfg_error;
    struct packed {
      logic        d;
    } owner_sw_cfg_error;
    struct packed {
      logic        d;
    } hw_cfg_error;
    struct packed {
      logic        d;
    } secret0_error;
    struct packed {
      logic        d;
    } secret1_error;
    struct packed {
      logic        d;
    } secret2_error;
    struct packed {
      logic        d;
    } life_cycle_error;
    struct packed {
      logic        d;
    } dai_error;
    struct packed {
      logic        d;
    } lci_error;
    struct packed {
      logic        d;
    } timeout_error;
    struct packed {
      logic        d;
    } lfsr_fsm_error;
    struct packed {
      logic        d;
    } scrambling_fsm_error;
    struct packed {
      logic        d;
    } key_deriv_fsm_error;
    struct packed {
      logic        d;
    } bus_integ_error;
    struct packed {
      logic        d;
    } dai_idle;
    struct packed {
      logic        d;
    } check_pending;
  } otp_ctrl_hw2reg_status_reg_t;

  typedef struct packed {
    logic [2:0]  d;
  } otp_ctrl_hw2reg_err_code_mreg_t;

  typedef struct packed {
    logic        d;
  } otp_ctrl_hw2reg_direct_access_regwen_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_direct_access_rdata_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_vendor_test_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_creator_sw_cfg_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_owner_sw_cfg_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_hw_cfg_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_secret0_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_secret1_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } otp_ctrl_hw2reg_secret2_digest_mreg_t;

  // Register -> HW type for core interface
  typedef struct packed {
    otp_ctrl_reg2hw_intr_state_reg_t intr_state; // [201:200]
    otp_ctrl_reg2hw_intr_enable_reg_t intr_enable; // [199:198]
    otp_ctrl_reg2hw_intr_test_reg_t intr_test; // [197:194]
    otp_ctrl_reg2hw_alert_test_reg_t alert_test; // [193:184]
    otp_ctrl_reg2hw_direct_access_cmd_reg_t direct_access_cmd; // [183:178]
    otp_ctrl_reg2hw_direct_access_address_reg_t direct_access_address; // [177:167]
    otp_ctrl_reg2hw_direct_access_wdata_mreg_t [1:0] direct_access_wdata; // [166:103]
    otp_ctrl_reg2hw_check_trigger_reg_t check_trigger; // [102:99]
    otp_ctrl_reg2hw_check_timeout_reg_t check_timeout; // [98:67]
    otp_ctrl_reg2hw_integrity_check_period_reg_t integrity_check_period; // [66:35]
    otp_ctrl_reg2hw_consistency_check_period_reg_t consistency_check_period; // [34:3]
    otp_ctrl_reg2hw_vendor_test_read_lock_reg_t vendor_test_read_lock; // [2:2]
    otp_ctrl_reg2hw_creator_sw_cfg_read_lock_reg_t creator_sw_cfg_read_lock; // [1:1]
    otp_ctrl_reg2hw_owner_sw_cfg_read_lock_reg_t owner_sw_cfg_read_lock; // [0:0]
  } otp_ctrl_core_reg2hw_t;

  // HW -> register type for core interface
  typedef struct packed {
    otp_ctrl_hw2reg_intr_state_reg_t intr_state; // [563:560]
    otp_ctrl_hw2reg_status_reg_t status; // [559:543]
    otp_ctrl_hw2reg_err_code_mreg_t [9:0] err_code; // [542:513]
    otp_ctrl_hw2reg_direct_access_regwen_reg_t direct_access_regwen; // [512:512]
    otp_ctrl_hw2reg_direct_access_rdata_mreg_t [1:0] direct_access_rdata; // [511:448]
    otp_ctrl_hw2reg_vendor_test_digest_mreg_t [1:0] vendor_test_digest; // [447:384]
    otp_ctrl_hw2reg_creator_sw_cfg_digest_mreg_t [1:0] creator_sw_cfg_digest; // [383:320]
    otp_ctrl_hw2reg_owner_sw_cfg_digest_mreg_t [1:0] owner_sw_cfg_digest; // [319:256]
    otp_ctrl_hw2reg_hw_cfg_digest_mreg_t [1:0] hw_cfg_digest; // [255:192]
    otp_ctrl_hw2reg_secret0_digest_mreg_t [1:0] secret0_digest; // [191:128]
    otp_ctrl_hw2reg_secret1_digest_mreg_t [1:0] secret1_digest; // [127:64]
    otp_ctrl_hw2reg_secret2_digest_mreg_t [1:0] secret2_digest; // [63:0]
  } otp_ctrl_core_hw2reg_t;

  // Register offsets for core interface
  parameter logic [CoreAw-1:0] OTP_CTRL_INTR_STATE_OFFSET = 13'h 0;
  parameter logic [CoreAw-1:0] OTP_CTRL_INTR_ENABLE_OFFSET = 13'h 4;
  parameter logic [CoreAw-1:0] OTP_CTRL_INTR_TEST_OFFSET = 13'h 8;
  parameter logic [CoreAw-1:0] OTP_CTRL_ALERT_TEST_OFFSET = 13'h c;
  parameter logic [CoreAw-1:0] OTP_CTRL_STATUS_OFFSET = 13'h 10;
  parameter logic [CoreAw-1:0] OTP_CTRL_ERR_CODE_OFFSET = 13'h 14;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_REGWEN_OFFSET = 13'h 18;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_CMD_OFFSET = 13'h 1c;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_ADDRESS_OFFSET = 13'h 20;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_WDATA_0_OFFSET = 13'h 24;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_WDATA_1_OFFSET = 13'h 28;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_RDATA_0_OFFSET = 13'h 2c;
  parameter logic [CoreAw-1:0] OTP_CTRL_DIRECT_ACCESS_RDATA_1_OFFSET = 13'h 30;
  parameter logic [CoreAw-1:0] OTP_CTRL_CHECK_TRIGGER_REGWEN_OFFSET = 13'h 34;
  parameter logic [CoreAw-1:0] OTP_CTRL_CHECK_TRIGGER_OFFSET = 13'h 38;
  parameter logic [CoreAw-1:0] OTP_CTRL_CHECK_REGWEN_OFFSET = 13'h 3c;
  parameter logic [CoreAw-1:0] OTP_CTRL_CHECK_TIMEOUT_OFFSET = 13'h 40;
  parameter logic [CoreAw-1:0] OTP_CTRL_INTEGRITY_CHECK_PERIOD_OFFSET = 13'h 44;
  parameter logic [CoreAw-1:0] OTP_CTRL_CONSISTENCY_CHECK_PERIOD_OFFSET = 13'h 48;
  parameter logic [CoreAw-1:0] OTP_CTRL_VENDOR_TEST_READ_LOCK_OFFSET = 13'h 4c;
  parameter logic [CoreAw-1:0] OTP_CTRL_CREATOR_SW_CFG_READ_LOCK_OFFSET = 13'h 50;
  parameter logic [CoreAw-1:0] OTP_CTRL_OWNER_SW_CFG_READ_LOCK_OFFSET = 13'h 54;
  parameter logic [CoreAw-1:0] OTP_CTRL_VENDOR_TEST_DIGEST_0_OFFSET = 13'h 58;
  parameter logic [CoreAw-1:0] OTP_CTRL_VENDOR_TEST_DIGEST_1_OFFSET = 13'h 5c;
  parameter logic [CoreAw-1:0] OTP_CTRL_CREATOR_SW_CFG_DIGEST_0_OFFSET = 13'h 60;
  parameter logic [CoreAw-1:0] OTP_CTRL_CREATOR_SW_CFG_DIGEST_1_OFFSET = 13'h 64;
  parameter logic [CoreAw-1:0] OTP_CTRL_OWNER_SW_CFG_DIGEST_0_OFFSET = 13'h 68;
  parameter logic [CoreAw-1:0] OTP_CTRL_OWNER_SW_CFG_DIGEST_1_OFFSET = 13'h 6c;
  parameter logic [CoreAw-1:0] OTP_CTRL_HW_CFG_DIGEST_0_OFFSET = 13'h 70;
  parameter logic [CoreAw-1:0] OTP_CTRL_HW_CFG_DIGEST_1_OFFSET = 13'h 74;
  parameter logic [CoreAw-1:0] OTP_CTRL_SECRET0_DIGEST_0_OFFSET = 13'h 78;
  parameter logic [CoreAw-1:0] OTP_CTRL_SECRET0_DIGEST_1_OFFSET = 13'h 7c;
  parameter logic [CoreAw-1:0] OTP_CTRL_SECRET1_DIGEST_0_OFFSET = 13'h 80;
  parameter logic [CoreAw-1:0] OTP_CTRL_SECRET1_DIGEST_1_OFFSET = 13'h 84;
  parameter logic [CoreAw-1:0] OTP_CTRL_SECRET2_DIGEST_0_OFFSET = 13'h 88;
  parameter logic [CoreAw-1:0] OTP_CTRL_SECRET2_DIGEST_1_OFFSET = 13'h 8c;

  // Reset values for hwext registers and their fields for core interface
  parameter logic [1:0] OTP_CTRL_INTR_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] OTP_CTRL_INTR_TEST_OTP_OPERATION_DONE_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_INTR_TEST_OTP_ERROR_RESVAL = 1'h 0;
  parameter logic [4:0] OTP_CTRL_ALERT_TEST_RESVAL = 5'h 0;
  parameter logic [0:0] OTP_CTRL_ALERT_TEST_FATAL_MACRO_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_ALERT_TEST_FATAL_CHECK_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_ALERT_TEST_FATAL_BUS_INTEG_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_ALERT_TEST_FATAL_PRIM_OTP_ALERT_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_ALERT_TEST_RECOV_PRIM_OTP_ALERT_RESVAL = 1'h 0;
  parameter logic [16:0] OTP_CTRL_STATUS_RESVAL = 17'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_VENDOR_TEST_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_CREATOR_SW_CFG_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_OWNER_SW_CFG_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_HW_CFG_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_SECRET0_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_SECRET1_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_SECRET2_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_LIFE_CYCLE_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_DAI_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_LCI_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_TIMEOUT_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_LFSR_FSM_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_SCRAMBLING_FSM_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_KEY_DERIV_FSM_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_BUS_INTEG_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_DAI_IDLE_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_STATUS_CHECK_PENDING_RESVAL = 1'h 0;
  parameter logic [29:0] OTP_CTRL_ERR_CODE_RESVAL = 30'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_0_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_1_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_2_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_3_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_4_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_5_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_6_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_7_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_8_RESVAL = 3'h 0;
  parameter logic [2:0] OTP_CTRL_ERR_CODE_ERR_CODE_9_RESVAL = 3'h 0;
  parameter logic [0:0] OTP_CTRL_DIRECT_ACCESS_REGWEN_RESVAL = 1'h 1;
  parameter logic [0:0] OTP_CTRL_DIRECT_ACCESS_REGWEN_DIRECT_ACCESS_REGWEN_RESVAL = 1'h 1;
  parameter logic [2:0] OTP_CTRL_DIRECT_ACCESS_CMD_RESVAL = 3'h 0;
  parameter logic [0:0] OTP_CTRL_DIRECT_ACCESS_CMD_RD_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_DIRECT_ACCESS_CMD_WR_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_DIRECT_ACCESS_CMD_DIGEST_RESVAL = 1'h 0;
  parameter logic [31:0] OTP_CTRL_DIRECT_ACCESS_RDATA_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_DIRECT_ACCESS_RDATA_0_DIRECT_ACCESS_RDATA_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_DIRECT_ACCESS_RDATA_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_DIRECT_ACCESS_RDATA_1_DIRECT_ACCESS_RDATA_1_RESVAL = 32'h 0;
  parameter logic [1:0] OTP_CTRL_CHECK_TRIGGER_RESVAL = 2'h 0;
  parameter logic [0:0] OTP_CTRL_CHECK_TRIGGER_INTEGRITY_RESVAL = 1'h 0;
  parameter logic [0:0] OTP_CTRL_CHECK_TRIGGER_CONSISTENCY_RESVAL = 1'h 0;
  parameter logic [31:0] OTP_CTRL_VENDOR_TEST_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_VENDOR_TEST_DIGEST_0_VENDOR_TEST_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_VENDOR_TEST_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_VENDOR_TEST_DIGEST_1_VENDOR_TEST_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_CREATOR_SW_CFG_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_CREATOR_SW_CFG_DIGEST_0_CREATOR_SW_CFG_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_CREATOR_SW_CFG_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_CREATOR_SW_CFG_DIGEST_1_CREATOR_SW_CFG_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_OWNER_SW_CFG_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_OWNER_SW_CFG_DIGEST_0_OWNER_SW_CFG_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_OWNER_SW_CFG_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_OWNER_SW_CFG_DIGEST_1_OWNER_SW_CFG_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_HW_CFG_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_HW_CFG_DIGEST_0_HW_CFG_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_HW_CFG_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_HW_CFG_DIGEST_1_HW_CFG_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET0_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET0_DIGEST_0_SECRET0_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET0_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET0_DIGEST_1_SECRET0_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET1_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET1_DIGEST_0_SECRET1_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET1_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET1_DIGEST_1_SECRET1_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET2_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET2_DIGEST_0_SECRET2_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET2_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] OTP_CTRL_SECRET2_DIGEST_1_SECRET2_DIGEST_1_RESVAL = 32'h 0;

  // Window parameters for core interface
  parameter logic [CoreAw-1:0] OTP_CTRL_SW_CFG_WINDOW_OFFSET = 13'h 1000;
  parameter int unsigned       OTP_CTRL_SW_CFG_WINDOW_SIZE   = 'h 800;

  // Register index for core interface
  typedef enum int {
    OTP_CTRL_INTR_STATE,
    OTP_CTRL_INTR_ENABLE,
    OTP_CTRL_INTR_TEST,
    OTP_CTRL_ALERT_TEST,
    OTP_CTRL_STATUS,
    OTP_CTRL_ERR_CODE,
    OTP_CTRL_DIRECT_ACCESS_REGWEN,
    OTP_CTRL_DIRECT_ACCESS_CMD,
    OTP_CTRL_DIRECT_ACCESS_ADDRESS,
    OTP_CTRL_DIRECT_ACCESS_WDATA_0,
    OTP_CTRL_DIRECT_ACCESS_WDATA_1,
    OTP_CTRL_DIRECT_ACCESS_RDATA_0,
    OTP_CTRL_DIRECT_ACCESS_RDATA_1,
    OTP_CTRL_CHECK_TRIGGER_REGWEN,
    OTP_CTRL_CHECK_TRIGGER,
    OTP_CTRL_CHECK_REGWEN,
    OTP_CTRL_CHECK_TIMEOUT,
    OTP_CTRL_INTEGRITY_CHECK_PERIOD,
    OTP_CTRL_CONSISTENCY_CHECK_PERIOD,
    OTP_CTRL_VENDOR_TEST_READ_LOCK,
    OTP_CTRL_CREATOR_SW_CFG_READ_LOCK,
    OTP_CTRL_OWNER_SW_CFG_READ_LOCK,
    OTP_CTRL_VENDOR_TEST_DIGEST_0,
    OTP_CTRL_VENDOR_TEST_DIGEST_1,
    OTP_CTRL_CREATOR_SW_CFG_DIGEST_0,
    OTP_CTRL_CREATOR_SW_CFG_DIGEST_1,
    OTP_CTRL_OWNER_SW_CFG_DIGEST_0,
    OTP_CTRL_OWNER_SW_CFG_DIGEST_1,
    OTP_CTRL_HW_CFG_DIGEST_0,
    OTP_CTRL_HW_CFG_DIGEST_1,
    OTP_CTRL_SECRET0_DIGEST_0,
    OTP_CTRL_SECRET0_DIGEST_1,
    OTP_CTRL_SECRET1_DIGEST_0,
    OTP_CTRL_SECRET1_DIGEST_1,
    OTP_CTRL_SECRET2_DIGEST_0,
    OTP_CTRL_SECRET2_DIGEST_1
  } otp_ctrl_core_id_e;

  // Register width information to check illegal writes for core interface
  parameter logic [3:0] OTP_CTRL_CORE_PERMIT [36] = '{
    4'b 0001, // index[ 0] OTP_CTRL_INTR_STATE
    4'b 0001, // index[ 1] OTP_CTRL_INTR_ENABLE
    4'b 0001, // index[ 2] OTP_CTRL_INTR_TEST
    4'b 0001, // index[ 3] OTP_CTRL_ALERT_TEST
    4'b 0111, // index[ 4] OTP_CTRL_STATUS
    4'b 1111, // index[ 5] OTP_CTRL_ERR_CODE
    4'b 0001, // index[ 6] OTP_CTRL_DIRECT_ACCESS_REGWEN
    4'b 0001, // index[ 7] OTP_CTRL_DIRECT_ACCESS_CMD
    4'b 0011, // index[ 8] OTP_CTRL_DIRECT_ACCESS_ADDRESS
    4'b 1111, // index[ 9] OTP_CTRL_DIRECT_ACCESS_WDATA_0
    4'b 1111, // index[10] OTP_CTRL_DIRECT_ACCESS_WDATA_1
    4'b 1111, // index[11] OTP_CTRL_DIRECT_ACCESS_RDATA_0
    4'b 1111, // index[12] OTP_CTRL_DIRECT_ACCESS_RDATA_1
    4'b 0001, // index[13] OTP_CTRL_CHECK_TRIGGER_REGWEN
    4'b 0001, // index[14] OTP_CTRL_CHECK_TRIGGER
    4'b 0001, // index[15] OTP_CTRL_CHECK_REGWEN
    4'b 1111, // index[16] OTP_CTRL_CHECK_TIMEOUT
    4'b 1111, // index[17] OTP_CTRL_INTEGRITY_CHECK_PERIOD
    4'b 1111, // index[18] OTP_CTRL_CONSISTENCY_CHECK_PERIOD
    4'b 0001, // index[19] OTP_CTRL_VENDOR_TEST_READ_LOCK
    4'b 0001, // index[20] OTP_CTRL_CREATOR_SW_CFG_READ_LOCK
    4'b 0001, // index[21] OTP_CTRL_OWNER_SW_CFG_READ_LOCK
    4'b 1111, // index[22] OTP_CTRL_VENDOR_TEST_DIGEST_0
    4'b 1111, // index[23] OTP_CTRL_VENDOR_TEST_DIGEST_1
    4'b 1111, // index[24] OTP_CTRL_CREATOR_SW_CFG_DIGEST_0
    4'b 1111, // index[25] OTP_CTRL_CREATOR_SW_CFG_DIGEST_1
    4'b 1111, // index[26] OTP_CTRL_OWNER_SW_CFG_DIGEST_0
    4'b 1111, // index[27] OTP_CTRL_OWNER_SW_CFG_DIGEST_1
    4'b 1111, // index[28] OTP_CTRL_HW_CFG_DIGEST_0
    4'b 1111, // index[29] OTP_CTRL_HW_CFG_DIGEST_1
    4'b 1111, // index[30] OTP_CTRL_SECRET0_DIGEST_0
    4'b 1111, // index[31] OTP_CTRL_SECRET0_DIGEST_1
    4'b 1111, // index[32] OTP_CTRL_SECRET1_DIGEST_0
    4'b 1111, // index[33] OTP_CTRL_SECRET1_DIGEST_1
    4'b 1111, // index[34] OTP_CTRL_SECRET2_DIGEST_0
    4'b 1111  // index[35] OTP_CTRL_SECRET2_DIGEST_1
  };

  ///////////////////////////////////////////////
  // Typedefs for registers for prim interface //
  ///////////////////////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } field0;
    struct packed {
      logic        q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic [9:0] q;
    } field3;
    struct packed {
      logic [10:0] q;
    } field4;
  } otp_ctrl_reg2hw_csr0_reg_t;

  typedef struct packed {
    struct packed {
      logic [6:0]  q;
    } field0;
    struct packed {
      logic        q;
    } field1;
    struct packed {
      logic [6:0]  q;
    } field2;
    struct packed {
      logic        q;
    } field3;
    struct packed {
      logic [15:0] q;
    } field4;
  } otp_ctrl_reg2hw_csr1_reg_t;

  typedef struct packed {
    logic        q;
  } otp_ctrl_reg2hw_csr2_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  q;
    } field0;
    struct packed {
      logic [9:0] q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic        q;
    } field3;
    struct packed {
      logic        q;
    } field4;
    struct packed {
      logic        q;
    } field5;
    struct packed {
      logic        q;
    } field6;
    struct packed {
      logic        q;
    } field7;
    struct packed {
      logic        q;
    } field8;
  } otp_ctrl_reg2hw_csr3_reg_t;

  typedef struct packed {
    struct packed {
      logic [9:0] q;
    } field0;
    struct packed {
      logic        q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic        q;
    } field3;
  } otp_ctrl_reg2hw_csr4_reg_t;

  typedef struct packed {
    struct packed {
      logic [5:0]  q;
    } field0;
    struct packed {
      logic [1:0]  q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic [2:0]  q;
    } field3;
    struct packed {
      logic        q;
    } field4;
    struct packed {
      logic        q;
    } field5;
    struct packed {
      logic [15:0] q;
    } field6;
  } otp_ctrl_reg2hw_csr5_reg_t;

  typedef struct packed {
    struct packed {
      logic [9:0] q;
    } field0;
    struct packed {
      logic        q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic [15:0] q;
    } field3;
  } otp_ctrl_reg2hw_csr6_reg_t;

  typedef struct packed {
    struct packed {
      logic [5:0]  q;
    } field0;
    struct packed {
      logic [2:0]  q;
    } field1;
    struct packed {
      logic        q;
    } field2;
    struct packed {
      logic        q;
    } field3;
  } otp_ctrl_reg2hw_csr7_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  d;
      logic        de;
    } field0;
    struct packed {
      logic [9:0] d;
      logic        de;
    } field1;
    struct packed {
      logic        d;
      logic        de;
    } field2;
    struct packed {
      logic        d;
      logic        de;
    } field3;
    struct packed {
      logic        d;
      logic        de;
    } field4;
    struct packed {
      logic        d;
      logic        de;
    } field5;
    struct packed {
      logic        d;
      logic        de;
    } field6;
    struct packed {
      logic        d;
      logic        de;
    } field7;
    struct packed {
      logic        d;
      logic        de;
    } field8;
  } otp_ctrl_hw2reg_csr3_reg_t;

  typedef struct packed {
    struct packed {
      logic [5:0]  d;
      logic        de;
    } field0;
    struct packed {
      logic [1:0]  d;
      logic        de;
    } field1;
    struct packed {
      logic        d;
      logic        de;
    } field2;
    struct packed {
      logic [2:0]  d;
      logic        de;
    } field3;
    struct packed {
      logic        d;
      logic        de;
    } field4;
    struct packed {
      logic        d;
      logic        de;
    } field5;
    struct packed {
      logic [15:0] d;
      logic        de;
    } field6;
  } otp_ctrl_hw2reg_csr5_reg_t;

  typedef struct packed {
    struct packed {
      logic [5:0]  d;
      logic        de;
    } field0;
    struct packed {
      logic [2:0]  d;
      logic        de;
    } field1;
    struct packed {
      logic        d;
      logic        de;
    } field2;
    struct packed {
      logic        d;
      logic        de;
    } field3;
  } otp_ctrl_hw2reg_csr7_reg_t;

  // Register -> HW type for prim interface
  typedef struct packed {
    otp_ctrl_reg2hw_csr0_reg_t csr0; // [158:135]
    otp_ctrl_reg2hw_csr1_reg_t csr1; // [134:103]
    otp_ctrl_reg2hw_csr2_reg_t csr2; // [102:102]
    otp_ctrl_reg2hw_csr3_reg_t csr3; // [101:82]
    otp_ctrl_reg2hw_csr4_reg_t csr4; // [81:69]
    otp_ctrl_reg2hw_csr5_reg_t csr5; // [68:39]
    otp_ctrl_reg2hw_csr6_reg_t csr6; // [38:11]
    otp_ctrl_reg2hw_csr7_reg_t csr7; // [10:0]
  } otp_ctrl_prim_reg2hw_t;

  // HW -> register type for prim interface
  typedef struct packed {
    otp_ctrl_hw2reg_csr3_reg_t csr3; // [80:52]
    otp_ctrl_hw2reg_csr5_reg_t csr5; // [51:15]
    otp_ctrl_hw2reg_csr7_reg_t csr7; // [14:0]
  } otp_ctrl_prim_hw2reg_t;

  // Register offsets for prim interface
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR0_OFFSET = 5'h 0;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR1_OFFSET = 5'h 4;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR2_OFFSET = 5'h 8;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR3_OFFSET = 5'h c;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR4_OFFSET = 5'h 10;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR5_OFFSET = 5'h 14;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR6_OFFSET = 5'h 18;
  parameter logic [PrimAw-1:0] OTP_CTRL_CSR7_OFFSET = 5'h 1c;

  // Register index for prim interface
  typedef enum int {
    OTP_CTRL_CSR0,
    OTP_CTRL_CSR1,
    OTP_CTRL_CSR2,
    OTP_CTRL_CSR3,
    OTP_CTRL_CSR4,
    OTP_CTRL_CSR5,
    OTP_CTRL_CSR6,
    OTP_CTRL_CSR7
  } otp_ctrl_prim_id_e;

  // Register width information to check illegal writes for prim interface
  parameter logic [3:0] OTP_CTRL_PRIM_PERMIT [8] = '{
    4'b 1111, // index[0] OTP_CTRL_CSR0
    4'b 1111, // index[1] OTP_CTRL_CSR1
    4'b 0001, // index[2] OTP_CTRL_CSR2
    4'b 0111, // index[3] OTP_CTRL_CSR3
    4'b 0011, // index[4] OTP_CTRL_CSR4
    4'b 1111, // index[5] OTP_CTRL_CSR5
    4'b 1111, // index[6] OTP_CTRL_CSR6
    4'b 0011  // index[7] OTP_CTRL_CSR7
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package top_pkg;

localparam int TL_AW=32;
localparam int TL_DW=32;    // = TL_DBW * 8; TL_DBW must be a power-of-two
localparam int TL_AIW=8;    // a_source, d_source
localparam int TL_DIW=1;    // d_sink
localparam int TL_AUW=21;   // a_user
localparam int TL_DUW=14;   // d_user
localparam int TL_DBW=(TL_DW>>3);
localparam int TL_SZW=$clog2($clog2(TL_DBW)+1);

localparam int TL_DW64=64;    // = TL_DBW * 8; TL_DBW must be a power-of-two
localparam int TL_DBW64=(TL_DW64>>3);
localparam int TL_SZW64=$clog2($clog2(TL_DBW64)+1); //2

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// tl_main package generated by `tlgen.py` tool

package tl_main_rot_pkg;

   // localparam logic [31:0] ADDR_SPACE_ROM_CTRL__ROM_ROT        = 32'h 00008000;
  // localparam logic [31:0] ADDR_SPACE_ROM_CTRL__REGS_ROT       = 32'h 411e0000;
  // localparam logic [31:0] ADDR_SPACE_HMAC_ROT                 = 32'h 41110000;
  // localparam logic [31:0] ADDR_SPACE_KMAC_ROT                 = 32'h 41120000;
  // localparam logic [31:0] ADDR_SPACE_ENTROPY_SRC_ROT          = 32'h 41160000;
  // localparam logic [31:0] ADDR_SPACE_CSRNG_ROT                = 32'h 41150000;
  // localparam logic [31:0] ADDR_SPACE_EDN0_ROT                 = 32'h 41170000;
  // localparam logic [31:0] ADDR_SPACE_KEYMGR_ROT               = 32'h 41140000;

  localparam logic [31:0] ADDR_SPACE_ROM_CTRL__ROM_ROT        = 32'h 3b200000;
  localparam logic [31:0] ADDR_SPACE_RSTMGR_ROT               = 32'h 3b010000;
  localparam logic [31:0] ADDR_SPACE_ROM_CTRL__REGS_ROT       = 32'h 3b1e0000;
  localparam logic [31:0] ADDR_SPACE_HMAC_ROT                 = 32'h 3b110000;
  localparam logic [31:0] ADDR_SPACE_KMAC_ROT                 = 32'h 3b120000;
  localparam logic [31:0] ADDR_SPACE_ENTROPY_SRC_ROT          = 32'h 3b160000;
  localparam logic [31:0] ADDR_SPACE_CSRNG_ROT                = 32'h 3b150000;
  localparam logic [31:0] ADDR_SPACE_EDN0_ROT                 = 32'h 3b190000;
  localparam logic [31:0] ADDR_SPACE_KEYMGR_ROT               = 32'h 3b140000;
  localparam logic [31:0] ADDR_SPACE_OTBN_ROT                 = 32'h 3b130000;
  localparam logic [31:0] ADDR_SPACE_SM3                      = 32'h 3b1a0000;
  localparam logic [31:0] ADDR_SPACE_SM4                      = 32'h 3b1b0000;
  localparam logic [31:0] ADDR_SPACE_RS_ENCODE                = 32'h 3b170000;
  localparam logic [31:0] ADDR_SPACE_RS_DECODE                = 32'h 3b180000;
  localparam logic [31:0] ADDR_SPACE_PUF                      = 32'h 3b1c0000;
  localparam logic [31:0] ADDR_SPACE_PUF2                     = 32'h 3b1d0000;
  
  // localparam logic [31:0] ADDR_SPACE_ROM_CTRL__ROM_ROT        = 32'h 44008000;
  // localparam logic [31:0] ADDR_SPACE_ROM_CTRL__REGS_ROT       = 32'h 411e0000;
  // localparam logic [31:0] ADDR_SPACE_HMAC_ROT                 = 32'h 41110000;
  // localparam logic [31:0] ADDR_SPACE_KMAC_ROT                 = 32'h 41120000;
  // localparam logic [31:0] ADDR_SPACE_ENTROPY_SRC_ROT          = 32'h 41160000;
  // localparam logic [31:0] ADDR_SPACE_CSRNG_ROT                = 32'h 41150000;
  // localparam logic [31:0] ADDR_SPACE_EDN0_ROT                 = 32'h 41190000;
  // localparam logic [31:0] ADDR_SPACE_KEYMGR_ROT               = 32'h 41140000;
  
  localparam logic [31:0] ADDR_MASK_ROM_CTRL__ROM_ROT        = 32'h 00007fff;
  localparam logic [31:0] ADDR_MASK_ROM_CTRL__REGS_ROT       = 32'h 0000007f;
  localparam logic [31:0] ADDR_MASK_HMAC_ROT                 = 32'h 00000fff;
  localparam logic [31:0] ADDR_MASK_KMAC_ROT                 = 32'h 00000fff;
  localparam logic [31:0] ADDR_MASK_ENTROPY_SRC_ROT          = 32'h 000000ff;
  localparam logic [31:0] ADDR_MASK_CSRNG_ROT                = 32'h 0000007f;
  localparam logic [31:0] ADDR_MASK_EDN0_ROT                 = 32'h 0000007f;
  localparam logic [31:0] ADDR_MASK_KEYMGR_ROT               = 32'h 000000ff;
  localparam logic [31:0] ADDR_MASK_OTBN_ROT                 = 32'h 0000ffff;
  localparam logic [31:0] ADDR_MASK_SM3                      = 32'h 0000003f;
  localparam logic [31:0] ADDR_MASK_SM4                      = 32'h 0000003f;
  localparam logic [31:0] ADDR_MASK_RS_ENCODE                = 32'h 000001ff;
  localparam logic [31:0] ADDR_MASK_RS_DECODE                = 32'h 000001ff;
  localparam logic [31:0] ADDR_MASK_PUF                      = 32'h 0000003f;
  localparam logic [31:0] ADDR_MASK_PUF2                     = 32'h 0000003f;

  localparam int N_HOST   = 1;
  localparam int N_DEVICE = 15;

  typedef enum int {
    TlRomCtrlRom = 0,
    TlRomCtrlRegs = 1,
    TlHmac = 2,
    TlKmac = 3,
    TlEntropySrc = 4,
    TlCsrng = 5,
    TlEdn0 = 6,
    TlKeymgr = 7,
    TlOtbn = 8,
    TlSm3 = 9,
    TlSm4 = 10,
    TlRsEncode = 11,
    TlRsDecode = 12,
    TlPuf = 13,
    TlPuf2 = 14
  } tl_device_e;

  typedef enum int {
    TlRvCoreIbexCorei = 0,
    TlRvCoreIbexCored = 1,
    TlRvDmSba = 2
  } tl_host_e;

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`ifdef UVM
  `include "uvm_macros.svh"
`endif

// UVM speficic macros
`ifndef gfn
`ifdef UVM
  // verilog_lint: waive macro-name-style
  `define gfn get_full_name()
`else
  // verilog_lint: waive macro-name-style
  `define gfn $sformatf("%m")
`endif
`endif

`ifndef gtn
  // verilog_lint: waive macro-name-style
  `define gtn get_type_name()
`endif

`ifndef gn
  // verilog_lint: waive macro-name-style
  `define gn get_name()
`endif

`ifndef gmv
  // verilog_lint: waive macro-name-style
  `define gmv(csr) csr.get_mirrored_value()
`endif

// cast base class obj holding extended class handle to extended class handle;
// throw error if cast fails
`ifndef downcast
  // verilog_lint: waive macro-name-style
  `define downcast(EXT_, BASE_, MSG_="", SEV_=fatal, ID_=`gfn) \
    begin \
      if (!$cast(EXT_, BASE_)) begin \
        `dv_``SEV_($sformatf({"Cast failed: base class variable %0s ", \
                              "does not hold extended class %0s handle %s"}, \
                              `"BASE_`", `"EXT_`", MSG_), ID_) \
      end \
    end
`endif

// Note, UVM provides a macro `uvm_new_func -- which only applies to uvm_components
`ifndef uvm_object_new
  `define uvm_object_new \
    function new (string name=""); \
      super.new(name); \
    endfunction : new
`endif

`ifndef uvm_create_obj
  `define uvm_create_obj(_type_name_, _inst_name_) \
    _inst_name_ = _type_name_::type_id::create(`"_inst_name_`");
`endif

`ifndef uvm_component_new
  `define uvm_component_new \
    function new (string name="", uvm_component parent=null); \
      super.new(name, parent); \
    endfunction : new
`endif

`ifndef uvm_create_comp
  `define uvm_create_comp(_type_name_, _inst_name_) \
    _inst_name_ = _type_name_::type_id::create(`"_inst_name_`", this);
`endif

// Convert arbitrary text / expression to string.
`ifndef DV_STRINGIFY
  `define DV_STRINGIFY(I_) `"I_`"
`endif

`ifndef DUT_HIER_STR
  `define DUT_HIER_STR `DV_STRINGIFY(`DUT_HIER)
`endif

// Common check macros used by DV_CHECK error and fatal macros.
// Note: Should not be called by user code
`ifndef DV_CHECK
  `define DV_CHECK(T_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if (T_) ; else begin \
        `dv_``SEV_($sformatf("Check failed (%s) %s ", `"T_`", MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_EQ
  `define DV_CHECK_EQ(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) == (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s == %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_NE
  `define DV_CHECK_NE(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) != (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s != %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_CASE_EQ
  `define DV_CHECK_CASE_EQ(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) === (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s === %s (0x%0h [%0b] vs 0x%0h [%0b]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_CASE_NE
  `define DV_CHECK_CASE_NE(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) !== (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s !== %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_LT
  `define DV_CHECK_LT(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) < (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s < %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_GT
  `define DV_CHECK_GT(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) > (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s > %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_LE
  `define DV_CHECK_LE(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) <= (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s <= %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_GE
  `define DV_CHECK_GE(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) >= (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed %s >= %s (%0d [0x%0h] vs %0d [0x%0h]) %s", \
                             `"ACT_`", `"EXP_`", ACT_, ACT_, EXP_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_STREQ
  `define DV_CHECK_STREQ(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) == (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed \"%s\" == \"%s\" %s", ACT_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_STRNE
  `define DV_CHECK_STRNE(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      if ((ACT_) != (EXP_)) ; else begin \
        `dv_``SEV_($sformatf("Check failed \"%s\" != \"%s\" %s", ACT_, EXP_, MSG_), ID_) \
      end \
    end
`endif

`ifndef DV_CHECK_Q_EQ
  `define DV_CHECK_Q_EQ(ACT_, EXP_, MSG_="", SEV_=error, ID_=`gfn) \
    begin \
      `DV_CHECK_EQ(ACT_.size(), EXP_.size(), MSG_, SEV_, ID_) \
      foreach (ACT_[i]) begin \
        `DV_CHECK_EQ(ACT_[i], EXP_[i], $sformatf("for i = %0d %s", i, MSG_), SEV_, ID_) \
      end \
    end
`endif

// Fatal version of the checks
`ifndef DV_CHECK_FATAL
  `define DV_CHECK_FATAL(T_, MSG_="", ID_=`gfn) \
    `DV_CHECK(T_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_EQ_FATAL
  `define DV_CHECK_EQ_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_EQ(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_NE_FATAL
  `define DV_CHECK_NE_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_NE(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_LT_FATAL
  `define DV_CHECK_LT_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_LT(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_GT_FATAL
  `define DV_CHECK_GT_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_GT(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_LE_FATAL
  `define DV_CHECK_LE_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_LE(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_GE_FATAL
  `define DV_CHECK_GE_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_GE(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_STREQ_FATAL
  `define DV_CHECK_STREQ_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_STREQ(ACT_, EXP_, MSG_, fatal, ID_)
`endif

`ifndef DV_CHECK_STRNE_FATAL
  `define DV_CHECK_STRNE_FATAL(ACT_, EXP_, MSG_="", ID_=`gfn) \
    `DV_CHECK_STRNE(ACT_, EXP_, MSG_, fatal, ID_)
`endif

// Shorthand for common foo.randomize() + fatal check
`ifndef DV_CHECK_RANDOMIZE_FATAL
  `define DV_CHECK_RANDOMIZE_FATAL(VAR_, MSG_="Randomization failed!", ID_=`gfn) \
    `DV_CHECK_FATAL(VAR_.randomize(), MSG_, ID_)
`endif

// Shorthand for common foo.randomize() with { } + fatal check
`ifndef DV_CHECK_RANDOMIZE_WITH_FATAL
  `define DV_CHECK_RANDOMIZE_WITH_FATAL(VAR_, WITH_C_, MSG_="Randomization failed!", ID_=`gfn) \
    `DV_CHECK_FATAL(VAR_.randomize() with {WITH_C_}, MSG_, ID_)
`endif

// Shorthand for common std::randomize(foo) + fatal check
`ifndef DV_CHECK_STD_RANDOMIZE_FATAL
  `define DV_CHECK_STD_RANDOMIZE_FATAL(VAR_, MSG_="Randomization failed!", ID_=`gfn) \
    `DV_CHECK_FATAL(std::randomize(VAR_), MSG_, ID_)
`endif

// Shorthand for common std::randomize(foo) with { } + fatal check
`ifndef DV_CHECK_STD_RANDOMIZE_WITH_FATAL
  `define DV_CHECK_STD_RANDOMIZE_WITH_FATAL(VAR_, WITH_C_, MSG_="Randomization failed!",ID_=`gfn) \
    `DV_CHECK_FATAL(std::randomize(VAR_) with {WITH_C_}, MSG_, ID_)
`endif

// Shorthand for common cls_inst.randomize(member) + fatal check
// Randomizes a specific member of a class instance.
`ifndef DV_CHECK_MEMBER_RANDOMIZE_FATAL
  `define DV_CHECK_MEMBER_RANDOMIZE_FATAL(VAR_, CLS_INST_=this, MSG_="Randomization failed!", ID_=`gfn) \
    `DV_CHECK_FATAL(CLS_INST_.randomize(VAR_), MSG_, ID_)
`endif

// Shorthand for common cls_inst.randomize(member) with { } + fatal check
// Randomizes a specific member of a class instance with inline constraints.
`ifndef DV_CHECK_MEMBER_RANDOMIZE_WITH_FATAL
  `define DV_CHECK_MEMBER_RANDOMIZE_WITH_FATAL(VAR_, C_, CLS_INST_=this, MSG_="Randomization failed!", ID_=`gfn) \
    `DV_CHECK_FATAL(CLS_INST_.randomize(VAR_) with {C_}, MSG_, ID_)
`endif

// print static/dynamic 1d array or queue
`ifndef DV_PRINT_ARR_CONTENTS
`define DV_PRINT_ARR_CONTENTS(ARR_, V_=uvm_pkg::UVM_MEDIUM, ID_=`gfn) \
  begin \
    foreach (ARR_[i]) begin \
      `dv_info($sformatf("%s[%0d] = %0d (0x%0h)", `"ARR_`", i, ARR_[i], ARR_[i]), V_, ID_) \
    end \
  end
`endif

// print non-empty tlm fifos that were uncompared at end of test
`ifndef DV_EOT_PRINT_TLM_FIFO_CONTENTS
`define DV_EOT_PRINT_TLM_FIFO_CONTENTS(TYP_, FIFO_, SEV_=error, ID_=`gfn) \
  begin \
    while (!FIFO_.is_empty()) begin \
      TYP_ item; \
      void'(FIFO_.try_get(item)); \
      `dv_``SEV_($sformatf("%s item uncompared:\n%s", `"FIFO_`", item.sprint()), ID_) \
    end \
  end
`endif

// print non-empty tlm fifos that were uncompared at end of test
`ifndef DV_EOT_PRINT_TLM_FIFO_ARR_CONTENTS
`define DV_EOT_PRINT_TLM_FIFO_ARR_CONTENTS(TYP_, FIFO_, SEV_=error, ID_=`gfn) \
  begin \
    foreach (FIFO_[i]) begin \
      while (!FIFO_[i].is_empty()) begin \
        TYP_ item; \
        void'(FIFO_[i].try_get(item)); \
        `dv_``SEV_($sformatf("%s[%0d] item uncompared:\n%s", `"FIFO_`", i, item.sprint()), ID_) \
      end \
    end \
  end
`endif

// print non-empty tlm fifos that were uncompared at end of test
`ifndef DV_EOT_PRINT_Q_CONTENTS
`define DV_EOT_PRINT_Q_CONTENTS(TYP_, Q_, SEV_=error, ID_=`gfn) \
  begin \
    while (Q_.size() != 0) begin \
      TYP_ item = Q_.pop_front(); \
      `dv_``SEV_($sformatf("%s item uncompared:\n%s", `"Q_`", item.sprint()), ID_) \
    end \
  end
`endif

// print non-empty tlm fifos that were uncompared at end of test
`ifndef DV_EOT_PRINT_Q_ARR_CONTENTS
`define DV_EOT_PRINT_Q_ARR_CONTENTS(TYP_, Q_, SEV_=error, ID_=`gfn) \
  begin \
    foreach (Q_[i]) begin \
      while (Q_[i].size() != 0) begin \
        TYP_ item = Q_[i].pop_front(); \
        `dv_``SEV_($sformatf("%s[%0d] item uncompared:\n%s", `"Q_`", i, item.sprint()), ID_) \
      end \
    end \
  end
`endif

// check for non-empty mailbox and print items that were uncompared at end of test
`ifndef DV_EOT_PRINT_MAILBOX_CONTENTS
`define DV_EOT_PRINT_MAILBOX_CONTENTS(TYP_, MAILBOX_, SEV_=error, ID_=`gfn) \
  begin \
    while (MAILBOX_.num() != 0) begin \
      TYP_ item; \
      void'(MAILBOX_.try_get(item)); \
      `dv_``SEV_($sformatf("%s item uncompared:\n%s", `"MAILBOX_`", item.sprint()), ID_) \
    end \
  end
`endif

// get parity - implemented as a macro so that it can be invoked in constraints as well
`ifndef GET_PARITY
  `define GET_PARITY(val, odd=0) (^val ^ odd)
`endif

// Wait a task or statement with exit condition
// Kill the thread when either the wait statement is completed or exit condition occurs
// input WAIT_ need to be a statement. Here are some examples
// `DV_SPINWAIT(wait(...);, "Wait for ...")
// `DV_SPINWAIT(
//              while (1) begin
//                ...
//              end)
`ifndef DV_SPINWAIT_EXIT
`define DV_SPINWAIT_EXIT(WAIT_, EXIT_, MSG_ = "exit condition occurred!", ID_ =`gfn) \
  begin \
    fork begin \
      fork \
        begin \
          WAIT_ \
        end \
        begin \
          EXIT_ \
          if (MSG_ != "") begin \
            `dv_info(MSG_, uvm_pkg::UVM_HIGH, ID_) \
          end \
        end \
      join_any \
      disable fork; \
    end join \
  end
`endif

// macro that waits for a given delay and then reports an error
`ifndef DV_WAIT_TIMEOUT
`define DV_WAIT_TIMEOUT(TIMEOUT_NS_, ID_  = `gfn, ERROR_MSG_ = "timeout occurred!", REPORT_FATAL_ = 1) \
  begin \
    #(TIMEOUT_NS_ * 1ns); \
    if (REPORT_FATAL_) `dv_fatal(ERROR_MSG_, ID_) \
    else               `dv_error(ERROR_MSG_, ID_) \
  end
`endif

// wait a task or statement with timer watchdog
`ifndef DV_SPINWAIT
`define DV_SPINWAIT(WAIT_, MSG_ = "timeout occurred!", TIMEOUT_NS_ = default_spinwait_timeout_ns, ID_ =`gfn) \
  `DV_SPINWAIT_EXIT(WAIT_, `DV_WAIT_TIMEOUT(TIMEOUT_NS_, ID_, MSG_);, "", ID_)
`endif

// a shorthand of `DV_SPINWAIT(wait(...))
`ifndef DV_WAIT
`define DV_WAIT(WAIT_COND_, MSG_ = "wait timeout occurred!", TIMEOUT_NS_ = default_spinwait_timeout_ns, ID_ =`gfn) \
  `DV_SPINWAIT(wait (WAIT_COND_);, MSG_, TIMEOUT_NS_, ID_)
`endif

// Control assertions in the DUT.
//
// This macro is invoked in top level testbench that instantiates the DUT. It spawns off an initial
// block that forever waits for a resource of type bit named by the string arg ~LABEL_~ that
// can be set by any entity in the testbench. Based on the value set, it enables or disables the
// assertions at the hierarchy of the provided path. The entity setting the resource value invokes
// uvm_config_db#(bit)::set(...) and this macro calls the corresponding get.
//
// LABEL_ : Name of the assertion control resource bit (string).
// HIER_  : Path to the module within which the assertion is controlled.
// LEVELS_: Number of levels within the module to control the assertions.
// SCOPE_ : Hierarchical string path to the testbench where this macro is invoked, example: %m.
// ID_    : Identifier string used for UVM logs.
`ifndef DV_ASSERT_CTRL
`define DV_ASSERT_CTRL(LABEL_, HIER_, LEVELS_ = 0, SCOPE_ = "", ID_ = $sformatf("%m")) \
  initial begin \
    bit assert_en; \
    forever begin \
      uvm_config_db#(bit)::wait_modified(null, SCOPE_, LABEL_); \
      if (!uvm_config_db#(bit)::get(null, SCOPE_, LABEL_, assert_en)) begin \
        `uvm_fatal(ID_, $sformatf("Failed to get \"%0s\" from uvm_config_db", LABEL_)) \
      end \
      if (assert_en) begin \
        `uvm_info(ID_, $sformatf("Enabling assertions: %0s", `DV_STRINGIFY(HIER_)), UVM_LOW) \
        $asserton(LEVELS_, HIER_); \
      end else begin \
        `uvm_info(ID_, $sformatf("Disabling assertions: %0s", `DV_STRINGIFY(HIER_)), UVM_LOW) \
        $assertoff(LEVELS_, HIER_); \
        $assertkill(LEVELS_, HIER_); \
      end \
    end \
  end
`endif

// Retrieves a plusarg value representing an enum literal.
//
// The plusarg is parsed as a string, which needs to be converted into the enum literal whose name
// matches the string. This functionality is provided by the UVM helper function below.
//
// ENUM_: The enum type.
// VAR_: The enum variable to which the plusarg value will be set (must be declared already).
// PLUSARG_: the name of the plusarg (as raw text). This is typically the same as the enum variable.
// CHECK_EXISTS_: Throws a fatal error if the plusarg is not set.
`ifndef DV_GET_ENUM_PLUSARG
`define DV_GET_ENUM_PLUSARG(ENUM_, VAR_, PLUSARG_, CHECK_EXISTS_ = 0, ID_ = `gfn) \
  begin \
    string str; \
    if ($value$plusargs(`"``PLUSARG_``=%0s`", str)) begin \
      if (!uvm_enum_wrapper#(ENUM_)::from_name(str, VAR_)) begin \
        `uvm_fatal(ID_, $sformatf(`"Cannot find %s from enum ``ENUM_```", VAR_.name())) \
      end \
    end else if (CHECK_EXISTS_) begin \
      `uvm_fatal(ID_, `"Please pass the plusarg +``PLUSARG_``=<``ENUM_``-literal>`") \
    end \
  end
`endif

// Retrieves a queue of plusarg value from a string.
//
// The plusarg is parsed as a string, which needs to be converted into a queue of string which given delimiter.
// This functionality is provided by the UVM helper function below.
//
// QUEUE_: The queue of string to which the plusarg value will be set (must be declared already).
// PLUSARG_: the name of the plusarg (as raw text). This is typically the same as the enum variable.
// DELIMITER_: the delimiter that separate each item in the plusarg string value.
// CHECK_EXISTS_: Throws a fatal error if the plusarg is not set.
`ifndef DV_GET_QUEUE_PLUSARG
`define DV_GET_QUEUE_PLUSARG(QUEUE_, PLUSARG_, DELIMITER_ = ",", CHECK_EXISTS_ = 0, ID_ = `gfn) \
  begin \
    string str; \
    if ($value$plusargs(`"``PLUSARG_``=%0s`", str)) begin \
      str_split(str, QUEUE_, DELIMITER_); \
    end else if (CHECK_EXISTS_) begin \
      `uvm_fatal(ID_, `"Please pass the plusarg +``PLUSARG_``=<``ENUM_``-literal>`") \
    end \
  end
`endif

// Enable / disable assertions at a module hierarchy identified by LABEL_.
//
// This goes in conjunction with `DV_ASSERT_CTRL() macro above, but is invoked in the entity that is
// sending the req to turn on / off the assertions. Note that piece of code invoking this macro
// does not have the information on the actual hierarchical path to the module or the levels - this
// is 'wrapped' into the LABEL_ instead. DV user needs to uniquify the label sufficienly enough to
// reflect it.
//
// LABEL_ : Name of the assertion control resource bit (string).
// VALUE_ : Value of the control bit - 1 - enable assertions, 0 - disable assertions.
// SCOPE_ : Hierarchical string path to the testbench where this macro is invoked, example: %m.
`ifndef DV_ASSERT_CTRL_REQ
`define DV_ASSERT_CTRL_REQ(LABEL_, VALUE_, SCOPE_="") \
  begin \
    uvm_config_db#(bit)::set(null, SCOPE_, LABEL_, VALUE_); \
  end
`endif

// Macros for logging (info, warning, error and fatal severities).
//
// These are meant to be invoked in modules and interfaces that are shared between DV and Verilator
// testbenches. We waive the lint requirement for these to be in uppercase, since they are
// UVM-adjacent.
`ifdef UVM
`ifndef dv_info
  // verilog_lint: waive macro-name-style
  `define dv_info(MSG_,  VERBOSITY_ = uvm_pkg::UVM_LOW, ID_ = $sformatf("%m")) \
    if (uvm_pkg::uvm_report_enabled(VERBOSITY_, uvm_pkg::UVM_INFO, ID_)) begin \
        uvm_pkg::uvm_report_info(ID_, MSG_, VERBOSITY_, `uvm_file, `uvm_line, "", 1); \
    end
`endif

`ifndef dv_warning
  // verilog_lint: waive macro-name-style
  `define dv_warning(MSG_, ID_ = $sformatf("%m")) \
    if (uvm_pkg::uvm_report_enabled(uvm_pkg::UVM_NONE, uvm_pkg::UVM_WARNING, ID_)) begin \
        uvm_pkg::uvm_report_warning(ID_, MSG_, uvm_pkg::UVM_NONE, `uvm_file, `uvm_line, "", 1); \
    end
`endif

`ifndef dv_error
  // verilog_lint: waive macro-name-style
  `define dv_error(MSG_, ID_ = $sformatf("%m")) \
    if (uvm_pkg::uvm_report_enabled(uvm_pkg::UVM_NONE, uvm_pkg::UVM_ERROR, ID_)) begin \
        uvm_pkg::uvm_report_error(ID_, MSG_, uvm_pkg::UVM_NONE, `uvm_file, `uvm_line, "", 1); \
    end
`endif

`ifndef dv_fatal
  // verilog_lint: waive macro-name-style
  `define dv_fatal(MSG_, ID_ = $sformatf("%m")) \
    if (uvm_pkg::uvm_report_enabled(uvm_pkg::UVM_NONE, uvm_pkg::UVM_FATAL, ID_)) begin \
        uvm_pkg::uvm_report_fatal(ID_, MSG_, uvm_pkg::UVM_NONE, `uvm_file, `uvm_line, "", 1); \
    end
`endif

`else // UVM

`ifndef dv_info
  // verilog_lint: waive macro-name-style
  `define dv_info(MSG_, VERBOSITY = DUMMY_, ID_ = $sformatf("%m")) \
    $display("%0t: (%0s:%0d) [%0s] %0s", $time, `__FILE__, `__LINE__, ID_, MSG_);
`endif

`ifndef dv_warning
  // verilog_lint: waive macro-name-style
  `define dv_warning(MSG_, ID_ = $sformatf("%m")) \
    $warning("%0t: (%0s:%0d) [%0s] %0s", $time, `__FILE__, `__LINE__, ID_, MSG_);
`endif

`ifndef dv_error
  // verilog_lint: waive macro-name-style
  `define dv_error(MSG_, ID_ = $sformatf("%m")) \
    $error("%0t: (%0s:%0d) [%0s] %0s", $time, `__FILE__, `__LINE__, ID_, MSG_);
`endif

`ifndef dv_fatal
  // verilog_lint: waive macro-name-style
  `define dv_fatal(MSG_, ID_ = $sformatf("%m")) \
    $fatal(1, "%0t: (%0s:%0d) [%0s] %0s", $time, `__FILE__, `__LINE__, ID_, MSG_);
`endif

`endif // UVM

// Macros for constrain clk with common frequencies
//
// Nominal clock frequency range is 24Mhz - 100Mhz and use higher weights on 24, 25, 48, 50, 100,
// To mimic manufacturing conditions (when clocks are uncalibrated), we need to be able to go as
// low as 5MHz.
`ifndef DV_COMMON_CLK_CONSTRAINT
`define DV_COMMON_CLK_CONSTRAINT(FREQ_) \
  FREQ_ dist { \
    [5:23]  :/ 2, \
    [24:25] :/ 2, \
    [26:47] :/ 1, \
    [48:50] :/ 2, \
    [51:95] :/ 1, \
    96      :/ 1, \
    [97:99] :/ 1, \
    100     :/ 1  \
  };
`endif

// Enables build-time randomization of fixed design constants.
//
// This is meant to be overridden externally by passing `+define+BUILD_SEED=<value>`.
`ifndef BUILD_SEED
  `define BUILD_SEED 1
`endif

// Max value out of 2 given expressions.
//
// Duplicate of dv_utils_pkg::max2() function, but this is better because
// it can consume different data types directly without the need for casting.
`ifndef DV_MAX2
  `define DV_MAX2(a, b) ((a) > (b) ? (a) : (b))
`endif

// Creates a signal probe function to sample / force / release an internal signal.
//
// If there is a need to sample / force an internal signal, then it must be done in the testbench,
// or in an interface bound to the DUT. This macro creates a standardized signal probe function
// meant to be invoked an interface. The generated function can then be invoked in test sequences
// or other UVM classes. The macro takes 2 arguments - name of the function and the hierarchical
// path to the signal. If invoked in an interface which is bound to the DUT, the signal can be a
// partial hierarchical path within the DUT. The generated function accepts 2 arguments - the first
// indicates the probe action (sample, force or release) of type dv_utils_pkg::signal_probe_e. The
// second argument is the value to be forced. If sample action is chosen, then it returns the
// sampled value (for other actions as well).
//
// The suggested naming convention for the function is:
//   signal_probe_<DUT_or_IP_block_name>_<signal_name>
//
// This macro must be invoked in an interface or module.
`ifndef DV_CREATE_SIGNAL_PROBE_FUNCTION
`define DV_CREATE_SIGNAL_PROBE_FUNCTION(FUNC_NAME_, SIGNAL_PATH_, SIGNAL_WIDTH_ = uvm_pkg::UVM_HDL_MAX_WIDTH) \
  function static logic [SIGNAL_WIDTH_-1:0] FUNC_NAME_(dv_utils_pkg::signal_probe_e kind,     \
                                                       logic [SIGNAL_WIDTH_-1:0] value = '0); \
    case (kind)                                                                               \
      dv_utils_pkg::SignalProbeSample: ;                                                      \
      dv_utils_pkg::SignalProbeForce: force SIGNAL_PATH_ = value;                             \
      dv_utils_pkg::SignalProbeRelease: release SIGNAL_PATH_;                                 \
      default: `uvm_fatal(`"FUNC_NAME_`", $sformatf("Bad value: %0d", kind))                  \
    endcase                                                                                   \
    return SIGNAL_PATH_;                                                                      \
  endfunction
`endif

// Usage:`OTDBG(( string ))
// This macro has unque keyword 'OTDBG'and timestemp only.
// Use for the temporary print to distinguish from `uvm_info.
// Do not leave this macro in other source files in the remote repo.
`ifndef OTDBG
  `define OTDBG(x) \
  $write($sformatf("%t:OTDBG:",$time));\
  $display($sformatf x);
`endif


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Interface: pins_if
// Description: Pin interface for driving and sampling individual pins such as interrupts, alerts
// and gpios.
`ifndef SYNTHESIS

interface pins_if #(
  parameter int Width = 1,
  parameter bit [8*4-1:0] PullStrength = "Pull"
) (
  inout [Width-1:0] pins
);

  `include "prim_assert.sv"

  `ASSERT_INIT(PullStrengthParamValid, PullStrength inside {"Weak", "Pull"})

  logic [Width-1:0] pins_o;       // value to be driven out
  bit   [Width-1:0] pins_oe = '0; // output enable
  bit   [Width-1:0] pins_pd = '0; // pull down enable
  bit   [Width-1:0] pins_pu = '0; // pull up enable

  // function to set pin output enable for specific pin (useful for single pin interface)
  function automatic void drive_en_pin(int idx = 0, bit val);
    pins_oe[idx] = val;
  endfunction

  // function to set pin output enable for all pins
  function automatic void drive_en(bit [Width-1:0] val);
    pins_oe = val;
  endfunction

  // function to drive a specific pin with a value (useful for single pin interface)
  function automatic void drive_pin(int idx = 0, logic val);
    pins_oe[idx] = 1'b1;
    pins_o[idx] = val;
  endfunction // drive_pin

  // function to drive all pins
  function automatic void drive(logic [Width-1:0] val);
    pins_oe = {Width{1'b1}};
    pins_o = val;
  endfunction // drive

  // function to drive all pull down values
  function automatic void set_pulldown_en(bit [Width-1:0] val);
    pins_pd = val;
  endfunction // set_pulldown_en

  // function to drive all pull up values
  function automatic void set_pullup_en(bit [Width-1:0] val);
    pins_pu = val;
  endfunction // set_pullup_en

  // function to drive the pull down value on a specific pin
  function automatic void set_pulldown_en_pin(int idx = 0, bit val);
    pins_pd[idx] = val;
  endfunction // set_pulldown_en_pin

  // function to drive the pull up value on a specific pin
  function automatic void set_pullup_en_pin(int idx = 0, bit val);
    pins_pu[idx] = val;
  endfunction // set_pullup_en_pin

  // function to sample a specific pin (useful for single pin interface)
  function automatic logic sample_pin(int idx = 0);
    return pins[idx];
  endfunction

  // function to sample all pins
  function automatic logic [Width-1:0] sample();
    return pins;
  endfunction

  // Fully disconnect this interface, including the pulls.
  function automatic void disconnect();
    pins_oe = {Width{1'b0}};
    pins_pu = {Width{1'b0}};
    pins_pd = {Width{1'b0}};
  endfunction

  // make connections
  for (genvar i = 0; i < Width; i++) begin : gen_each_pin
`ifdef VERILATOR
    assign pins[i] = pins_oe[i] ? pins_o[i] :
                     pins_pu[i] ? 1'b1 :
                     pins_pd[i] ? 1'b0 : 1'bz;
`else
    // Drive the pin based on whether pullup / pulldown is enabled.
    //
    // If output is not enabled, then the pin is pulled up or down with the `PullStrength` strength
    // Pullup has priority over pulldown.
    if (PullStrength == "Pull") begin : gen_pull_strength_pull
      assign (pull0, pull1) pins[i] = ~pins_oe[i] ? (pins_pu[i] ? 1'b1 :
                                                     pins_pd[i] ? 1'b0 : 1'bz) : 1'bz;
    end : gen_pull_strength_pull
    else if (PullStrength == "Weak") begin : gen_pull_strength_weak
      assign (weak0, weak1) pins[i] = ~pins_oe[i] ? (pins_pu[i] ? 1'b1 :
                                                     pins_pd[i] ? 1'b0 : 1'bz) : 1'bz;
    end : gen_pull_strength_weak

    // If output enable is 1, strong driver assigns pin to 'value to be driven out';
    // the external strong driver can still affect pin, if exists.
    // Else if output enable is 0, weak pullup or pulldown is applied to pin.
    // By doing this, we make sure that weak pullup or pulldown does not override
    // any 'x' value on pin, that may result due to conflicting values
    // between 'value to be driven out' and the external driver's value.
    assign pins[i] = pins_oe[i] ? pins_o[i] : 1'bz;
`endif
  end : gen_each_pin

endinterface
`endif


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// State definitions for entropy_src_ack_sm, provided as a separate package for use in DV

package entropy_src_ack_sm_pkg;

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 3 -n 6 \
  //      -s 1236774883 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (33.33%)
  //  4: |||||||||||||||||||| (33.33%)
  //  5: |||||||||||||||||||| (33.33%)
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 5
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4
  //
  localparam int StateWidth = 6;
  typedef enum logic [StateWidth-1:0] {
    Idle  = 6'b011101, // idle
    Wait  = 6'b101100, // wait until the fifo has an entry
    Error = 6'b000010  // illegal state reached and hang
  } state_e;

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// State definitions for entropy_src_main_sm, provided as a separate package for use in DV

package entropy_src_main_sm_pkg;

// Encoding generated with:
// $ ./util/design/sparse-fsm-encode.py -d 3 -m 21 -n 9 \
//      -s 2359261201 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||| (19.05%)
//  4: |||||||||||||||||||| (30.48%)
//  5: ||||||||||||||||| (26.19%)
//  6: |||||||||| (15.71%)
//  7: ||| (5.71%)
//  8: | (2.38%)
//  9:  (0.48%)
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 9
// Minimum Hamming weight: 1
// Maximum Hamming weight: 8
//

  localparam int StateWidth = 9;

  typedef enum logic [StateWidth-1:0] {
    Idle              = 9'b011110101, // idle
    BootHTRunning     = 9'b111010010, // boot mode, wait for health test done pulse
    BootPostHTChk     = 9'b101101110, // boot mode, wait for post health test packer not empty state
    BootPhaseDone     = 9'b010001110, // boot mode, stay here until master enable is off
    StartupHTStart    = 9'b000101100, // startup mode, pulse the sha3 start input
    StartupPhase1     = 9'b100000001, // startup mode, look for first test pass/fail
    StartupPass1      = 9'b110100101, // startup mode, look for first test pass/fail, done if pass
    StartupFail1      = 9'b000010111, // startup mode, look for second fail, alert if fail
    ContHTStart       = 9'b001000000, // continuous test mode, pulse the sha3 start input
    ContHTRunning     = 9'b110100010, // continuous test mode, wait for health test done pulse
    FWInsertStart     = 9'b011000011, // fw ov mode, start the sha3 block
    FWInsertMsg       = 9'b001011001, // fw ov mode, insert fw message into sha3 block
    Sha3MsgDone       = 9'b100001111, // sha3 mode, all input messages added, ready to process
    Sha3Prep          = 9'b011111000, // sha3 mode, request csrng arb to reduce power
    Sha3Process       = 9'b010111111, // sha3 mode, pulse the sha3 process input
    Sha3Valid         = 9'b101110001, // sha3 mode, wait for sha3 valid indication
    Sha3Done          = 9'b110011000, // sha3 mode, capture sha3 result, pulse done input
    Sha3Quiesce       = 9'b111001101, // sha3 mode, goto alert state or continuous check mode
    AlertState        = 9'b111111011, // if some alert condition occurs, pulse an alert indication
    AlertHang         = 9'b101011100, // after pulsing alert signal, hang here until sw handles
    Error             = 9'b100111101  // illegal state reached and hang
  } state_e;

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package entropy_src_pkg;

  //-------------------------
  // Entropy Interface
  //-------------------------

  parameter int  RNG_BUS_WIDTH   = 4;
  parameter int  CSRNG_BUS_WIDTH = 384;
  parameter int  FIPS_BUS_WIDTH  = 1;
  parameter int  FIPS_CSRNG_BUS_WIDTH = FIPS_BUS_WIDTH + CSRNG_BUS_WIDTH;

  // es entropy i/f
  typedef struct packed {
    logic es_ack;
    logic [CSRNG_BUS_WIDTH-1:0] es_bits;
    logic [FIPS_BUS_WIDTH-1:0] es_fips;
  } entropy_src_hw_if_rsp_t;

  typedef struct packed {
    logic es_req;
  } entropy_src_hw_if_req_t;

  parameter entropy_src_hw_if_req_t ENTROPY_SRC_HW_IF_REQ_DEFAULT = '{default: '0};
  parameter entropy_src_hw_if_rsp_t ENTROPY_SRC_HW_IF_RSP_DEFAULT = '{default: '0};


  // csrng block encrypt request/ack i/f
  typedef struct packed {
    logic cs_aes_halt_req;
  } cs_aes_halt_req_t;

  typedef struct packed {
    logic cs_aes_halt_ack;
  } cs_aes_halt_rsp_t;

  parameter cs_aes_halt_req_t CS_AES_HALT_REQ_DEFAULT = '{default: '0};
  parameter cs_aes_halt_rsp_t CS_AES_HALT_RSP_DEFAULT = '{default: '0};

  // ast rng i/f
  typedef struct packed {
    logic rng_enable;
  } entropy_src_rng_req_t;

  typedef struct packed {
    logic rng_valid;
    logic [RNG_BUS_WIDTH-1:0] rng_b;
  } entropy_src_rng_rsp_t;

  parameter entropy_src_rng_req_t ENTROPY_SRC_RNG_REQ_DEFAULT = '{default: '0};
  parameter entropy_src_rng_rsp_t ENTROPY_SRC_RNG_RSP_DEFAULT = '{default: '0};

  // external health test i/f
  typedef struct packed {
    logic [RNG_BUS_WIDTH-1:0] entropy_bit;
    logic entropy_bit_valid;
    logic clear;
    logic active;
    logic [15:0] thresh_hi;
    logic [15:0] thresh_lo;
    logic [15:0] health_test_window;
    logic window_wrap_pulse;
    logic threshold_scope;
  } entropy_src_xht_req_t;

  typedef struct packed {
    logic[15:0] test_cnt_hi;
    logic[15:0] test_cnt_lo;
    logic continuous_test;
    logic test_fail_hi_pulse;
    logic test_fail_lo_pulse;
  } entropy_src_xht_rsp_t;

  parameter entropy_src_xht_req_t ENTROPY_SRC_XHT_REQ_DEFAULT = '{default: '0};
  parameter entropy_src_xht_rsp_t ENTROPY_SRC_XHT_RSP_DEFAULT =
      '{test_cnt_lo: 16'hffff, default: '0};

endpackage : entropy_src_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Constants for use in primitives

// This file is auto-generated.

package prim_pkg;

  // Implementation target specialization
  typedef enum integer {
    ImplGeneric
  } impl_e;
endpackage : prim_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Some generally useful macros for RTL.

// Determine if __actual equals __expected with a margin of __allowed_less and __allowed_more, i.e.,
// if __actual is in the interval [__expected - __allowed_less, __expected + __allowed_more], where
// lower and upper bounds are inclusive.
//
// The caller is responsible for ensuring that the data types are such that
// (1) __actual + __allowed_less
// (2) __expected + __allowed_more
// are well defined and do not overflow and
// (3) (1) >= __expected
// (4) __actual <= (2)
// are well defined and meaningful.  Subtractions are deliberately not used, in order to prevent
// underflows.
`define WITHIN_MARGIN(__actual, __expected, __allowed_less, __allowed_more) \
  (((__actual) + (__allowed_less) >= (__expected)) &&                       \
   ((__actual) <= (__expected) + (__allowed_more)))

// Coverage pragmas, used around code for which we want to disable coverage collection.
// Don't forget to add a closing ON pragma after the code to be skipped.
//
// Some notes:
// - The first line is for VCS, the second for xcelium. It is okay to issue both regardless of
//   the tool used.
// - For xcelium it is possible to discriminate between metrics to be disabled as follows
//   //pragma coverage <metric> = on/off
//   where metric can be block | expr | toggle | fsm.

// TODO(https://github.com/chipsalliance/verible/issues/1498) Verible seems to get confused
// by these macros, so the code will inline these directives until this is fixed.
/*
`ifndef PRAGMA_COVERAGE_OFF
`define PRAGMA_COVERAGE_OFF \
/``/VCS coverage off \
/``/ pragma coverage off
`endif

`ifndef PRAGMA_COVERAGE_ON
`define PRAGMA_COVERAGE_ON \
/``/VCS coverage on \
/``/ pragma coverage on
`endif
*/


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package prim_ram_1p_pkg;

  typedef struct packed {
    logic       cfg_en;
    logic [3:0] cfg;
  } cfg_t;

  typedef struct packed {
    cfg_t ram_cfg;  // configuration for ram
    cfg_t rf_cfg;   // configuration for regfile
  } ram_1p_cfg_t;

  parameter ram_1p_cfg_t RAM_1P_CFG_DEFAULT = '0;

endpackage // prim_ram_1p_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package prim_rom_pkg;

  typedef struct packed {
    logic       cfg_en;
    logic [3:0] cfg;
  } rom_cfg_t;

  parameter rom_cfg_t ROM_CFG_DEFAULT = '0;

endpackage // prim_rom_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This package holds common constants and functions for PRESENT- and
// PRINCE-based scrambling devices.
//
// See also: prim_present, prim_prince
//
// References: - https://en.wikipedia.org/wiki/PRESENT
//             - https://en.wikipedia.org/wiki/Prince_(cipher)
//             - http://www.lightweightcrypto.org/present/present_ches2007.pdf
//             - https://eprint.iacr.org/2012/529.pdf
//             - https://eprint.iacr.org/2015/372.pdf
//             - https://eprint.iacr.org/2014/656.pdf

package prim_cipher_pkg;

  ///////////////////
  // PRINCE Cipher //
  ///////////////////

  parameter logic [15:0][3:0] PRINCE_SBOX4 = {4'h4, 4'hD, 4'h5, 4'hE,
                                              4'h0, 4'h8, 4'h7, 4'h6,
                                              4'h1, 4'h9, 4'hC, 4'hA,
                                              4'h2, 4'h3, 4'hF, 4'hB};

  parameter logic [15:0][3:0] PRINCE_SBOX4_INV = {4'h1, 4'hC, 4'hE, 4'h5,
                                                  4'h0, 4'h4, 4'h6, 4'hA,
                                                  4'h9, 4'h8, 4'hD, 4'hF,
                                                  4'h2, 4'h3, 4'h7, 4'hB};
  // nibble permutations
  parameter logic [15:0][3:0] PRINCE_SHIFT_ROWS64  = '{4'hF, 4'hA, 4'h5, 4'h0,
                                                       4'hB, 4'h6, 4'h1, 4'hC,
                                                       4'h7, 4'h2, 4'hD, 4'h8,
                                                       4'h3, 4'hE, 4'h9, 4'h4};

  parameter logic [15:0][3:0] PRINCE_SHIFT_ROWS64_INV = '{4'hF, 4'h2, 4'h5, 4'h8,
                                                          4'hB, 4'hE, 4'h1, 4'h4,
                                                          4'h7, 4'hA, 4'hD, 4'h0,
                                                          4'h3, 4'h6, 4'h9, 4'hC};

  // these are the round constants
  parameter logic [11:0][63:0] PRINCE_ROUND_CONST = {64'hC0AC29B7C97C50DD,
                                                     64'hD3B5A399CA0C2399,
                                                     64'h64A51195E0E3610D,
                                                     64'hC882D32F25323C54,
                                                     64'h85840851F1AC43AA,
                                                     64'h7EF84F78FD955CB1,
                                                     64'hBE5466CF34E90C6C,
                                                     64'h452821E638D01377,
                                                     64'h082EFA98EC4E6C89,
                                                     64'hA4093822299F31D0,
                                                     64'h13198A2E03707344,
                                                     64'h0000000000000000};

  // tweak constant for key modification between enc/dec modes
  parameter logic [63:0] PRINCE_ALPHA_CONST = 64'hC0AC29B7C97C50DD;

  // masking constants for shift rows function below
  parameter logic [15:0] PRINCE_SHIFT_ROWS_CONST0 = 16'h7BDE;
  parameter logic [15:0] PRINCE_SHIFT_ROWS_CONST1 = 16'hBDE7;
  parameter logic [15:0] PRINCE_SHIFT_ROWS_CONST2 = 16'hDE7B;
  parameter logic [15:0] PRINCE_SHIFT_ROWS_CONST3 = 16'hE7BD;

  // nibble shifts
  function automatic logic [31:0] prince_shiftrows_32bit(logic [31:0]      state_in,
                                                         logic [15:0][3:0] shifts );
    logic [31:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 32/2; k++) begin
      // operate on pairs of 2bit instead of nibbles
      state_out[k*2  +: 2] = state_in[shifts[k]*2  +: 2];
    end
    return state_out;
  endfunction : prince_shiftrows_32bit

  function automatic logic [63:0] prince_shiftrows_64bit(logic [63:0]      state_in,
                                                         logic [15:0][3:0] shifts );
    logic [63:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 64/4; k++) begin
      state_out[k*4  +: 4] = state_in[shifts[k]*4  +: 4];
    end
    return state_out;
  endfunction : prince_shiftrows_64bit

  // XOR reduction of four nibbles in a 16bit subvector
  function automatic logic [3:0] prince_nibble_red16(logic [15:0] vect);
    return vect[0 +: 4] ^ vect[4 +: 4] ^ vect[8 +: 4] ^ vect[12 +: 4];
  endfunction : prince_nibble_red16

  // M prime multiplication
  function automatic logic [31:0] prince_mult_prime_32bit(logic [31:0] state_in);
    logic [31:0] state_out;
    // M0
    state_out[0  +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST3);
    state_out[4  +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST2);
    state_out[8  +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST1);
    state_out[12 +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST0);
    // M1
    state_out[16 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST0);
    state_out[20 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST3);
    state_out[24 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST2);
    state_out[28 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST1);
    return state_out;
  endfunction : prince_mult_prime_32bit

  // M prime multiplication
  function automatic logic [63:0] prince_mult_prime_64bit(logic [63:0] state_in);
    logic [63:0] state_out;
    // M0
    state_out[0  +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST3);
    state_out[4  +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST2);
    state_out[8  +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST1);
    state_out[12 +: 4] = prince_nibble_red16(state_in[ 0 +: 16] & PRINCE_SHIFT_ROWS_CONST0);
    // M1
    state_out[16 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST0);
    state_out[20 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST3);
    state_out[24 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST2);
    state_out[28 +: 4] = prince_nibble_red16(state_in[16 +: 16] & PRINCE_SHIFT_ROWS_CONST1);
    // M1
    state_out[32 +: 4] = prince_nibble_red16(state_in[32 +: 16] & PRINCE_SHIFT_ROWS_CONST0);
    state_out[36 +: 4] = prince_nibble_red16(state_in[32 +: 16] & PRINCE_SHIFT_ROWS_CONST3);
    state_out[40 +: 4] = prince_nibble_red16(state_in[32 +: 16] & PRINCE_SHIFT_ROWS_CONST2);
    state_out[44 +: 4] = prince_nibble_red16(state_in[32 +: 16] & PRINCE_SHIFT_ROWS_CONST1);
    // M0
    state_out[48 +: 4] = prince_nibble_red16(state_in[48 +: 16] & PRINCE_SHIFT_ROWS_CONST3);
    state_out[52 +: 4] = prince_nibble_red16(state_in[48 +: 16] & PRINCE_SHIFT_ROWS_CONST2);
    state_out[56 +: 4] = prince_nibble_red16(state_in[48 +: 16] & PRINCE_SHIFT_ROWS_CONST1);
    state_out[60 +: 4] = prince_nibble_red16(state_in[48 +: 16] & PRINCE_SHIFT_ROWS_CONST0);
    return state_out;
  endfunction : prince_mult_prime_64bit


  ////////////////////
  // PRESENT Cipher //
  ////////////////////

  // this is the sbox from the present cipher
  parameter logic [15:0][3:0] PRESENT_SBOX4 = {4'h2, 4'h1, 4'h7, 4'h4,
                                               4'h8, 4'hF, 4'hE, 4'h3,
                                               4'hD, 4'hA, 4'h0, 4'h9,
                                               4'hB, 4'h6, 4'h5, 4'hC};

  parameter logic [15:0][3:0] PRESENT_SBOX4_INV = {4'hA, 4'h9, 4'h7, 4'h0,
                                                   4'h3, 4'h6, 4'h4, 4'hB,
                                                   4'hD, 4'h2, 4'h1, 4'hC,
                                                   4'h8, 4'hF, 4'hE, 4'h5};

  // these are modified permutation indices for a 32bit version that
  // follow the same pattern as for the 64bit version
  parameter logic [31:0][4:0] PRESENT_PERM32 = {5'd31, 5'd23, 5'd15, 5'd07,
                                                5'd30, 5'd22, 5'd14, 5'd06,
                                                5'd29, 5'd21, 5'd13, 5'd05,
                                                5'd28, 5'd20, 5'd12, 5'd04,
                                                5'd27, 5'd19, 5'd11, 5'd03,
                                                5'd26, 5'd18, 5'd10, 5'd02,
                                                5'd25, 5'd17, 5'd09, 5'd01,
                                                5'd24, 5'd16, 5'd08, 5'd00};

  parameter logic [31:0][4:0] PRESENT_PERM32_INV = {5'd31, 5'd27, 5'd23, 5'd19,
                                                    5'd15, 5'd11, 5'd07, 5'd03,
                                                    5'd30, 5'd26, 5'd22, 5'd18,
                                                    5'd14, 5'd10, 5'd06, 5'd02,
                                                    5'd29, 5'd25, 5'd21, 5'd17,
                                                    5'd13, 5'd09, 5'd05, 5'd01,
                                                    5'd28, 5'd24, 5'd20, 5'd16,
                                                    5'd12, 5'd08, 5'd04, 5'd00};

  // these are the permutation indices of the present cipher
  parameter logic [63:0][5:0] PRESENT_PERM64 = {6'd63, 6'd47, 6'd31, 6'd15,
                                                6'd62, 6'd46, 6'd30, 6'd14,
                                                6'd61, 6'd45, 6'd29, 6'd13,
                                                6'd60, 6'd44, 6'd28, 6'd12,
                                                6'd59, 6'd43, 6'd27, 6'd11,
                                                6'd58, 6'd42, 6'd26, 6'd10,
                                                6'd57, 6'd41, 6'd25, 6'd09,
                                                6'd56, 6'd40, 6'd24, 6'd08,
                                                6'd55, 6'd39, 6'd23, 6'd07,
                                                6'd54, 6'd38, 6'd22, 6'd06,
                                                6'd53, 6'd37, 6'd21, 6'd05,
                                                6'd52, 6'd36, 6'd20, 6'd04,
                                                6'd51, 6'd35, 6'd19, 6'd03,
                                                6'd50, 6'd34, 6'd18, 6'd02,
                                                6'd49, 6'd33, 6'd17, 6'd01,
                                                6'd48, 6'd32, 6'd16, 6'd00};

  parameter logic [63:0][5:0] PRESENT_PERM64_INV = {6'd63, 6'd59, 6'd55, 6'd51,
                                                    6'd47, 6'd43, 6'd39, 6'd35,
                                                    6'd31, 6'd27, 6'd23, 6'd19,
                                                    6'd15, 6'd11, 6'd07, 6'd03,
                                                    6'd62, 6'd58, 6'd54, 6'd50,
                                                    6'd46, 6'd42, 6'd38, 6'd34,
                                                    6'd30, 6'd26, 6'd22, 6'd18,
                                                    6'd14, 6'd10, 6'd06, 6'd02,
                                                    6'd61, 6'd57, 6'd53, 6'd49,
                                                    6'd45, 6'd41, 6'd37, 6'd33,
                                                    6'd29, 6'd25, 6'd21, 6'd17,
                                                    6'd13, 6'd09, 6'd05, 6'd01,
                                                    6'd60, 6'd56, 6'd52, 6'd48,
                                                    6'd44, 6'd40, 6'd36, 6'd32,
                                                    6'd28, 6'd24, 6'd20, 6'd16,
                                                    6'd12, 6'd08, 6'd04, 6'd00};

  // forward key schedule
  function automatic logic [63:0] present_update_key64(logic [63:0] key_in,
                                                       logic [4:0]  round_idx);
    logic [63:0] key_out;
    // rotate by 61 to the left
    key_out = {key_in[63-61:0], key_in[63:64-61]};
    // sbox on uppermost 4 bits
    key_out[63 -: 4] = PRESENT_SBOX4[key_out[63 -: 4]];
    // xor in round counter on bits 19 to 15
    key_out[19:15] ^= round_idx;
    return key_out;
  endfunction : present_update_key64

  function automatic logic [79:0] present_update_key80(logic [79:0] key_in,
                                                       logic [4:0]  round_idx);
    logic [79:0] key_out;
    // rotate by 61 to the left
    key_out = {key_in[79-61:0], key_in[79:80-61]};
    // sbox on uppermost 4 bits
    key_out[79 -: 4] = PRESENT_SBOX4[key_out[79 -: 4]];
    // xor in round counter on bits 19 to 15
    key_out[19:15] ^= round_idx;
    return key_out;
  endfunction : present_update_key80

  function automatic logic [127:0] present_update_key128(logic [127:0] key_in,
                                                         logic [4:0]   round_idx);
    logic [127:0] key_out;
    // rotate by 61 to the left
    key_out = {key_in[127-61:0], key_in[127:128-61]};
    // sbox on uppermost 4 bits
    key_out[127 -: 4] = PRESENT_SBOX4[key_out[127 -: 4]];
    // sbox on second nibble from top
    key_out[123 -: 4] = PRESENT_SBOX4[key_out[123 -: 4]];
    // xor in round counter on bits 66 to 62
    key_out[66:62] ^= round_idx;
    return key_out;
  endfunction : present_update_key128


  // inverse key schedule
  function automatic logic [63:0] present_inv_update_key64(logic [63:0] key_in,
                                                           logic [4:0]  round_idx);
    logic [63:0] key_out = key_in;
    // xor in round counter on bits 19 to 15
    key_out[19:15] ^= round_idx;
    // sbox on uppermost 4 bits
    key_out[63 -: 4] = PRESENT_SBOX4_INV[key_out[63 -: 4]];
    // rotate by 61 to the right
    key_out = {key_out[60:0], key_out[63:61]};
    return key_out;
  endfunction : present_inv_update_key64

  function automatic logic [79:0] present_inv_update_key80(logic [79:0] key_in,
                                                           logic [4:0]  round_idx);
    logic [79:0] key_out = key_in;
    // xor in round counter on bits 19 to 15
    key_out[19:15] ^= round_idx;
    // sbox on uppermost 4 bits
    key_out[79 -: 4] = PRESENT_SBOX4_INV[key_out[79 -: 4]];
    // rotate by 61 to the right
    key_out = {key_out[60:0], key_out[79:61]};
    return key_out;
  endfunction : present_inv_update_key80

  function automatic logic [127:0] present_inv_update_key128(logic [127:0] key_in,
                                                             logic [4:0]   round_idx);
    logic [127:0] key_out = key_in;
    // xor in round counter on bits 66 to 62
    key_out[66:62] ^= round_idx;
    // sbox on second highest nibble
    key_out[123 -: 4] = PRESENT_SBOX4_INV[key_out[123 -: 4]];
    // sbox on uppermost 4 bits
    key_out[127 -: 4] = PRESENT_SBOX4_INV[key_out[127 -: 4]];
    // rotate by 61 to the right
    key_out = {key_out[60:0], key_out[127:61]};
    return key_out;
  endfunction : present_inv_update_key128


  // these functions can be used to derive the DEC key from the ENC key by
  // stepping the key by the correct number of rounds using the keyschedule functions above.
  function automatic logic [63:0] present_get_dec_key64(logic [63:0] key_in,
                                                        // total number of rounds employed
                                                        logic [4:0]  round_cnt);
    logic [63:0] key_out;
    key_out = key_in;
    for (int unsigned k = 0; k < round_cnt; k++) begin
      key_out = present_update_key64(key_out, 5'(k + 1));
    end
    return key_out;
  endfunction : present_get_dec_key64

  function automatic logic [79:0] present_get_dec_key80(logic [79:0] key_in,
                                                        // total number of rounds employed
                                                        logic [4:0]  round_cnt);
    logic [79:0] key_out;
    key_out = key_in;
    for (int unsigned k = 0; k < round_cnt; k++) begin
      key_out = present_update_key80(key_out, 5'(k + 1));
    end
    return key_out;
  endfunction : present_get_dec_key80

  function automatic logic [127:0] present_get_dec_key128(logic [127:0] key_in,
                                                          // total number of rounds employed
                                                          logic [4:0]   round_cnt);
    logic [127:0] key_out;
    key_out = key_in;
    for (int unsigned k = 0; k < round_cnt; k++) begin
      key_out = present_update_key128(key_out, 5'(k + 1));
    end
    return key_out;
  endfunction : present_get_dec_key128

  /////////////////////////
  // Common Subfunctions //
  /////////////////////////

  function automatic logic [7:0] sbox4_8bit(logic [7:0] state_in, logic [15:0][3:0] sbox4);
    logic [7:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 8/4; k++) begin
      state_out[k*4  +: 4] = sbox4[state_in[k*4  +: 4]];
    end
    return state_out;
  endfunction : sbox4_8bit

  function automatic logic [15:0] sbox4_16bit(logic [15:0] state_in, logic [15:0][3:0] sbox4);
    logic [15:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 2; k++) begin
      state_out[k*8  +: 8] = sbox4_8bit(state_in[k*8  +: 8], sbox4);
    end
    return state_out;
  endfunction : sbox4_16bit

  function automatic logic [31:0] sbox4_32bit(logic [31:0] state_in, logic [15:0][3:0] sbox4);
    logic [31:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 4; k++) begin
      state_out[k*8  +: 8] = sbox4_8bit(state_in[k*8  +: 8], sbox4);
    end
    return state_out;
  endfunction : sbox4_32bit

  function automatic logic [63:0] sbox4_64bit(logic [63:0] state_in, logic [15:0][3:0] sbox4);
    logic [63:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 8; k++) begin
      state_out[k*8  +: 8] = sbox4_8bit(state_in[k*8  +: 8], sbox4);
    end
    return state_out;
  endfunction : sbox4_64bit

  function automatic logic [7:0] perm_8bit(logic [7:0] state_in, logic [7:0][2:0] perm);
    logic [7:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 8; k++) begin
      state_out[perm[k]] = state_in[k];
    end
    return state_out;
  endfunction : perm_8bit

    function automatic logic [15:0] perm_16bit(logic [15:0] state_in, logic [15:0][3:0] perm);
    logic [15:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 16; k++) begin
      state_out[perm[k]] = state_in[k];
    end
    return state_out;
  endfunction : perm_16bit

  function automatic logic [31:0] perm_32bit(logic [31:0] state_in, logic [31:0][4:0] perm);
    logic [31:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 32; k++) begin
      state_out[perm[k]] = state_in[k];
    end
    return state_out;
  endfunction : perm_32bit

  function automatic logic [63:0] perm_64bit(logic [63:0] state_in, logic [63:0][5:0] perm);
    logic [63:0] state_out;
    // note that if simulation performance becomes an issue, this loop can be unrolled
    for (int k = 0; k < 64; k++) begin
      state_out[perm[k]] = state_in[k];
    end
    return state_out;
  endfunction : perm_64bit

endpackage : prim_cipher_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// CRC32 calculator
//
// This module takes in n-bits data words (n defined by BytePerWord parameter) and updates an
// internally stored CRC with each valid data word. The polynomial used is the standard CRC32 IEEE
// one. An interface is provided to set the internal CRC to an arbitrary value. The output CRC is an
// inverted version of the internally stored CRC and the input CRC is inverted before being stored.
// This is done so results match existing widely used software libraries (e.g. the crc32
// functionality available in Python). Note that a initial CRC of 0x0 (corresponding to an internal
// CRC of 0xffffffff) must be used to match results generated elsewhere.


module prim_crc32 #(
  parameter int unsigned BytesPerWord = 4
) (
  input  logic                      clk_i,
  input  logic                      rst_ni,

  input  logic                      set_crc_i,
  input  logic [31:0]               crc_in_i,

  input  logic                      data_valid_i,
  input  logic [BytesPerWord*8-1:0] data_i,

  output logic [31:0]               crc_out_o
);
  // Generated using hw/ip/prim/util/prim_crc32_table_gen.py
  function automatic logic [31:0] crc32_byte_calc(logic [7:0] b);
    unique case (b)
      8'hff:   crc32_byte_calc = 32'h2d02ef8d;
      8'hfe:   crc32_byte_calc = 32'h5a05df1b;
      8'hfd:   crc32_byte_calc = 32'hc30c8ea1;
      8'hfc:   crc32_byte_calc = 32'hb40bbe37;
      8'hfb:   crc32_byte_calc = 32'h2a6f2b94;
      8'hfa:   crc32_byte_calc = 32'h5d681b02;
      8'hf9:   crc32_byte_calc = 32'hc4614ab8;
      8'hf8:   crc32_byte_calc = 32'hb3667a2e;
      8'hf7:   crc32_byte_calc = 32'h23d967bf;
      8'hf6:   crc32_byte_calc = 32'h54de5729;
      8'hf5:   crc32_byte_calc = 32'hcdd70693;
      8'hf4:   crc32_byte_calc = 32'hbad03605;
      8'hf3:   crc32_byte_calc = 32'h24b4a3a6;
      8'hf2:   crc32_byte_calc = 32'h53b39330;
      8'hf1:   crc32_byte_calc = 32'hcabac28a;
      8'hf0:   crc32_byte_calc = 32'hbdbdf21c;
      8'hef:   crc32_byte_calc = 32'h30b5ffe9;
      8'hee:   crc32_byte_calc = 32'h47b2cf7f;
      8'hed:   crc32_byte_calc = 32'hdebb9ec5;
      8'hec:   crc32_byte_calc = 32'ha9bcae53;
      8'heb:   crc32_byte_calc = 32'h37d83bf0;
      8'hea:   crc32_byte_calc = 32'h40df0b66;
      8'he9:   crc32_byte_calc = 32'hd9d65adc;
      8'he8:   crc32_byte_calc = 32'haed16a4a;
      8'he7:   crc32_byte_calc = 32'h3e6e77db;
      8'he6:   crc32_byte_calc = 32'h4969474d;
      8'he5:   crc32_byte_calc = 32'hd06016f7;
      8'he4:   crc32_byte_calc = 32'ha7672661;
      8'he3:   crc32_byte_calc = 32'h3903b3c2;
      8'he2:   crc32_byte_calc = 32'h4e048354;
      8'he1:   crc32_byte_calc = 32'hd70dd2ee;
      8'he0:   crc32_byte_calc = 32'ha00ae278;
      8'hdf:   crc32_byte_calc = 32'h166ccf45;
      8'hde:   crc32_byte_calc = 32'h616bffd3;
      8'hdd:   crc32_byte_calc = 32'hf862ae69;
      8'hdc:   crc32_byte_calc = 32'h8f659eff;
      8'hdb:   crc32_byte_calc = 32'h11010b5c;
      8'hda:   crc32_byte_calc = 32'h66063bca;
      8'hd9:   crc32_byte_calc = 32'hff0f6a70;
      8'hd8:   crc32_byte_calc = 32'h88085ae6;
      8'hd7:   crc32_byte_calc = 32'h18b74777;
      8'hd6:   crc32_byte_calc = 32'h6fb077e1;
      8'hd5:   crc32_byte_calc = 32'hf6b9265b;
      8'hd4:   crc32_byte_calc = 32'h81be16cd;
      8'hd3:   crc32_byte_calc = 32'h1fda836e;
      8'hd2:   crc32_byte_calc = 32'h68ddb3f8;
      8'hd1:   crc32_byte_calc = 32'hf1d4e242;
      8'hd0:   crc32_byte_calc = 32'h86d3d2d4;
      8'hcf:   crc32_byte_calc = 32'h0bdbdf21;
      8'hce:   crc32_byte_calc = 32'h7cdcefb7;
      8'hcd:   crc32_byte_calc = 32'he5d5be0d;
      8'hcc:   crc32_byte_calc = 32'h92d28e9b;
      8'hcb:   crc32_byte_calc = 32'h0cb61b38;
      8'hca:   crc32_byte_calc = 32'h7bb12bae;
      8'hc9:   crc32_byte_calc = 32'he2b87a14;
      8'hc8:   crc32_byte_calc = 32'h95bf4a82;
      8'hc7:   crc32_byte_calc = 32'h05005713;
      8'hc6:   crc32_byte_calc = 32'h72076785;
      8'hc5:   crc32_byte_calc = 32'heb0e363f;
      8'hc4:   crc32_byte_calc = 32'h9c0906a9;
      8'hc3:   crc32_byte_calc = 32'h026d930a;
      8'hc2:   crc32_byte_calc = 32'h756aa39c;
      8'hc1:   crc32_byte_calc = 32'hec63f226;
      8'hc0:   crc32_byte_calc = 32'h9b64c2b0;
      8'hbf:   crc32_byte_calc = 32'h5bdeae1d;
      8'hbe:   crc32_byte_calc = 32'h2cd99e8b;
      8'hbd:   crc32_byte_calc = 32'hb5d0cf31;
      8'hbc:   crc32_byte_calc = 32'hc2d7ffa7;
      8'hbb:   crc32_byte_calc = 32'h5cb36a04;
      8'hba:   crc32_byte_calc = 32'h2bb45a92;
      8'hb9:   crc32_byte_calc = 32'hb2bd0b28;
      8'hb8:   crc32_byte_calc = 32'hc5ba3bbe;
      8'hb7:   crc32_byte_calc = 32'h5505262f;
      8'hb6:   crc32_byte_calc = 32'h220216b9;
      8'hb5:   crc32_byte_calc = 32'hbb0b4703;
      8'hb4:   crc32_byte_calc = 32'hcc0c7795;
      8'hb3:   crc32_byte_calc = 32'h5268e236;
      8'hb2:   crc32_byte_calc = 32'h256fd2a0;
      8'hb1:   crc32_byte_calc = 32'hbc66831a;
      8'hb0:   crc32_byte_calc = 32'hcb61b38c;
      8'haf:   crc32_byte_calc = 32'h4669be79;
      8'hae:   crc32_byte_calc = 32'h316e8eef;
      8'had:   crc32_byte_calc = 32'ha867df55;
      8'hac:   crc32_byte_calc = 32'hdf60efc3;
      8'hab:   crc32_byte_calc = 32'h41047a60;
      8'haa:   crc32_byte_calc = 32'h36034af6;
      8'ha9:   crc32_byte_calc = 32'haf0a1b4c;
      8'ha8:   crc32_byte_calc = 32'hd80d2bda;
      8'ha7:   crc32_byte_calc = 32'h48b2364b;
      8'ha6:   crc32_byte_calc = 32'h3fb506dd;
      8'ha5:   crc32_byte_calc = 32'ha6bc5767;
      8'ha4:   crc32_byte_calc = 32'hd1bb67f1;
      8'ha3:   crc32_byte_calc = 32'h4fdff252;
      8'ha2:   crc32_byte_calc = 32'h38d8c2c4;
      8'ha1:   crc32_byte_calc = 32'ha1d1937e;
      8'ha0:   crc32_byte_calc = 32'hd6d6a3e8;
      8'h9f:   crc32_byte_calc = 32'h60b08ed5;
      8'h9e:   crc32_byte_calc = 32'h17b7be43;
      8'h9d:   crc32_byte_calc = 32'h8ebeeff9;
      8'h9c:   crc32_byte_calc = 32'hf9b9df6f;
      8'h9b:   crc32_byte_calc = 32'h67dd4acc;
      8'h9a:   crc32_byte_calc = 32'h10da7a5a;
      8'h99:   crc32_byte_calc = 32'h89d32be0;
      8'h98:   crc32_byte_calc = 32'hfed41b76;
      8'h97:   crc32_byte_calc = 32'h6e6b06e7;
      8'h96:   crc32_byte_calc = 32'h196c3671;
      8'h95:   crc32_byte_calc = 32'h806567cb;
      8'h94:   crc32_byte_calc = 32'hf762575d;
      8'h93:   crc32_byte_calc = 32'h6906c2fe;
      8'h92:   crc32_byte_calc = 32'h1e01f268;
      8'h91:   crc32_byte_calc = 32'h8708a3d2;
      8'h90:   crc32_byte_calc = 32'hf00f9344;
      8'h8f:   crc32_byte_calc = 32'h7d079eb1;
      8'h8e:   crc32_byte_calc = 32'h0a00ae27;
      8'h8d:   crc32_byte_calc = 32'h9309ff9d;
      8'h8c:   crc32_byte_calc = 32'he40ecf0b;
      8'h8b:   crc32_byte_calc = 32'h7a6a5aa8;
      8'h8a:   crc32_byte_calc = 32'h0d6d6a3e;
      8'h89:   crc32_byte_calc = 32'h94643b84;
      8'h88:   crc32_byte_calc = 32'he3630b12;
      8'h87:   crc32_byte_calc = 32'h73dc1683;
      8'h86:   crc32_byte_calc = 32'h04db2615;
      8'h85:   crc32_byte_calc = 32'h9dd277af;
      8'h84:   crc32_byte_calc = 32'head54739;
      8'h83:   crc32_byte_calc = 32'h74b1d29a;
      8'h82:   crc32_byte_calc = 32'h03b6e20c;
      8'h81:   crc32_byte_calc = 32'h9abfb3b6;
      8'h80:   crc32_byte_calc = 32'hedb88320;
      8'h7f:   crc32_byte_calc = 32'hc0ba6cad;
      8'h7e:   crc32_byte_calc = 32'hb7bd5c3b;
      8'h7d:   crc32_byte_calc = 32'h2eb40d81;
      8'h7c:   crc32_byte_calc = 32'h59b33d17;
      8'h7b:   crc32_byte_calc = 32'hc7d7a8b4;
      8'h7a:   crc32_byte_calc = 32'hb0d09822;
      8'h79:   crc32_byte_calc = 32'h29d9c998;
      8'h78:   crc32_byte_calc = 32'h5edef90e;
      8'h77:   crc32_byte_calc = 32'hce61e49f;
      8'h76:   crc32_byte_calc = 32'hb966d409;
      8'h75:   crc32_byte_calc = 32'h206f85b3;
      8'h74:   crc32_byte_calc = 32'h5768b525;
      8'h73:   crc32_byte_calc = 32'hc90c2086;
      8'h72:   crc32_byte_calc = 32'hbe0b1010;
      8'h71:   crc32_byte_calc = 32'h270241aa;
      8'h70:   crc32_byte_calc = 32'h5005713c;
      8'h6f:   crc32_byte_calc = 32'hdd0d7cc9;
      8'h6e:   crc32_byte_calc = 32'haa0a4c5f;
      8'h6d:   crc32_byte_calc = 32'h33031de5;
      8'h6c:   crc32_byte_calc = 32'h44042d73;
      8'h6b:   crc32_byte_calc = 32'hda60b8d0;
      8'h6a:   crc32_byte_calc = 32'had678846;
      8'h69:   crc32_byte_calc = 32'h346ed9fc;
      8'h68:   crc32_byte_calc = 32'h4369e96a;
      8'h67:   crc32_byte_calc = 32'hd3d6f4fb;
      8'h66:   crc32_byte_calc = 32'ha4d1c46d;
      8'h65:   crc32_byte_calc = 32'h3dd895d7;
      8'h64:   crc32_byte_calc = 32'h4adfa541;
      8'h63:   crc32_byte_calc = 32'hd4bb30e2;
      8'h62:   crc32_byte_calc = 32'ha3bc0074;
      8'h61:   crc32_byte_calc = 32'h3ab551ce;
      8'h60:   crc32_byte_calc = 32'h4db26158;
      8'h5f:   crc32_byte_calc = 32'hfbd44c65;
      8'h5e:   crc32_byte_calc = 32'h8cd37cf3;
      8'h5d:   crc32_byte_calc = 32'h15da2d49;
      8'h5c:   crc32_byte_calc = 32'h62dd1ddf;
      8'h5b:   crc32_byte_calc = 32'hfcb9887c;
      8'h5a:   crc32_byte_calc = 32'h8bbeb8ea;
      8'h59:   crc32_byte_calc = 32'h12b7e950;
      8'h58:   crc32_byte_calc = 32'h65b0d9c6;
      8'h57:   crc32_byte_calc = 32'hf50fc457;
      8'h56:   crc32_byte_calc = 32'h8208f4c1;
      8'h55:   crc32_byte_calc = 32'h1b01a57b;
      8'h54:   crc32_byte_calc = 32'h6c0695ed;
      8'h53:   crc32_byte_calc = 32'hf262004e;
      8'h52:   crc32_byte_calc = 32'h856530d8;
      8'h51:   crc32_byte_calc = 32'h1c6c6162;
      8'h50:   crc32_byte_calc = 32'h6b6b51f4;
      8'h4f:   crc32_byte_calc = 32'he6635c01;
      8'h4e:   crc32_byte_calc = 32'h91646c97;
      8'h4d:   crc32_byte_calc = 32'h086d3d2d;
      8'h4c:   crc32_byte_calc = 32'h7f6a0dbb;
      8'h4b:   crc32_byte_calc = 32'he10e9818;
      8'h4a:   crc32_byte_calc = 32'h9609a88e;
      8'h49:   crc32_byte_calc = 32'h0f00f934;
      8'h48:   crc32_byte_calc = 32'h7807c9a2;
      8'h47:   crc32_byte_calc = 32'he8b8d433;
      8'h46:   crc32_byte_calc = 32'h9fbfe4a5;
      8'h45:   crc32_byte_calc = 32'h06b6b51f;
      8'h44:   crc32_byte_calc = 32'h71b18589;
      8'h43:   crc32_byte_calc = 32'hefd5102a;
      8'h42:   crc32_byte_calc = 32'h98d220bc;
      8'h41:   crc32_byte_calc = 32'h01db7106;
      8'h40:   crc32_byte_calc = 32'h76dc4190;
      8'h3f:   crc32_byte_calc = 32'hb6662d3d;
      8'h3e:   crc32_byte_calc = 32'hc1611dab;
      8'h3d:   crc32_byte_calc = 32'h58684c11;
      8'h3c:   crc32_byte_calc = 32'h2f6f7c87;
      8'h3b:   crc32_byte_calc = 32'hb10be924;
      8'h3a:   crc32_byte_calc = 32'hc60cd9b2;
      8'h39:   crc32_byte_calc = 32'h5f058808;
      8'h38:   crc32_byte_calc = 32'h2802b89e;
      8'h37:   crc32_byte_calc = 32'hb8bda50f;
      8'h36:   crc32_byte_calc = 32'hcfba9599;
      8'h35:   crc32_byte_calc = 32'h56b3c423;
      8'h34:   crc32_byte_calc = 32'h21b4f4b5;
      8'h33:   crc32_byte_calc = 32'hbfd06116;
      8'h32:   crc32_byte_calc = 32'hc8d75180;
      8'h31:   crc32_byte_calc = 32'h51de003a;
      8'h30:   crc32_byte_calc = 32'h26d930ac;
      8'h2f:   crc32_byte_calc = 32'habd13d59;
      8'h2e:   crc32_byte_calc = 32'hdcd60dcf;
      8'h2d:   crc32_byte_calc = 32'h45df5c75;
      8'h2c:   crc32_byte_calc = 32'h32d86ce3;
      8'h2b:   crc32_byte_calc = 32'hacbcf940;
      8'h2a:   crc32_byte_calc = 32'hdbbbc9d6;
      8'h29:   crc32_byte_calc = 32'h42b2986c;
      8'h28:   crc32_byte_calc = 32'h35b5a8fa;
      8'h27:   crc32_byte_calc = 32'ha50ab56b;
      8'h26:   crc32_byte_calc = 32'hd20d85fd;
      8'h25:   crc32_byte_calc = 32'h4b04d447;
      8'h24:   crc32_byte_calc = 32'h3c03e4d1;
      8'h23:   crc32_byte_calc = 32'ha2677172;
      8'h22:   crc32_byte_calc = 32'hd56041e4;
      8'h21:   crc32_byte_calc = 32'h4c69105e;
      8'h20:   crc32_byte_calc = 32'h3b6e20c8;
      8'h1f:   crc32_byte_calc = 32'h8d080df5;
      8'h1e:   crc32_byte_calc = 32'hfa0f3d63;
      8'h1d:   crc32_byte_calc = 32'h63066cd9;
      8'h1c:   crc32_byte_calc = 32'h14015c4f;
      8'h1b:   crc32_byte_calc = 32'h8a65c9ec;
      8'h1a:   crc32_byte_calc = 32'hfd62f97a;
      8'h19:   crc32_byte_calc = 32'h646ba8c0;
      8'h18:   crc32_byte_calc = 32'h136c9856;
      8'h17:   crc32_byte_calc = 32'h83d385c7;
      8'h16:   crc32_byte_calc = 32'hf4d4b551;
      8'h15:   crc32_byte_calc = 32'h6ddde4eb;
      8'h14:   crc32_byte_calc = 32'h1adad47d;
      8'h13:   crc32_byte_calc = 32'h84be41de;
      8'h12:   crc32_byte_calc = 32'hf3b97148;
      8'h11:   crc32_byte_calc = 32'h6ab020f2;
      8'h10:   crc32_byte_calc = 32'h1db71064;
      8'h0f:   crc32_byte_calc = 32'h90bf1d91;
      8'h0e:   crc32_byte_calc = 32'he7b82d07;
      8'h0d:   crc32_byte_calc = 32'h7eb17cbd;
      8'h0c:   crc32_byte_calc = 32'h09b64c2b;
      8'h0b:   crc32_byte_calc = 32'h97d2d988;
      8'h0a:   crc32_byte_calc = 32'he0d5e91e;
      8'h09:   crc32_byte_calc = 32'h79dcb8a4;
      8'h08:   crc32_byte_calc = 32'h0edb8832;
      8'h07:   crc32_byte_calc = 32'h9e6495a3;
      8'h06:   crc32_byte_calc = 32'he963a535;
      8'h05:   crc32_byte_calc = 32'h706af48f;
      8'h04:   crc32_byte_calc = 32'h076dc419;
      8'h03:   crc32_byte_calc = 32'h990951ba;
      8'h02:   crc32_byte_calc = 32'hee0e612c;
      8'h01:   crc32_byte_calc = 32'h77073096;
      8'h00:   crc32_byte_calc = 32'h00000000;
      default: crc32_byte_calc = '0;
    endcase
  endfunction

  logic [31:0] crc_d, crc_q;
  logic        crc_en;
  logic [31:0] crc_stages[BytesPerWord + 1];

  assign crc_en = set_crc_i | data_valid_i;

  assign crc_stages[0] = crc_q;

  for (genvar i = 0;i < BytesPerWord; ++i) begin : g_crc_stages
    assign crc_stages[i + 1] =
      {8'h00, crc_stages[i][31:8]} ^
      crc32_byte_calc(crc_stages[i][7:0] ^ data_i[i * 8 +: 8]);
  end

  always_comb begin
    if (set_crc_i) begin
      crc_d = ~crc_in_i;
    end else begin
      crc_d = crc_stages[BytesPerWord];
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      crc_q <= 32'hFFFFFFFF;
    end else if (crc_en) begin
      crc_q <= crc_d;
    end
  end

  assign crc_out_o = ~crc_q;
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_and2 #(
  parameter int Width = 1
) (
  input        [Width-1:0] in0_i,
  input        [Width-1:0] in1_i,
  output logic [Width-1:0] out_o
);

  assign out_o = in0_i & in1_i;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_buf #(
  parameter int Width = 1
) (
  input        [Width-1:0] in_i,
  output logic [Width-1:0] out_o
);

  logic [Width-1:0] inv;
  assign inv = ~in_i;
  assign out_o = ~inv;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_flop #(
  parameter int               Width      = 1,
  parameter logic [Width-1:0] ResetValue = 0
) (
  input                    clk_i,
  input                    rst_ni,
  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_o
);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      q_o <= ResetValue;
    end else begin
      q_o <= d_i;
    end
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_xnor2 #(
  parameter int Width = 1
) (
  input        [Width-1:0] in0_i,
  input        [Width-1:0] in1_i,
  output logic [Width-1:0] out_o
);

  assign out_o = !(in0_i ^ in1_i);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_xor2 #(
  parameter int Width = 1
) (
  input        [Width-1:0] in0_i,
  input        [Width-1:0] in1_i,
  output logic [Width-1:0] out_o
);

  assign out_o = in0_i ^ in1_i;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package prim_pad_wrapper_pkg;

  typedef enum logic [2:0] {
    BidirStd = 3'h0,     // Standard bidirectional pad
    BidirTol = 3'h1,     // Voltage tolerant pad
    BidirOd = 3'h2,      // Open-drain capable pad
    InputStd = 3'h3,     // Input-only pad
    AnalogIn0 = 3'h4,    // Analog input pad
    AnalogIn1 = 3'h5,    // Analog input pad
    DualBidirTol = 3'h6  // Dual Voltage tolerant pad
  } pad_type_e;

  typedef enum logic [1:0] {
    NoScan = 2'h0,
    ScanIn = 2'h1,
    ScanOut = 2'h2
  } scan_role_e;

  // Pad attributes
  parameter int DriveStrDw = 4;
  parameter int SlewRateDw = 2;

  typedef struct packed {
    logic [DriveStrDw-1:0] drive_strength; // Drive strength (0000: weakest, 1111: strongest).
    logic [SlewRateDw-1:0] slew_rate;      // Slew rate (0: slowest, 11: fastest).
    logic od_en;                           // Open-drain enable
    logic schmitt_en;                      // Schmitt trigger enable.
    logic keep_en;                         // Keeper enable.
    logic pull_select;                     // Pull direction (0: pull down, 1: pull up).
    logic pull_en;                         // Pull enable.
    logic virt_od_en;                      // Virtual open drain enable.
    logic invert;                          // Input/output inversion.
  } pad_attr_t;

  parameter int AttrDw = $bits(pad_attr_t);

  // Power OK signals (library dependent)
  parameter int PokDw = 8;

  typedef logic [PokDw-1:0] pad_pok_t;

endpackage : prim_pad_wrapper_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED package generated by
// util/design/secded_gen.py from util/design/data/secded_cfg.hjson

package prim_secded_pkg;

  typedef enum int {
    SecdedNone,
    Secded_22_16,
    Secded_28_22,
    Secded_39_32,
    Secded_64_57,
    Secded_72_64,
    SecdedHamming_22_16,
    SecdedHamming_39_32,
    SecdedHamming_72_64,
    SecdedHamming_76_68,
    SecdedInv_22_16,
    SecdedInv_28_22,
    SecdedInv_39_32,
    SecdedInv_64_57,
    SecdedInv_72_64,
    SecdedInvHamming_22_16,
    SecdedInvHamming_39_32,
    SecdedInvHamming_72_64,
    SecdedInvHamming_76_68
  } prim_secded_e;

  function automatic int get_ecc_data_width(prim_secded_e ecc_type);
    case (ecc_type)
      Secded_22_16: return 16;
      Secded_28_22: return 22;
      Secded_39_32: return 32;
      Secded_64_57: return 57;
      Secded_72_64: return 64;
      SecdedHamming_22_16: return 16;
      SecdedHamming_39_32: return 32;
      SecdedHamming_72_64: return 64;
      SecdedHamming_76_68: return 68;
      SecdedInv_22_16: return 16;
      SecdedInv_28_22: return 22;
      SecdedInv_39_32: return 32;
      SecdedInv_64_57: return 57;
      SecdedInv_72_64: return 64;
      SecdedInvHamming_22_16: return 16;
      SecdedInvHamming_39_32: return 32;
      SecdedInvHamming_72_64: return 64;
      SecdedInvHamming_76_68: return 68;
      // Return a non-zero width to avoid VCS compile issues
      default: return 32;
    endcase
  endfunction

  function automatic int get_ecc_parity_width(prim_secded_e ecc_type);
    case (ecc_type)
      Secded_22_16: return 6;
      Secded_28_22: return 6;
      Secded_39_32: return 7;
      Secded_64_57: return 7;
      Secded_72_64: return 8;
      SecdedHamming_22_16: return 6;
      SecdedHamming_39_32: return 7;
      SecdedHamming_72_64: return 8;
      SecdedHamming_76_68: return 8;
      SecdedInv_22_16: return 6;
      SecdedInv_28_22: return 6;
      SecdedInv_39_32: return 7;
      SecdedInv_64_57: return 7;
      SecdedInv_72_64: return 8;
      SecdedInvHamming_22_16: return 6;
      SecdedInvHamming_39_32: return 7;
      SecdedInvHamming_72_64: return 8;
      SecdedInvHamming_76_68: return 8;
      default: return 0;
    endcase
  endfunction

  parameter logic [5:0] Secded2216ZeroEcc = 6'h0;
  parameter logic [21:0] Secded2216ZeroWord = 22'h0;

  typedef struct packed {
    logic [15:0] data;
    logic [5:0] syndrome;
    logic [1:0]  err;
  } secded_22_16_t;

  parameter logic [5:0] Secded2822ZeroEcc = 6'h0;
  parameter logic [27:0] Secded2822ZeroWord = 28'h0;

  typedef struct packed {
    logic [21:0] data;
    logic [5:0] syndrome;
    logic [1:0]  err;
  } secded_28_22_t;

  parameter logic [6:0] Secded3932ZeroEcc = 7'h0;
  parameter logic [38:0] Secded3932ZeroWord = 39'h0;

  typedef struct packed {
    logic [31:0] data;
    logic [6:0] syndrome;
    logic [1:0]  err;
  } secded_39_32_t;

  parameter logic [6:0] Secded6457ZeroEcc = 7'h0;
  parameter logic [63:0] Secded6457ZeroWord = 64'h0;

  typedef struct packed {
    logic [56:0] data;
    logic [6:0] syndrome;
    logic [1:0]  err;
  } secded_64_57_t;

  parameter logic [7:0] Secded7264ZeroEcc = 8'h0;
  parameter logic [71:0] Secded7264ZeroWord = 72'h0;

  typedef struct packed {
    logic [63:0] data;
    logic [7:0] syndrome;
    logic [1:0]  err;
  } secded_72_64_t;

  parameter logic [5:0] SecdedHamming2216ZeroEcc = 6'h0;
  parameter logic [21:0] SecdedHamming2216ZeroWord = 22'h0;

  typedef struct packed {
    logic [15:0] data;
    logic [5:0] syndrome;
    logic [1:0]  err;
  } secded_hamming_22_16_t;

  parameter logic [6:0] SecdedHamming3932ZeroEcc = 7'h0;
  parameter logic [38:0] SecdedHamming3932ZeroWord = 39'h0;

  typedef struct packed {
    logic [31:0] data;
    logic [6:0] syndrome;
    logic [1:0]  err;
  } secded_hamming_39_32_t;

  parameter logic [7:0] SecdedHamming7264ZeroEcc = 8'h0;
  parameter logic [71:0] SecdedHamming7264ZeroWord = 72'h0;

  typedef struct packed {
    logic [63:0] data;
    logic [7:0] syndrome;
    logic [1:0]  err;
  } secded_hamming_72_64_t;

  parameter logic [7:0] SecdedHamming7668ZeroEcc = 8'h0;
  parameter logic [75:0] SecdedHamming7668ZeroWord = 76'h0;

  typedef struct packed {
    logic [67:0] data;
    logic [7:0] syndrome;
    logic [1:0]  err;
  } secded_hamming_76_68_t;

  parameter logic [5:0] SecdedInv2216ZeroEcc = 6'h2A;
  parameter logic [21:0] SecdedInv2216ZeroWord = 22'h2A0000;

  typedef struct packed {
    logic [15:0] data;
    logic [5:0] syndrome;
    logic [1:0]  err;
  } secded_inv_22_16_t;

  parameter logic [5:0] SecdedInv2822ZeroEcc = 6'h2A;
  parameter logic [27:0] SecdedInv2822ZeroWord = 28'hA800000;

  typedef struct packed {
    logic [21:0] data;
    logic [5:0] syndrome;
    logic [1:0]  err;
  } secded_inv_28_22_t;

  parameter logic [6:0] SecdedInv3932ZeroEcc = 7'h2A;
  parameter logic [38:0] SecdedInv3932ZeroWord = 39'h2A00000000;

  typedef struct packed {
    logic [31:0] data;
    logic [6:0] syndrome;
    logic [1:0]  err;
  } secded_inv_39_32_t;

  parameter logic [6:0] SecdedInv6457ZeroEcc = 7'h2A;
  parameter logic [63:0] SecdedInv6457ZeroWord = 64'h5400000000000000;

  typedef struct packed {
    logic [56:0] data;
    logic [6:0] syndrome;
    logic [1:0]  err;
  } secded_inv_64_57_t;

  parameter logic [7:0] SecdedInv7264ZeroEcc = 8'hAA;
  parameter logic [71:0] SecdedInv7264ZeroWord = 72'hAA0000000000000000;

  typedef struct packed {
    logic [63:0] data;
    logic [7:0] syndrome;
    logic [1:0]  err;
  } secded_inv_72_64_t;

  parameter logic [5:0] SecdedInvHamming2216ZeroEcc = 6'h2A;
  parameter logic [21:0] SecdedInvHamming2216ZeroWord = 22'h2A0000;

  typedef struct packed {
    logic [15:0] data;
    logic [5:0] syndrome;
    logic [1:0]  err;
  } secded_inv_hamming_22_16_t;

  parameter logic [6:0] SecdedInvHamming3932ZeroEcc = 7'h2A;
  parameter logic [38:0] SecdedInvHamming3932ZeroWord = 39'h2A00000000;

  typedef struct packed {
    logic [31:0] data;
    logic [6:0] syndrome;
    logic [1:0]  err;
  } secded_inv_hamming_39_32_t;

  parameter logic [7:0] SecdedInvHamming7264ZeroEcc = 8'hAA;
  parameter logic [71:0] SecdedInvHamming7264ZeroWord = 72'hAA0000000000000000;

  typedef struct packed {
    logic [63:0] data;
    logic [7:0] syndrome;
    logic [1:0]  err;
  } secded_inv_hamming_72_64_t;

  parameter logic [7:0] SecdedInvHamming7668ZeroEcc = 8'hAA;
  parameter logic [75:0] SecdedInvHamming7668ZeroWord = 76'hAA00000000000000000;

  typedef struct packed {
    logic [67:0] data;
    logic [7:0] syndrome;
    logic [1:0]  err;
  } secded_inv_hamming_76_68_t;

  function automatic logic [21:0]
      prim_secded_22_16_enc (logic [15:0] data_i);
    logic [21:0] data_o;
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00496E);
    data_o[17] = ^(data_o & 22'h00F20B);
    data_o[18] = ^(data_o & 22'h008ED8);
    data_o[19] = ^(data_o & 22'h007714);
    data_o[20] = ^(data_o & 22'h00ACA5);
    data_o[21] = ^(data_o & 22'h0011F3);
    return data_o;
  endfunction

  function automatic secded_22_16_t
      prim_secded_22_16_dec (logic [21:0] data_i);
    logic [15:0] data_o;
    logic [5:0] syndrome_o;
    logic [1:0]  err_o;

    secded_22_16_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 22'h01496E);
    syndrome_o[1] = ^(data_i & 22'h02F20B);
    syndrome_o[2] = ^(data_i & 22'h048ED8);
    syndrome_o[3] = ^(data_i & 22'h087714);
    syndrome_o[4] = ^(data_i & 22'h10ACA5);
    syndrome_o[5] = ^(data_i & 22'h2011F3);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h32) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h23) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h19) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h7) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h2c) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h31) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h34) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'he) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h1c) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h15) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h2a) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'hb) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h16) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [27:0]
      prim_secded_28_22_enc (logic [21:0] data_i);
    logic [27:0] data_o;
    data_o = 28'(data_i);
    data_o[22] = ^(data_o & 28'h03003FF);
    data_o[23] = ^(data_o & 28'h010FC0F);
    data_o[24] = ^(data_o & 28'h0271C71);
    data_o[25] = ^(data_o & 28'h03B6592);
    data_o[26] = ^(data_o & 28'h03DAAA4);
    data_o[27] = ^(data_o & 28'h03ED348);
    return data_o;
  endfunction

  function automatic secded_28_22_t
      prim_secded_28_22_dec (logic [27:0] data_i);
    logic [21:0] data_o;
    logic [5:0] syndrome_o;
    logic [1:0]  err_o;

    secded_28_22_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 28'h07003FF);
    syndrome_o[1] = ^(data_i & 28'h090FC0F);
    syndrome_o[2] = ^(data_i & 28'h1271C71);
    syndrome_o[3] = ^(data_i & 28'h23B6592);
    syndrome_o[4] = ^(data_i & 28'h43DAAA4);
    syndrome_o[5] = ^(data_i & 28'h83ED348);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'hd) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h19) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h31) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'he) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h16) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h26) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h2a) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h32) ^ data_i[15];
    data_o[16] = (syndrome_o == 6'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 6'h2c) ^ data_i[17];
    data_o[18] = (syndrome_o == 6'h34) ^ data_i[18];
    data_o[19] = (syndrome_o == 6'h38) ^ data_i[19];
    data_o[20] = (syndrome_o == 6'h3b) ^ data_i[20];
    data_o[21] = (syndrome_o == 6'h3d) ^ data_i[21];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [38:0]
      prim_secded_39_32_enc (logic [31:0] data_i);
    logic [38:0] data_o;
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h002606BD25);
    data_o[33] = ^(data_o & 39'h00DEBA8050);
    data_o[34] = ^(data_o & 39'h00413D89AA);
    data_o[35] = ^(data_o & 39'h0031234ED1);
    data_o[36] = ^(data_o & 39'h00C2C1323B);
    data_o[37] = ^(data_o & 39'h002DCC624C);
    data_o[38] = ^(data_o & 39'h0098505586);
    return data_o;
  endfunction

  function automatic secded_39_32_t
      prim_secded_39_32_dec (logic [38:0] data_i);
    logic [31:0] data_o;
    logic [6:0] syndrome_o;
    logic [1:0]  err_o;

    secded_39_32_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 39'h012606BD25);
    syndrome_o[1] = ^(data_i & 39'h02DEBA8050);
    syndrome_o[2] = ^(data_i & 39'h04413D89AA);
    syndrome_o[3] = ^(data_i & 39'h0831234ED1);
    syndrome_o[4] = ^(data_i & 39'h10C2C1323B);
    syndrome_o[5] = ^(data_i & 39'h202DCC624C);
    syndrome_o[6] = ^(data_i & 39'h4098505586);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h19) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h54) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h61) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h34) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h1a) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h2a) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h38) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h49) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'hd) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h51) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h31) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h68) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h7) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'hb) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h25) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h26) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h46) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h70) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h32) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h2c) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h13) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h23) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h29) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h16) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h52) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [63:0]
      prim_secded_64_57_enc (logic [56:0] data_i);
    logic [63:0] data_o;
    data_o = 64'(data_i);
    data_o[57] = ^(data_o & 64'h0103FFF800007FFF);
    data_o[58] = ^(data_o & 64'h017C1FF801FF801F);
    data_o[59] = ^(data_o & 64'h01BDE1F87E0781E1);
    data_o[60] = ^(data_o & 64'h01DEEE3B8E388E22);
    data_o[61] = ^(data_o & 64'h01EF76CDB2C93244);
    data_o[62] = ^(data_o & 64'h01F7BB56D5525488);
    data_o[63] = ^(data_o & 64'h01FBDDA769A46910);
    return data_o;
  endfunction

  function automatic secded_64_57_t
      prim_secded_64_57_dec (logic [63:0] data_i);
    logic [56:0] data_o;
    logic [6:0] syndrome_o;
    logic [1:0]  err_o;

    secded_64_57_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 64'h0303FFF800007FFF);
    syndrome_o[1] = ^(data_i & 64'h057C1FF801FF801F);
    syndrome_o[2] = ^(data_i & 64'h09BDE1F87E0781E1);
    syndrome_o[3] = ^(data_i & 64'h11DEEE3B8E388E22);
    syndrome_o[4] = ^(data_i & 64'h21EF76CDB2C93244);
    syndrome_o[5] = ^(data_i & 64'h41F7BB56D5525488);
    syndrome_o[6] = ^(data_i & 64'h81FBDDA769A46910);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'hd) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h15) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h25) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h19) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h29) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h49) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h31) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h51) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h61) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'he) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h16) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h26) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h46) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h1a) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h2a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h4a) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h32) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h52) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h62) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h1c) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h2c) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h4c) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h34) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h54) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h64) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h38) ^ data_i[31];
    data_o[32] = (syndrome_o == 7'h58) ^ data_i[32];
    data_o[33] = (syndrome_o == 7'h68) ^ data_i[33];
    data_o[34] = (syndrome_o == 7'h70) ^ data_i[34];
    data_o[35] = (syndrome_o == 7'h1f) ^ data_i[35];
    data_o[36] = (syndrome_o == 7'h2f) ^ data_i[36];
    data_o[37] = (syndrome_o == 7'h4f) ^ data_i[37];
    data_o[38] = (syndrome_o == 7'h37) ^ data_i[38];
    data_o[39] = (syndrome_o == 7'h57) ^ data_i[39];
    data_o[40] = (syndrome_o == 7'h67) ^ data_i[40];
    data_o[41] = (syndrome_o == 7'h3b) ^ data_i[41];
    data_o[42] = (syndrome_o == 7'h5b) ^ data_i[42];
    data_o[43] = (syndrome_o == 7'h6b) ^ data_i[43];
    data_o[44] = (syndrome_o == 7'h73) ^ data_i[44];
    data_o[45] = (syndrome_o == 7'h3d) ^ data_i[45];
    data_o[46] = (syndrome_o == 7'h5d) ^ data_i[46];
    data_o[47] = (syndrome_o == 7'h6d) ^ data_i[47];
    data_o[48] = (syndrome_o == 7'h75) ^ data_i[48];
    data_o[49] = (syndrome_o == 7'h79) ^ data_i[49];
    data_o[50] = (syndrome_o == 7'h3e) ^ data_i[50];
    data_o[51] = (syndrome_o == 7'h5e) ^ data_i[51];
    data_o[52] = (syndrome_o == 7'h6e) ^ data_i[52];
    data_o[53] = (syndrome_o == 7'h76) ^ data_i[53];
    data_o[54] = (syndrome_o == 7'h7a) ^ data_i[54];
    data_o[55] = (syndrome_o == 7'h7c) ^ data_i[55];
    data_o[56] = (syndrome_o == 7'h7f) ^ data_i[56];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [71:0]
      prim_secded_72_64_enc (logic [63:0] data_i);
    logic [71:0] data_o;
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00B9000000001FFFFF);
    data_o[65] = ^(data_o & 72'h005E00000FFFE0003F);
    data_o[66] = ^(data_o & 72'h0067003FF003E007C1);
    data_o[67] = ^(data_o & 72'h00CD0FC0F03C207842);
    data_o[68] = ^(data_o & 72'h00B671C711C4438884);
    data_o[69] = ^(data_o & 72'h00B5B65926488C9108);
    data_o[70] = ^(data_o & 72'h00CBDAAA4A91152210);
    data_o[71] = ^(data_o & 72'h007AED348D221A4420);
    return data_o;
  endfunction

  function automatic secded_72_64_t
      prim_secded_72_64_dec (logic [71:0] data_i);
    logic [63:0] data_o;
    logic [7:0] syndrome_o;
    logic [1:0]  err_o;

    secded_72_64_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 72'h01B9000000001FFFFF);
    syndrome_o[1] = ^(data_i & 72'h025E00000FFFE0003F);
    syndrome_o[2] = ^(data_i & 72'h0467003FF003E007C1);
    syndrome_o[3] = ^(data_i & 72'h08CD0FC0F03C207842);
    syndrome_o[4] = ^(data_i & 72'h10B671C711C4438884);
    syndrome_o[5] = ^(data_i & 72'h20B5B65926488C9108);
    syndrome_o[6] = ^(data_i & 72'h40CBDAAA4A91152210);
    syndrome_o[7] = ^(data_i & 72'h807AED348D221A4420);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h83) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'hd) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h15) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h25) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h45) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h85) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h19) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h29) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h49) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h89) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h31) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h51) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h91) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h61) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'ha1) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'hc1) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h16) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h26) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h46) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h86) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'h1a) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'h2a) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'h8a) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'h32) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'h52) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'h92) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'h62) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha2) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'hc2) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'h1c) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'h2c) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'h4c) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'h8c) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'h34) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'h54) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'h94) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'h64) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'ha4) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hc4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'h38) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'h58) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'h98) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'h68) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'ha8) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hc8) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'h70) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hb0) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hd0) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'he0) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'h6d) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hd6) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'h3e) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hcb) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hb3) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hb5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hce) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'h79) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [21:0]
      prim_secded_hamming_22_16_enc (logic [15:0] data_i);
    logic [21:0] data_o;
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00AD5B);
    data_o[17] = ^(data_o & 22'h00366D);
    data_o[18] = ^(data_o & 22'h00C78E);
    data_o[19] = ^(data_o & 22'h0007F0);
    data_o[20] = ^(data_o & 22'h00F800);
    data_o[21] = ^(data_o & 22'h1FFFFF);
    return data_o;
  endfunction

  function automatic secded_hamming_22_16_t
      prim_secded_hamming_22_16_dec (logic [21:0] data_i);
    logic [15:0] data_o;
    logic [5:0] syndrome_o;
    logic [1:0]  err_o;

    secded_hamming_22_16_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 22'h01AD5B);
    syndrome_o[1] = ^(data_i & 22'h02366D);
    syndrome_o[2] = ^(data_i & 22'h04C78E);
    syndrome_o[3] = ^(data_i & 22'h0807F0);
    syndrome_o[4] = ^(data_i & 22'h10F800);
    syndrome_o[5] = ^(data_i & 22'h3FFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h23) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h25) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h26) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h27) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h29) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h2a) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h2b) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h2c) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h2d) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h2e) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h2f) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h31) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h32) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h33) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h34) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h35) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[5];
    err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [38:0]
      prim_secded_hamming_39_32_enc (logic [31:0] data_i);
    logic [38:0] data_o;
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h0056AAAD5B);
    data_o[33] = ^(data_o & 39'h009B33366D);
    data_o[34] = ^(data_o & 39'h00E3C3C78E);
    data_o[35] = ^(data_o & 39'h0003FC07F0);
    data_o[36] = ^(data_o & 39'h0003FFF800);
    data_o[37] = ^(data_o & 39'h00FC000000);
    data_o[38] = ^(data_o & 39'h3FFFFFFFFF);
    return data_o;
  endfunction

  function automatic secded_hamming_39_32_t
      prim_secded_hamming_39_32_dec (logic [38:0] data_i);
    logic [31:0] data_o;
    logic [6:0] syndrome_o;
    logic [1:0]  err_o;

    secded_hamming_39_32_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 39'h0156AAAD5B);
    syndrome_o[1] = ^(data_i & 39'h029B33366D);
    syndrome_o[2] = ^(data_i & 39'h04E3C3C78E);
    syndrome_o[3] = ^(data_i & 39'h0803FC07F0);
    syndrome_o[4] = ^(data_i & 39'h1003FFF800);
    syndrome_o[5] = ^(data_i & 39'h20FC000000);
    syndrome_o[6] = ^(data_i & 39'h7FFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h43) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h45) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h46) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h47) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h49) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h4a) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h4b) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h4d) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h4e) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h4f) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h51) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h52) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h53) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h54) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h55) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h56) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h57) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h58) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h59) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h5a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h5b) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h5c) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h5d) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h5e) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h5f) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h61) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h63) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h64) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h65) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h66) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[6];
    err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [71:0]
      prim_secded_hamming_72_64_enc (logic [63:0] data_i);
    logic [71:0] data_o;
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00AB55555556AAAD5B);
    data_o[65] = ^(data_o & 72'h00CD9999999B33366D);
    data_o[66] = ^(data_o & 72'h00F1E1E1E1E3C3C78E);
    data_o[67] = ^(data_o & 72'h0001FE01FE03FC07F0);
    data_o[68] = ^(data_o & 72'h0001FFFE0003FFF800);
    data_o[69] = ^(data_o & 72'h0001FFFFFFFC000000);
    data_o[70] = ^(data_o & 72'h00FE00000000000000);
    data_o[71] = ^(data_o & 72'h7FFFFFFFFFFFFFFFFF);
    return data_o;
  endfunction

  function automatic secded_hamming_72_64_t
      prim_secded_hamming_72_64_dec (logic [71:0] data_i);
    logic [63:0] data_o;
    logic [7:0] syndrome_o;
    logic [1:0]  err_o;

    secded_hamming_72_64_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 72'h01AB55555556AAAD5B);
    syndrome_o[1] = ^(data_i & 72'h02CD9999999B33366D);
    syndrome_o[2] = ^(data_i & 72'h04F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^(data_i & 72'h0801FE01FE03FC07F0);
    syndrome_o[4] = ^(data_i & 72'h1001FFFE0003FFF800);
    syndrome_o[5] = ^(data_i & 72'h2001FFFFFFFC000000);
    syndrome_o[6] = ^(data_i & 72'h40FE00000000000000);
    syndrome_o[7] = ^(data_i & 72'hFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [75:0]
      prim_secded_hamming_76_68_enc (logic [67:0] data_i);
    logic [75:0] data_o;
    data_o = 76'(data_i);
    data_o[68] = ^(data_o & 76'h00AAB55555556AAAD5B);
    data_o[69] = ^(data_o & 76'h00CCD9999999B33366D);
    data_o[70] = ^(data_o & 76'h000F1E1E1E1E3C3C78E);
    data_o[71] = ^(data_o & 76'h00F01FE01FE03FC07F0);
    data_o[72] = ^(data_o & 76'h00001FFFE0003FFF800);
    data_o[73] = ^(data_o & 76'h00001FFFFFFFC000000);
    data_o[74] = ^(data_o & 76'h00FFE00000000000000);
    data_o[75] = ^(data_o & 76'h7FFFFFFFFFFFFFFFFFF);
    return data_o;
  endfunction

  function automatic secded_hamming_76_68_t
      prim_secded_hamming_76_68_dec (logic [75:0] data_i);
    logic [67:0] data_o;
    logic [7:0] syndrome_o;
    logic [1:0]  err_o;

    secded_hamming_76_68_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 76'h01AAB55555556AAAD5B);
    syndrome_o[1] = ^(data_i & 76'h02CCD9999999B33366D);
    syndrome_o[2] = ^(data_i & 76'h040F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^(data_i & 76'h08F01FE01FE03FC07F0);
    syndrome_o[4] = ^(data_i & 76'h10001FFFE0003FFF800);
    syndrome_o[5] = ^(data_i & 76'h20001FFFFFFFC000000);
    syndrome_o[6] = ^(data_i & 76'h40FFE00000000000000);
    syndrome_o[7] = ^(data_i & 76'hFFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
    data_o[64] = (syndrome_o == 8'hc8) ^ data_i[64];
    data_o[65] = (syndrome_o == 8'hc9) ^ data_i[65];
    data_o[66] = (syndrome_o == 8'hca) ^ data_i[66];
    data_o[67] = (syndrome_o == 8'hcb) ^ data_i[67];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [21:0]
      prim_secded_inv_22_16_enc (logic [15:0] data_i);
    logic [21:0] data_o;
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00496E);
    data_o[17] = ^(data_o & 22'h00F20B);
    data_o[18] = ^(data_o & 22'h008ED8);
    data_o[19] = ^(data_o & 22'h007714);
    data_o[20] = ^(data_o & 22'h00ACA5);
    data_o[21] = ^(data_o & 22'h0011F3);
    data_o ^= 22'h2A0000;
    return data_o;
  endfunction

  function automatic secded_inv_22_16_t
      prim_secded_inv_22_16_dec (logic [21:0] data_i);
    logic [15:0] data_o;
    logic [5:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_22_16_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 22'h2A0000) & 22'h01496E);
    syndrome_o[1] = ^((data_i ^ 22'h2A0000) & 22'h02F20B);
    syndrome_o[2] = ^((data_i ^ 22'h2A0000) & 22'h048ED8);
    syndrome_o[3] = ^((data_i ^ 22'h2A0000) & 22'h087714);
    syndrome_o[4] = ^((data_i ^ 22'h2A0000) & 22'h10ACA5);
    syndrome_o[5] = ^((data_i ^ 22'h2A0000) & 22'h2011F3);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h32) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h23) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h19) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h7) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h2c) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h31) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h34) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'he) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h1c) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h15) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h2a) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'hb) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h16) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [27:0]
      prim_secded_inv_28_22_enc (logic [21:0] data_i);
    logic [27:0] data_o;
    data_o = 28'(data_i);
    data_o[22] = ^(data_o & 28'h03003FF);
    data_o[23] = ^(data_o & 28'h010FC0F);
    data_o[24] = ^(data_o & 28'h0271C71);
    data_o[25] = ^(data_o & 28'h03B6592);
    data_o[26] = ^(data_o & 28'h03DAAA4);
    data_o[27] = ^(data_o & 28'h03ED348);
    data_o ^= 28'hA800000;
    return data_o;
  endfunction

  function automatic secded_inv_28_22_t
      prim_secded_inv_28_22_dec (logic [27:0] data_i);
    logic [21:0] data_o;
    logic [5:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_28_22_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 28'hA800000) & 28'h07003FF);
    syndrome_o[1] = ^((data_i ^ 28'hA800000) & 28'h090FC0F);
    syndrome_o[2] = ^((data_i ^ 28'hA800000) & 28'h1271C71);
    syndrome_o[3] = ^((data_i ^ 28'hA800000) & 28'h23B6592);
    syndrome_o[4] = ^((data_i ^ 28'hA800000) & 28'h43DAAA4);
    syndrome_o[5] = ^((data_i ^ 28'hA800000) & 28'h83ED348);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'hd) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h19) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h31) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'he) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h16) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h26) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h2a) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h32) ^ data_i[15];
    data_o[16] = (syndrome_o == 6'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 6'h2c) ^ data_i[17];
    data_o[18] = (syndrome_o == 6'h34) ^ data_i[18];
    data_o[19] = (syndrome_o == 6'h38) ^ data_i[19];
    data_o[20] = (syndrome_o == 6'h3b) ^ data_i[20];
    data_o[21] = (syndrome_o == 6'h3d) ^ data_i[21];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [38:0]
      prim_secded_inv_39_32_enc (logic [31:0] data_i);
    logic [38:0] data_o;
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h002606BD25);
    data_o[33] = ^(data_o & 39'h00DEBA8050);
    data_o[34] = ^(data_o & 39'h00413D89AA);
    data_o[35] = ^(data_o & 39'h0031234ED1);
    data_o[36] = ^(data_o & 39'h00C2C1323B);
    data_o[37] = ^(data_o & 39'h002DCC624C);
    data_o[38] = ^(data_o & 39'h0098505586);
    data_o ^= 39'h2A00000000;
    return data_o;
  endfunction

  function automatic secded_inv_39_32_t
      prim_secded_inv_39_32_dec (logic [38:0] data_i);
    logic [31:0] data_o;
    logic [6:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_39_32_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 39'h2A00000000) & 39'h012606BD25);
    syndrome_o[1] = ^((data_i ^ 39'h2A00000000) & 39'h02DEBA8050);
    syndrome_o[2] = ^((data_i ^ 39'h2A00000000) & 39'h04413D89AA);
    syndrome_o[3] = ^((data_i ^ 39'h2A00000000) & 39'h0831234ED1);
    syndrome_o[4] = ^((data_i ^ 39'h2A00000000) & 39'h10C2C1323B);
    syndrome_o[5] = ^((data_i ^ 39'h2A00000000) & 39'h202DCC624C);
    syndrome_o[6] = ^((data_i ^ 39'h2A00000000) & 39'h4098505586);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h19) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h54) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h61) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h34) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h1a) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h2a) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h38) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h49) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'hd) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h51) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h31) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h68) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h7) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'hb) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h25) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h26) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h46) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h70) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h32) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h2c) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h13) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h23) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h29) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h16) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h52) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [63:0]
      prim_secded_inv_64_57_enc (logic [56:0] data_i);
    logic [63:0] data_o;
    data_o = 64'(data_i);
    data_o[57] = ^(data_o & 64'h0103FFF800007FFF);
    data_o[58] = ^(data_o & 64'h017C1FF801FF801F);
    data_o[59] = ^(data_o & 64'h01BDE1F87E0781E1);
    data_o[60] = ^(data_o & 64'h01DEEE3B8E388E22);
    data_o[61] = ^(data_o & 64'h01EF76CDB2C93244);
    data_o[62] = ^(data_o & 64'h01F7BB56D5525488);
    data_o[63] = ^(data_o & 64'h01FBDDA769A46910);
    data_o ^= 64'h5400000000000000;
    return data_o;
  endfunction

  function automatic secded_inv_64_57_t
      prim_secded_inv_64_57_dec (logic [63:0] data_i);
    logic [56:0] data_o;
    logic [6:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_64_57_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 64'h5400000000000000) & 64'h0303FFF800007FFF);
    syndrome_o[1] = ^((data_i ^ 64'h5400000000000000) & 64'h057C1FF801FF801F);
    syndrome_o[2] = ^((data_i ^ 64'h5400000000000000) & 64'h09BDE1F87E0781E1);
    syndrome_o[3] = ^((data_i ^ 64'h5400000000000000) & 64'h11DEEE3B8E388E22);
    syndrome_o[4] = ^((data_i ^ 64'h5400000000000000) & 64'h21EF76CDB2C93244);
    syndrome_o[5] = ^((data_i ^ 64'h5400000000000000) & 64'h41F7BB56D5525488);
    syndrome_o[6] = ^((data_i ^ 64'h5400000000000000) & 64'h81FBDDA769A46910);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'hd) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h15) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h25) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h19) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h29) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h49) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h31) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h51) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h61) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'he) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h16) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h26) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h46) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h1a) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h2a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h4a) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h32) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h52) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h62) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h1c) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h2c) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h4c) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h34) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h54) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h64) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h38) ^ data_i[31];
    data_o[32] = (syndrome_o == 7'h58) ^ data_i[32];
    data_o[33] = (syndrome_o == 7'h68) ^ data_i[33];
    data_o[34] = (syndrome_o == 7'h70) ^ data_i[34];
    data_o[35] = (syndrome_o == 7'h1f) ^ data_i[35];
    data_o[36] = (syndrome_o == 7'h2f) ^ data_i[36];
    data_o[37] = (syndrome_o == 7'h4f) ^ data_i[37];
    data_o[38] = (syndrome_o == 7'h37) ^ data_i[38];
    data_o[39] = (syndrome_o == 7'h57) ^ data_i[39];
    data_o[40] = (syndrome_o == 7'h67) ^ data_i[40];
    data_o[41] = (syndrome_o == 7'h3b) ^ data_i[41];
    data_o[42] = (syndrome_o == 7'h5b) ^ data_i[42];
    data_o[43] = (syndrome_o == 7'h6b) ^ data_i[43];
    data_o[44] = (syndrome_o == 7'h73) ^ data_i[44];
    data_o[45] = (syndrome_o == 7'h3d) ^ data_i[45];
    data_o[46] = (syndrome_o == 7'h5d) ^ data_i[46];
    data_o[47] = (syndrome_o == 7'h6d) ^ data_i[47];
    data_o[48] = (syndrome_o == 7'h75) ^ data_i[48];
    data_o[49] = (syndrome_o == 7'h79) ^ data_i[49];
    data_o[50] = (syndrome_o == 7'h3e) ^ data_i[50];
    data_o[51] = (syndrome_o == 7'h5e) ^ data_i[51];
    data_o[52] = (syndrome_o == 7'h6e) ^ data_i[52];
    data_o[53] = (syndrome_o == 7'h76) ^ data_i[53];
    data_o[54] = (syndrome_o == 7'h7a) ^ data_i[54];
    data_o[55] = (syndrome_o == 7'h7c) ^ data_i[55];
    data_o[56] = (syndrome_o == 7'h7f) ^ data_i[56];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [71:0]
      prim_secded_inv_72_64_enc (logic [63:0] data_i);
    logic [71:0] data_o;
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00B9000000001FFFFF);
    data_o[65] = ^(data_o & 72'h005E00000FFFE0003F);
    data_o[66] = ^(data_o & 72'h0067003FF003E007C1);
    data_o[67] = ^(data_o & 72'h00CD0FC0F03C207842);
    data_o[68] = ^(data_o & 72'h00B671C711C4438884);
    data_o[69] = ^(data_o & 72'h00B5B65926488C9108);
    data_o[70] = ^(data_o & 72'h00CBDAAA4A91152210);
    data_o[71] = ^(data_o & 72'h007AED348D221A4420);
    data_o ^= 72'hAA0000000000000000;
    return data_o;
  endfunction

  function automatic secded_inv_72_64_t
      prim_secded_inv_72_64_dec (logic [71:0] data_i);
    logic [63:0] data_o;
    logic [7:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_72_64_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 72'hAA0000000000000000) & 72'h01B9000000001FFFFF);
    syndrome_o[1] = ^((data_i ^ 72'hAA0000000000000000) & 72'h025E00000FFFE0003F);
    syndrome_o[2] = ^((data_i ^ 72'hAA0000000000000000) & 72'h0467003FF003E007C1);
    syndrome_o[3] = ^((data_i ^ 72'hAA0000000000000000) & 72'h08CD0FC0F03C207842);
    syndrome_o[4] = ^((data_i ^ 72'hAA0000000000000000) & 72'h10B671C711C4438884);
    syndrome_o[5] = ^((data_i ^ 72'hAA0000000000000000) & 72'h20B5B65926488C9108);
    syndrome_o[6] = ^((data_i ^ 72'hAA0000000000000000) & 72'h40CBDAAA4A91152210);
    syndrome_o[7] = ^((data_i ^ 72'hAA0000000000000000) & 72'h807AED348D221A4420);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h83) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'hd) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h15) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h25) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h45) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h85) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h19) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h29) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h49) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h89) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h31) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h51) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h91) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h61) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'ha1) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'hc1) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h16) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h26) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h46) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h86) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'h1a) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'h2a) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'h8a) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'h32) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'h52) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'h92) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'h62) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha2) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'hc2) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'h1c) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'h2c) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'h4c) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'h8c) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'h34) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'h54) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'h94) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'h64) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'ha4) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hc4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'h38) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'h58) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'h98) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'h68) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'ha8) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hc8) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'h70) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hb0) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hd0) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'he0) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'h6d) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hd6) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'h3e) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hcb) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hb3) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hb5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hce) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'h79) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [21:0]
      prim_secded_inv_hamming_22_16_enc (logic [15:0] data_i);
    logic [21:0] data_o;
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00AD5B);
    data_o[17] = ^(data_o & 22'h00366D);
    data_o[18] = ^(data_o & 22'h00C78E);
    data_o[19] = ^(data_o & 22'h0007F0);
    data_o[20] = ^(data_o & 22'h00F800);
    data_o[21] = ^(data_o & 22'h1FFFFF);
    data_o ^= 22'h2A0000;
    return data_o;
  endfunction

  function automatic secded_inv_hamming_22_16_t
      prim_secded_inv_hamming_22_16_dec (logic [21:0] data_i);
    logic [15:0] data_o;
    logic [5:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_hamming_22_16_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 22'h2A0000) & 22'h01AD5B);
    syndrome_o[1] = ^((data_i ^ 22'h2A0000) & 22'h02366D);
    syndrome_o[2] = ^((data_i ^ 22'h2A0000) & 22'h04C78E);
    syndrome_o[3] = ^((data_i ^ 22'h2A0000) & 22'h0807F0);
    syndrome_o[4] = ^((data_i ^ 22'h2A0000) & 22'h10F800);
    syndrome_o[5] = ^((data_i ^ 22'h2A0000) & 22'h3FFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h23) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h25) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h26) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h27) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h29) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h2a) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h2b) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h2c) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h2d) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h2e) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h2f) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h31) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h32) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h33) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h34) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h35) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[5];
    err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [38:0]
      prim_secded_inv_hamming_39_32_enc (logic [31:0] data_i);
    logic [38:0] data_o;
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h0056AAAD5B);
    data_o[33] = ^(data_o & 39'h009B33366D);
    data_o[34] = ^(data_o & 39'h00E3C3C78E);
    data_o[35] = ^(data_o & 39'h0003FC07F0);
    data_o[36] = ^(data_o & 39'h0003FFF800);
    data_o[37] = ^(data_o & 39'h00FC000000);
    data_o[38] = ^(data_o & 39'h3FFFFFFFFF);
    data_o ^= 39'h2A00000000;
    return data_o;
  endfunction

  function automatic secded_inv_hamming_39_32_t
      prim_secded_inv_hamming_39_32_dec (logic [38:0] data_i);
    logic [31:0] data_o;
    logic [6:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_hamming_39_32_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 39'h2A00000000) & 39'h0156AAAD5B);
    syndrome_o[1] = ^((data_i ^ 39'h2A00000000) & 39'h029B33366D);
    syndrome_o[2] = ^((data_i ^ 39'h2A00000000) & 39'h04E3C3C78E);
    syndrome_o[3] = ^((data_i ^ 39'h2A00000000) & 39'h0803FC07F0);
    syndrome_o[4] = ^((data_i ^ 39'h2A00000000) & 39'h1003FFF800);
    syndrome_o[5] = ^((data_i ^ 39'h2A00000000) & 39'h20FC000000);
    syndrome_o[6] = ^((data_i ^ 39'h2A00000000) & 39'h7FFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h43) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h45) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h46) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h47) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h49) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h4a) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h4b) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h4d) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h4e) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h4f) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h51) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h52) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h53) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h54) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h55) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h56) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h57) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h58) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h59) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h5a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h5b) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h5c) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h5d) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h5e) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h5f) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h61) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h63) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h64) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h65) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h66) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[6];
    err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [71:0]
      prim_secded_inv_hamming_72_64_enc (logic [63:0] data_i);
    logic [71:0] data_o;
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00AB55555556AAAD5B);
    data_o[65] = ^(data_o & 72'h00CD9999999B33366D);
    data_o[66] = ^(data_o & 72'h00F1E1E1E1E3C3C78E);
    data_o[67] = ^(data_o & 72'h0001FE01FE03FC07F0);
    data_o[68] = ^(data_o & 72'h0001FFFE0003FFF800);
    data_o[69] = ^(data_o & 72'h0001FFFFFFFC000000);
    data_o[70] = ^(data_o & 72'h00FE00000000000000);
    data_o[71] = ^(data_o & 72'h7FFFFFFFFFFFFFFFFF);
    data_o ^= 72'hAA0000000000000000;
    return data_o;
  endfunction

  function automatic secded_inv_hamming_72_64_t
      prim_secded_inv_hamming_72_64_dec (logic [71:0] data_i);
    logic [63:0] data_o;
    logic [7:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_hamming_72_64_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 72'hAA0000000000000000) & 72'h01AB55555556AAAD5B);
    syndrome_o[1] = ^((data_i ^ 72'hAA0000000000000000) & 72'h02CD9999999B33366D);
    syndrome_o[2] = ^((data_i ^ 72'hAA0000000000000000) & 72'h04F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^((data_i ^ 72'hAA0000000000000000) & 72'h0801FE01FE03FC07F0);
    syndrome_o[4] = ^((data_i ^ 72'hAA0000000000000000) & 72'h1001FFFE0003FFF800);
    syndrome_o[5] = ^((data_i ^ 72'hAA0000000000000000) & 72'h2001FFFFFFFC000000);
    syndrome_o[6] = ^((data_i ^ 72'hAA0000000000000000) & 72'h40FE00000000000000);
    syndrome_o[7] = ^((data_i ^ 72'hAA0000000000000000) & 72'hFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction

  function automatic logic [75:0]
      prim_secded_inv_hamming_76_68_enc (logic [67:0] data_i);
    logic [75:0] data_o;
    data_o = 76'(data_i);
    data_o[68] = ^(data_o & 76'h00AAB55555556AAAD5B);
    data_o[69] = ^(data_o & 76'h00CCD9999999B33366D);
    data_o[70] = ^(data_o & 76'h000F1E1E1E1E3C3C78E);
    data_o[71] = ^(data_o & 76'h00F01FE01FE03FC07F0);
    data_o[72] = ^(data_o & 76'h00001FFFE0003FFF800);
    data_o[73] = ^(data_o & 76'h00001FFFFFFFC000000);
    data_o[74] = ^(data_o & 76'h00FFE00000000000000);
    data_o[75] = ^(data_o & 76'h7FFFFFFFFFFFFFFFFFF);
    data_o ^= 76'hAA00000000000000000;
    return data_o;
  endfunction

  function automatic secded_inv_hamming_76_68_t
      prim_secded_inv_hamming_76_68_dec (logic [75:0] data_i);
    logic [67:0] data_o;
    logic [7:0] syndrome_o;
    logic [1:0]  err_o;

    secded_inv_hamming_76_68_t dec;

    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 76'hAA00000000000000000) & 76'h01AAB55555556AAAD5B);
    syndrome_o[1] = ^((data_i ^ 76'hAA00000000000000000) & 76'h02CCD9999999B33366D);
    syndrome_o[2] = ^((data_i ^ 76'hAA00000000000000000) & 76'h040F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^((data_i ^ 76'hAA00000000000000000) & 76'h08F01FE01FE03FC07F0);
    syndrome_o[4] = ^((data_i ^ 76'hAA00000000000000000) & 76'h10001FFFE0003FFF800);
    syndrome_o[5] = ^((data_i ^ 76'hAA00000000000000000) & 76'h20001FFFFFFFC000000);
    syndrome_o[6] = ^((data_i ^ 76'hAA00000000000000000) & 76'h40FFE00000000000000);
    syndrome_o[7] = ^((data_i ^ 76'hAA00000000000000000) & 76'hFFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
    data_o[64] = (syndrome_o == 8'hc8) ^ data_i[64];
    data_o[65] = (syndrome_o == 8'hc9) ^ data_i[65];
    data_o[66] = (syndrome_o == 8'hca) ^ data_i[66];
    data_o[67] = (syndrome_o == 8'hcb) ^ data_i[67];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];

    dec.data      = data_o;
    dec.syndrome  = syndrome_o;
    dec.err       = err_o;
    return dec;

  endfunction


endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_22_16_dec (
  input        [21:0] data_i,
  output logic [15:0] data_o,
  output logic [5:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 22'h01496E);
    syndrome_o[1] = ^(data_i & 22'h02F20B);
    syndrome_o[2] = ^(data_i & 22'h048ED8);
    syndrome_o[3] = ^(data_i & 22'h087714);
    syndrome_o[4] = ^(data_i & 22'h10ACA5);
    syndrome_o[5] = ^(data_i & 22'h2011F3);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h32) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h23) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h19) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h7) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h2c) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h31) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h34) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'he) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h1c) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h15) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h2a) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'hb) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h16) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_22_16_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_22_16_enc (
  input        [15:0] data_i,
  output logic [21:0] data_o
);

  always_comb begin : p_encode
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00496E);
    data_o[17] = ^(data_o & 22'h00F20B);
    data_o[18] = ^(data_o & 22'h008ED8);
    data_o[19] = ^(data_o & 22'h007714);
    data_o[20] = ^(data_o & 22'h00ACA5);
    data_o[21] = ^(data_o & 22'h0011F3);
  end

endmodule : prim_secded_22_16_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_28_22_dec (
  input        [27:0] data_i,
  output logic [21:0] data_o,
  output logic [5:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 28'h07003FF);
    syndrome_o[1] = ^(data_i & 28'h090FC0F);
    syndrome_o[2] = ^(data_i & 28'h1271C71);
    syndrome_o[3] = ^(data_i & 28'h23B6592);
    syndrome_o[4] = ^(data_i & 28'h43DAAA4);
    syndrome_o[5] = ^(data_i & 28'h83ED348);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'hd) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h19) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h31) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'he) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h16) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h26) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h2a) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h32) ^ data_i[15];
    data_o[16] = (syndrome_o == 6'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 6'h2c) ^ data_i[17];
    data_o[18] = (syndrome_o == 6'h34) ^ data_i[18];
    data_o[19] = (syndrome_o == 6'h38) ^ data_i[19];
    data_o[20] = (syndrome_o == 6'h3b) ^ data_i[20];
    data_o[21] = (syndrome_o == 6'h3d) ^ data_i[21];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_28_22_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_28_22_enc (
  input        [21:0] data_i,
  output logic [27:0] data_o
);

  always_comb begin : p_encode
    data_o = 28'(data_i);
    data_o[22] = ^(data_o & 28'h03003FF);
    data_o[23] = ^(data_o & 28'h010FC0F);
    data_o[24] = ^(data_o & 28'h0271C71);
    data_o[25] = ^(data_o & 28'h03B6592);
    data_o[26] = ^(data_o & 28'h03DAAA4);
    data_o[27] = ^(data_o & 28'h03ED348);
  end

endmodule : prim_secded_28_22_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_39_32_dec (
  input        [38:0] data_i,
  output logic [31:0] data_o,
  output logic [6:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 39'h012606BD25);
    syndrome_o[1] = ^(data_i & 39'h02DEBA8050);
    syndrome_o[2] = ^(data_i & 39'h04413D89AA);
    syndrome_o[3] = ^(data_i & 39'h0831234ED1);
    syndrome_o[4] = ^(data_i & 39'h10C2C1323B);
    syndrome_o[5] = ^(data_i & 39'h202DCC624C);
    syndrome_o[6] = ^(data_i & 39'h4098505586);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h19) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h54) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h61) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h34) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h1a) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h2a) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h38) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h49) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'hd) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h51) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h31) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h68) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h7) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'hb) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h25) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h26) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h46) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h70) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h32) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h2c) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h13) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h23) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h29) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h16) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h52) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_39_32_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_39_32_enc (
  input        [31:0] data_i,
  output logic [38:0] data_o
);

  always_comb begin : p_encode
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h002606BD25);
    data_o[33] = ^(data_o & 39'h00DEBA8050);
    data_o[34] = ^(data_o & 39'h00413D89AA);
    data_o[35] = ^(data_o & 39'h0031234ED1);
    data_o[36] = ^(data_o & 39'h00C2C1323B);
    data_o[37] = ^(data_o & 39'h002DCC624C);
    data_o[38] = ^(data_o & 39'h0098505586);
  end

endmodule : prim_secded_39_32_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_64_57_dec (
  input        [63:0] data_i,
  output logic [56:0] data_o,
  output logic [6:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 64'h0303FFF800007FFF);
    syndrome_o[1] = ^(data_i & 64'h057C1FF801FF801F);
    syndrome_o[2] = ^(data_i & 64'h09BDE1F87E0781E1);
    syndrome_o[3] = ^(data_i & 64'h11DEEE3B8E388E22);
    syndrome_o[4] = ^(data_i & 64'h21EF76CDB2C93244);
    syndrome_o[5] = ^(data_i & 64'h41F7BB56D5525488);
    syndrome_o[6] = ^(data_i & 64'h81FBDDA769A46910);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'hd) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h15) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h25) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h19) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h29) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h49) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h31) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h51) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h61) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'he) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h16) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h26) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h46) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h1a) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h2a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h4a) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h32) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h52) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h62) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h1c) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h2c) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h4c) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h34) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h54) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h64) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h38) ^ data_i[31];
    data_o[32] = (syndrome_o == 7'h58) ^ data_i[32];
    data_o[33] = (syndrome_o == 7'h68) ^ data_i[33];
    data_o[34] = (syndrome_o == 7'h70) ^ data_i[34];
    data_o[35] = (syndrome_o == 7'h1f) ^ data_i[35];
    data_o[36] = (syndrome_o == 7'h2f) ^ data_i[36];
    data_o[37] = (syndrome_o == 7'h4f) ^ data_i[37];
    data_o[38] = (syndrome_o == 7'h37) ^ data_i[38];
    data_o[39] = (syndrome_o == 7'h57) ^ data_i[39];
    data_o[40] = (syndrome_o == 7'h67) ^ data_i[40];
    data_o[41] = (syndrome_o == 7'h3b) ^ data_i[41];
    data_o[42] = (syndrome_o == 7'h5b) ^ data_i[42];
    data_o[43] = (syndrome_o == 7'h6b) ^ data_i[43];
    data_o[44] = (syndrome_o == 7'h73) ^ data_i[44];
    data_o[45] = (syndrome_o == 7'h3d) ^ data_i[45];
    data_o[46] = (syndrome_o == 7'h5d) ^ data_i[46];
    data_o[47] = (syndrome_o == 7'h6d) ^ data_i[47];
    data_o[48] = (syndrome_o == 7'h75) ^ data_i[48];
    data_o[49] = (syndrome_o == 7'h79) ^ data_i[49];
    data_o[50] = (syndrome_o == 7'h3e) ^ data_i[50];
    data_o[51] = (syndrome_o == 7'h5e) ^ data_i[51];
    data_o[52] = (syndrome_o == 7'h6e) ^ data_i[52];
    data_o[53] = (syndrome_o == 7'h76) ^ data_i[53];
    data_o[54] = (syndrome_o == 7'h7a) ^ data_i[54];
    data_o[55] = (syndrome_o == 7'h7c) ^ data_i[55];
    data_o[56] = (syndrome_o == 7'h7f) ^ data_i[56];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_64_57_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_64_57_enc (
  input        [56:0] data_i,
  output logic [63:0] data_o
);

  always_comb begin : p_encode
    data_o = 64'(data_i);
    data_o[57] = ^(data_o & 64'h0103FFF800007FFF);
    data_o[58] = ^(data_o & 64'h017C1FF801FF801F);
    data_o[59] = ^(data_o & 64'h01BDE1F87E0781E1);
    data_o[60] = ^(data_o & 64'h01DEEE3B8E388E22);
    data_o[61] = ^(data_o & 64'h01EF76CDB2C93244);
    data_o[62] = ^(data_o & 64'h01F7BB56D5525488);
    data_o[63] = ^(data_o & 64'h01FBDDA769A46910);
  end

endmodule : prim_secded_64_57_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_72_64_dec (
  input        [71:0] data_i,
  output logic [63:0] data_o,
  output logic [7:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 72'h01B9000000001FFFFF);
    syndrome_o[1] = ^(data_i & 72'h025E00000FFFE0003F);
    syndrome_o[2] = ^(data_i & 72'h0467003FF003E007C1);
    syndrome_o[3] = ^(data_i & 72'h08CD0FC0F03C207842);
    syndrome_o[4] = ^(data_i & 72'h10B671C711C4438884);
    syndrome_o[5] = ^(data_i & 72'h20B5B65926488C9108);
    syndrome_o[6] = ^(data_i & 72'h40CBDAAA4A91152210);
    syndrome_o[7] = ^(data_i & 72'h807AED348D221A4420);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h83) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'hd) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h15) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h25) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h45) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h85) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h19) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h29) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h49) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h89) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h31) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h51) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h91) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h61) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'ha1) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'hc1) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h16) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h26) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h46) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h86) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'h1a) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'h2a) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'h8a) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'h32) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'h52) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'h92) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'h62) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha2) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'hc2) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'h1c) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'h2c) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'h4c) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'h8c) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'h34) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'h54) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'h94) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'h64) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'ha4) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hc4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'h38) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'h58) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'h98) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'h68) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'ha8) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hc8) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'h70) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hb0) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hd0) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'he0) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'h6d) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hd6) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'h3e) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hcb) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hb3) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hb5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hce) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'h79) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_72_64_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_72_64_enc (
  input        [63:0] data_i,
  output logic [71:0] data_o
);

  always_comb begin : p_encode
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00B9000000001FFFFF);
    data_o[65] = ^(data_o & 72'h005E00000FFFE0003F);
    data_o[66] = ^(data_o & 72'h0067003FF003E007C1);
    data_o[67] = ^(data_o & 72'h00CD0FC0F03C207842);
    data_o[68] = ^(data_o & 72'h00B671C711C4438884);
    data_o[69] = ^(data_o & 72'h00B5B65926488C9108);
    data_o[70] = ^(data_o & 72'h00CBDAAA4A91152210);
    data_o[71] = ^(data_o & 72'h007AED348D221A4420);
  end

endmodule : prim_secded_72_64_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_hamming_22_16_dec (
  input        [21:0] data_i,
  output logic [15:0] data_o,
  output logic [5:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 22'h01AD5B);
    syndrome_o[1] = ^(data_i & 22'h02366D);
    syndrome_o[2] = ^(data_i & 22'h04C78E);
    syndrome_o[3] = ^(data_i & 22'h0807F0);
    syndrome_o[4] = ^(data_i & 22'h10F800);
    syndrome_o[5] = ^(data_i & 22'h3FFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h23) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h25) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h26) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h27) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h29) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h2a) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h2b) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h2c) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h2d) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h2e) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h2f) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h31) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h32) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h33) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h34) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h35) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[5];
    err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];
  end
endmodule : prim_secded_hamming_22_16_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_hamming_22_16_enc (
  input        [15:0] data_i,
  output logic [21:0] data_o
);

  always_comb begin : p_encode
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00AD5B);
    data_o[17] = ^(data_o & 22'h00366D);
    data_o[18] = ^(data_o & 22'h00C78E);
    data_o[19] = ^(data_o & 22'h0007F0);
    data_o[20] = ^(data_o & 22'h00F800);
    data_o[21] = ^(data_o & 22'h1FFFFF);
  end

endmodule : prim_secded_hamming_22_16_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_hamming_39_32_dec (
  input        [38:0] data_i,
  output logic [31:0] data_o,
  output logic [6:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 39'h0156AAAD5B);
    syndrome_o[1] = ^(data_i & 39'h029B33366D);
    syndrome_o[2] = ^(data_i & 39'h04E3C3C78E);
    syndrome_o[3] = ^(data_i & 39'h0803FC07F0);
    syndrome_o[4] = ^(data_i & 39'h1003FFF800);
    syndrome_o[5] = ^(data_i & 39'h20FC000000);
    syndrome_o[6] = ^(data_i & 39'h7FFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h43) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h45) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h46) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h47) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h49) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h4a) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h4b) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h4d) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h4e) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h4f) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h51) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h52) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h53) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h54) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h55) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h56) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h57) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h58) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h59) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h5a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h5b) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h5c) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h5d) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h5e) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h5f) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h61) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h63) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h64) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h65) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h66) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[6];
    err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];
  end
endmodule : prim_secded_hamming_39_32_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_hamming_39_32_enc (
  input        [31:0] data_i,
  output logic [38:0] data_o
);

  always_comb begin : p_encode
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h0056AAAD5B);
    data_o[33] = ^(data_o & 39'h009B33366D);
    data_o[34] = ^(data_o & 39'h00E3C3C78E);
    data_o[35] = ^(data_o & 39'h0003FC07F0);
    data_o[36] = ^(data_o & 39'h0003FFF800);
    data_o[37] = ^(data_o & 39'h00FC000000);
    data_o[38] = ^(data_o & 39'h3FFFFFFFFF);
  end

endmodule : prim_secded_hamming_39_32_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_hamming_72_64_dec (
  input        [71:0] data_i,
  output logic [63:0] data_o,
  output logic [7:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 72'h01AB55555556AAAD5B);
    syndrome_o[1] = ^(data_i & 72'h02CD9999999B33366D);
    syndrome_o[2] = ^(data_i & 72'h04F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^(data_i & 72'h0801FE01FE03FC07F0);
    syndrome_o[4] = ^(data_i & 72'h1001FFFE0003FFF800);
    syndrome_o[5] = ^(data_i & 72'h2001FFFFFFFC000000);
    syndrome_o[6] = ^(data_i & 72'h40FE00000000000000);
    syndrome_o[7] = ^(data_i & 72'hFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
  end
endmodule : prim_secded_hamming_72_64_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_hamming_72_64_enc (
  input        [63:0] data_i,
  output logic [71:0] data_o
);

  always_comb begin : p_encode
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00AB55555556AAAD5B);
    data_o[65] = ^(data_o & 72'h00CD9999999B33366D);
    data_o[66] = ^(data_o & 72'h00F1E1E1E1E3C3C78E);
    data_o[67] = ^(data_o & 72'h0001FE01FE03FC07F0);
    data_o[68] = ^(data_o & 72'h0001FFFE0003FFF800);
    data_o[69] = ^(data_o & 72'h0001FFFFFFFC000000);
    data_o[70] = ^(data_o & 72'h00FE00000000000000);
    data_o[71] = ^(data_o & 72'h7FFFFFFFFFFFFFFFFF);
  end

endmodule : prim_secded_hamming_72_64_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_hamming_76_68_dec (
  input        [75:0] data_i,
  output logic [67:0] data_o,
  output logic [7:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^(data_i & 76'h01AAB55555556AAAD5B);
    syndrome_o[1] = ^(data_i & 76'h02CCD9999999B33366D);
    syndrome_o[2] = ^(data_i & 76'h040F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^(data_i & 76'h08F01FE01FE03FC07F0);
    syndrome_o[4] = ^(data_i & 76'h10001FFFE0003FFF800);
    syndrome_o[5] = ^(data_i & 76'h20001FFFFFFFC000000);
    syndrome_o[6] = ^(data_i & 76'h40FFE00000000000000);
    syndrome_o[7] = ^(data_i & 76'hFFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
    data_o[64] = (syndrome_o == 8'hc8) ^ data_i[64];
    data_o[65] = (syndrome_o == 8'hc9) ^ data_i[65];
    data_o[66] = (syndrome_o == 8'hca) ^ data_i[66];
    data_o[67] = (syndrome_o == 8'hcb) ^ data_i[67];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
  end
endmodule : prim_secded_hamming_76_68_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_hamming_76_68_enc (
  input        [67:0] data_i,
  output logic [75:0] data_o
);

  always_comb begin : p_encode
    data_o = 76'(data_i);
    data_o[68] = ^(data_o & 76'h00AAB55555556AAAD5B);
    data_o[69] = ^(data_o & 76'h00CCD9999999B33366D);
    data_o[70] = ^(data_o & 76'h000F1E1E1E1E3C3C78E);
    data_o[71] = ^(data_o & 76'h00F01FE01FE03FC07F0);
    data_o[72] = ^(data_o & 76'h00001FFFE0003FFF800);
    data_o[73] = ^(data_o & 76'h00001FFFFFFFC000000);
    data_o[74] = ^(data_o & 76'h00FFE00000000000000);
    data_o[75] = ^(data_o & 76'h7FFFFFFFFFFFFFFFFFF);
  end

endmodule : prim_secded_hamming_76_68_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_22_16_dec (
  input        [21:0] data_i,
  output logic [15:0] data_o,
  output logic [5:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 22'h2A0000) & 22'h01496E);
    syndrome_o[1] = ^((data_i ^ 22'h2A0000) & 22'h02F20B);
    syndrome_o[2] = ^((data_i ^ 22'h2A0000) & 22'h048ED8);
    syndrome_o[3] = ^((data_i ^ 22'h2A0000) & 22'h087714);
    syndrome_o[4] = ^((data_i ^ 22'h2A0000) & 22'h10ACA5);
    syndrome_o[5] = ^((data_i ^ 22'h2A0000) & 22'h2011F3);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h32) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h23) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h19) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h7) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h2c) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h31) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h34) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'he) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h1c) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h15) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h2a) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'hb) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h16) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_inv_22_16_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_22_16_enc (
  input        [15:0] data_i,
  output logic [21:0] data_o
);

  always_comb begin : p_encode
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00496E);
    data_o[17] = ^(data_o & 22'h00F20B);
    data_o[18] = ^(data_o & 22'h008ED8);
    data_o[19] = ^(data_o & 22'h007714);
    data_o[20] = ^(data_o & 22'h00ACA5);
    data_o[21] = ^(data_o & 22'h0011F3);
    data_o ^= 22'h2A0000;
  end

endmodule : prim_secded_inv_22_16_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_28_22_dec (
  input        [27:0] data_i,
  output logic [21:0] data_o,
  output logic [5:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 28'hA800000) & 28'h07003FF);
    syndrome_o[1] = ^((data_i ^ 28'hA800000) & 28'h090FC0F);
    syndrome_o[2] = ^((data_i ^ 28'hA800000) & 28'h1271C71);
    syndrome_o[3] = ^((data_i ^ 28'hA800000) & 28'h23B6592);
    syndrome_o[4] = ^((data_i ^ 28'hA800000) & 28'h43DAAA4);
    syndrome_o[5] = ^((data_i ^ 28'hA800000) & 28'h83ED348);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'hd) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h25) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h19) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h29) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h31) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'he) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h16) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h26) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h1a) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h2a) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h32) ^ data_i[15];
    data_o[16] = (syndrome_o == 6'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 6'h2c) ^ data_i[17];
    data_o[18] = (syndrome_o == 6'h34) ^ data_i[18];
    data_o[19] = (syndrome_o == 6'h38) ^ data_i[19];
    data_o[20] = (syndrome_o == 6'h3b) ^ data_i[20];
    data_o[21] = (syndrome_o == 6'h3d) ^ data_i[21];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_inv_28_22_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_28_22_enc (
  input        [21:0] data_i,
  output logic [27:0] data_o
);

  always_comb begin : p_encode
    data_o = 28'(data_i);
    data_o[22] = ^(data_o & 28'h03003FF);
    data_o[23] = ^(data_o & 28'h010FC0F);
    data_o[24] = ^(data_o & 28'h0271C71);
    data_o[25] = ^(data_o & 28'h03B6592);
    data_o[26] = ^(data_o & 28'h03DAAA4);
    data_o[27] = ^(data_o & 28'h03ED348);
    data_o ^= 28'hA800000;
  end

endmodule : prim_secded_inv_28_22_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_39_32_dec (
  input        [38:0] data_i,
  output logic [31:0] data_o,
  output logic [6:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 39'h2A00000000) & 39'h012606BD25);
    syndrome_o[1] = ^((data_i ^ 39'h2A00000000) & 39'h02DEBA8050);
    syndrome_o[2] = ^((data_i ^ 39'h2A00000000) & 39'h04413D89AA);
    syndrome_o[3] = ^((data_i ^ 39'h2A00000000) & 39'h0831234ED1);
    syndrome_o[4] = ^((data_i ^ 39'h2A00000000) & 39'h10C2C1323B);
    syndrome_o[5] = ^((data_i ^ 39'h2A00000000) & 39'h202DCC624C);
    syndrome_o[6] = ^((data_i ^ 39'h2A00000000) & 39'h4098505586);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h19) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h54) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h61) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h34) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h1a) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h15) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h2a) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h38) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h49) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'hd) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h51) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h31) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h68) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h7) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h1c) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'hb) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h25) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h26) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h46) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h70) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h32) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h2c) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h13) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h23) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h29) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h16) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h52) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_inv_39_32_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_39_32_enc (
  input        [31:0] data_i,
  output logic [38:0] data_o
);

  always_comb begin : p_encode
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h002606BD25);
    data_o[33] = ^(data_o & 39'h00DEBA8050);
    data_o[34] = ^(data_o & 39'h00413D89AA);
    data_o[35] = ^(data_o & 39'h0031234ED1);
    data_o[36] = ^(data_o & 39'h00C2C1323B);
    data_o[37] = ^(data_o & 39'h002DCC624C);
    data_o[38] = ^(data_o & 39'h0098505586);
    data_o ^= 39'h2A00000000;
  end

endmodule : prim_secded_inv_39_32_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_64_57_dec (
  input        [63:0] data_i,
  output logic [56:0] data_o,
  output logic [6:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 64'h5400000000000000) & 64'h0303FFF800007FFF);
    syndrome_o[1] = ^((data_i ^ 64'h5400000000000000) & 64'h057C1FF801FF801F);
    syndrome_o[2] = ^((data_i ^ 64'h5400000000000000) & 64'h09BDE1F87E0781E1);
    syndrome_o[3] = ^((data_i ^ 64'h5400000000000000) & 64'h11DEEE3B8E388E22);
    syndrome_o[4] = ^((data_i ^ 64'h5400000000000000) & 64'h21EF76CDB2C93244);
    syndrome_o[5] = ^((data_i ^ 64'h5400000000000000) & 64'h41F7BB56D5525488);
    syndrome_o[6] = ^((data_i ^ 64'h5400000000000000) & 64'h81FBDDA769A46910);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'hd) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h15) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h25) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h45) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h19) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h29) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h49) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h31) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h51) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h61) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'he) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h16) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h26) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h46) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h1a) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h2a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h4a) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h32) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h52) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h62) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h1c) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h2c) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h4c) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h34) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h54) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h64) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h38) ^ data_i[31];
    data_o[32] = (syndrome_o == 7'h58) ^ data_i[32];
    data_o[33] = (syndrome_o == 7'h68) ^ data_i[33];
    data_o[34] = (syndrome_o == 7'h70) ^ data_i[34];
    data_o[35] = (syndrome_o == 7'h1f) ^ data_i[35];
    data_o[36] = (syndrome_o == 7'h2f) ^ data_i[36];
    data_o[37] = (syndrome_o == 7'h4f) ^ data_i[37];
    data_o[38] = (syndrome_o == 7'h37) ^ data_i[38];
    data_o[39] = (syndrome_o == 7'h57) ^ data_i[39];
    data_o[40] = (syndrome_o == 7'h67) ^ data_i[40];
    data_o[41] = (syndrome_o == 7'h3b) ^ data_i[41];
    data_o[42] = (syndrome_o == 7'h5b) ^ data_i[42];
    data_o[43] = (syndrome_o == 7'h6b) ^ data_i[43];
    data_o[44] = (syndrome_o == 7'h73) ^ data_i[44];
    data_o[45] = (syndrome_o == 7'h3d) ^ data_i[45];
    data_o[46] = (syndrome_o == 7'h5d) ^ data_i[46];
    data_o[47] = (syndrome_o == 7'h6d) ^ data_i[47];
    data_o[48] = (syndrome_o == 7'h75) ^ data_i[48];
    data_o[49] = (syndrome_o == 7'h79) ^ data_i[49];
    data_o[50] = (syndrome_o == 7'h3e) ^ data_i[50];
    data_o[51] = (syndrome_o == 7'h5e) ^ data_i[51];
    data_o[52] = (syndrome_o == 7'h6e) ^ data_i[52];
    data_o[53] = (syndrome_o == 7'h76) ^ data_i[53];
    data_o[54] = (syndrome_o == 7'h7a) ^ data_i[54];
    data_o[55] = (syndrome_o == 7'h7c) ^ data_i[55];
    data_o[56] = (syndrome_o == 7'h7f) ^ data_i[56];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_inv_64_57_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_64_57_enc (
  input        [56:0] data_i,
  output logic [63:0] data_o
);

  always_comb begin : p_encode
    data_o = 64'(data_i);
    data_o[57] = ^(data_o & 64'h0103FFF800007FFF);
    data_o[58] = ^(data_o & 64'h017C1FF801FF801F);
    data_o[59] = ^(data_o & 64'h01BDE1F87E0781E1);
    data_o[60] = ^(data_o & 64'h01DEEE3B8E388E22);
    data_o[61] = ^(data_o & 64'h01EF76CDB2C93244);
    data_o[62] = ^(data_o & 64'h01F7BB56D5525488);
    data_o[63] = ^(data_o & 64'h01FBDDA769A46910);
    data_o ^= 64'h5400000000000000;
  end

endmodule : prim_secded_inv_64_57_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_72_64_dec (
  input        [71:0] data_i,
  output logic [63:0] data_o,
  output logic [7:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 72'hAA0000000000000000) & 72'h01B9000000001FFFFF);
    syndrome_o[1] = ^((data_i ^ 72'hAA0000000000000000) & 72'h025E00000FFFE0003F);
    syndrome_o[2] = ^((data_i ^ 72'hAA0000000000000000) & 72'h0467003FF003E007C1);
    syndrome_o[3] = ^((data_i ^ 72'hAA0000000000000000) & 72'h08CD0FC0F03C207842);
    syndrome_o[4] = ^((data_i ^ 72'hAA0000000000000000) & 72'h10B671C711C4438884);
    syndrome_o[5] = ^((data_i ^ 72'hAA0000000000000000) & 72'h20B5B65926488C9108);
    syndrome_o[6] = ^((data_i ^ 72'hAA0000000000000000) & 72'h40CBDAAA4A91152210);
    syndrome_o[7] = ^((data_i ^ 72'hAA0000000000000000) & 72'h807AED348D221A4420);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h7) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'hb) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h13) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h23) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h43) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h83) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'hd) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h15) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h25) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h45) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h85) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h19) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h29) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h49) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h89) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h31) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h51) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h91) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h61) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'ha1) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'hc1) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'he) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h16) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h26) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h46) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h86) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'h1a) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'h2a) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'h4a) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'h8a) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'h32) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'h52) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'h92) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'h62) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha2) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'hc2) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'h1c) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'h2c) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'h4c) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'h8c) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'h34) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'h54) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'h94) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'h64) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'ha4) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hc4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'h38) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'h58) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'h98) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'h68) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'ha8) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hc8) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'h70) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hb0) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hd0) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'he0) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'h6d) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hd6) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'h3e) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hcb) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hb3) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hb5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hce) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'h79) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = ^syndrome_o;
    err_o[1] = ~err_o[0] & (|syndrome_o);
  end
endmodule : prim_secded_inv_72_64_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_72_64_enc (
  input        [63:0] data_i,
  output logic [71:0] data_o
);

  always_comb begin : p_encode
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00B9000000001FFFFF);
    data_o[65] = ^(data_o & 72'h005E00000FFFE0003F);
    data_o[66] = ^(data_o & 72'h0067003FF003E007C1);
    data_o[67] = ^(data_o & 72'h00CD0FC0F03C207842);
    data_o[68] = ^(data_o & 72'h00B671C711C4438884);
    data_o[69] = ^(data_o & 72'h00B5B65926488C9108);
    data_o[70] = ^(data_o & 72'h00CBDAAA4A91152210);
    data_o[71] = ^(data_o & 72'h007AED348D221A4420);
    data_o ^= 72'hAA0000000000000000;
  end

endmodule : prim_secded_inv_72_64_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_22_16_dec (
  input        [21:0] data_i,
  output logic [15:0] data_o,
  output logic [5:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 22'h2A0000) & 22'h01AD5B);
    syndrome_o[1] = ^((data_i ^ 22'h2A0000) & 22'h02366D);
    syndrome_o[2] = ^((data_i ^ 22'h2A0000) & 22'h04C78E);
    syndrome_o[3] = ^((data_i ^ 22'h2A0000) & 22'h0807F0);
    syndrome_o[4] = ^((data_i ^ 22'h2A0000) & 22'h10F800);
    syndrome_o[5] = ^((data_i ^ 22'h2A0000) & 22'h3FFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 6'h23) ^ data_i[0];
    data_o[1] = (syndrome_o == 6'h25) ^ data_i[1];
    data_o[2] = (syndrome_o == 6'h26) ^ data_i[2];
    data_o[3] = (syndrome_o == 6'h27) ^ data_i[3];
    data_o[4] = (syndrome_o == 6'h29) ^ data_i[4];
    data_o[5] = (syndrome_o == 6'h2a) ^ data_i[5];
    data_o[6] = (syndrome_o == 6'h2b) ^ data_i[6];
    data_o[7] = (syndrome_o == 6'h2c) ^ data_i[7];
    data_o[8] = (syndrome_o == 6'h2d) ^ data_i[8];
    data_o[9] = (syndrome_o == 6'h2e) ^ data_i[9];
    data_o[10] = (syndrome_o == 6'h2f) ^ data_i[10];
    data_o[11] = (syndrome_o == 6'h31) ^ data_i[11];
    data_o[12] = (syndrome_o == 6'h32) ^ data_i[12];
    data_o[13] = (syndrome_o == 6'h33) ^ data_i[13];
    data_o[14] = (syndrome_o == 6'h34) ^ data_i[14];
    data_o[15] = (syndrome_o == 6'h35) ^ data_i[15];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[5];
    err_o[1] = |syndrome_o[4:0] & ~syndrome_o[5];
  end
endmodule : prim_secded_inv_hamming_22_16_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_22_16_enc (
  input        [15:0] data_i,
  output logic [21:0] data_o
);

  always_comb begin : p_encode
    data_o = 22'(data_i);
    data_o[16] = ^(data_o & 22'h00AD5B);
    data_o[17] = ^(data_o & 22'h00366D);
    data_o[18] = ^(data_o & 22'h00C78E);
    data_o[19] = ^(data_o & 22'h0007F0);
    data_o[20] = ^(data_o & 22'h00F800);
    data_o[21] = ^(data_o & 22'h1FFFFF);
    data_o ^= 22'h2A0000;
  end

endmodule : prim_secded_inv_hamming_22_16_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_39_32_dec (
  input        [38:0] data_i,
  output logic [31:0] data_o,
  output logic [6:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 39'h2A00000000) & 39'h0156AAAD5B);
    syndrome_o[1] = ^((data_i ^ 39'h2A00000000) & 39'h029B33366D);
    syndrome_o[2] = ^((data_i ^ 39'h2A00000000) & 39'h04E3C3C78E);
    syndrome_o[3] = ^((data_i ^ 39'h2A00000000) & 39'h0803FC07F0);
    syndrome_o[4] = ^((data_i ^ 39'h2A00000000) & 39'h1003FFF800);
    syndrome_o[5] = ^((data_i ^ 39'h2A00000000) & 39'h20FC000000);
    syndrome_o[6] = ^((data_i ^ 39'h2A00000000) & 39'h7FFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 7'h43) ^ data_i[0];
    data_o[1] = (syndrome_o == 7'h45) ^ data_i[1];
    data_o[2] = (syndrome_o == 7'h46) ^ data_i[2];
    data_o[3] = (syndrome_o == 7'h47) ^ data_i[3];
    data_o[4] = (syndrome_o == 7'h49) ^ data_i[4];
    data_o[5] = (syndrome_o == 7'h4a) ^ data_i[5];
    data_o[6] = (syndrome_o == 7'h4b) ^ data_i[6];
    data_o[7] = (syndrome_o == 7'h4c) ^ data_i[7];
    data_o[8] = (syndrome_o == 7'h4d) ^ data_i[8];
    data_o[9] = (syndrome_o == 7'h4e) ^ data_i[9];
    data_o[10] = (syndrome_o == 7'h4f) ^ data_i[10];
    data_o[11] = (syndrome_o == 7'h51) ^ data_i[11];
    data_o[12] = (syndrome_o == 7'h52) ^ data_i[12];
    data_o[13] = (syndrome_o == 7'h53) ^ data_i[13];
    data_o[14] = (syndrome_o == 7'h54) ^ data_i[14];
    data_o[15] = (syndrome_o == 7'h55) ^ data_i[15];
    data_o[16] = (syndrome_o == 7'h56) ^ data_i[16];
    data_o[17] = (syndrome_o == 7'h57) ^ data_i[17];
    data_o[18] = (syndrome_o == 7'h58) ^ data_i[18];
    data_o[19] = (syndrome_o == 7'h59) ^ data_i[19];
    data_o[20] = (syndrome_o == 7'h5a) ^ data_i[20];
    data_o[21] = (syndrome_o == 7'h5b) ^ data_i[21];
    data_o[22] = (syndrome_o == 7'h5c) ^ data_i[22];
    data_o[23] = (syndrome_o == 7'h5d) ^ data_i[23];
    data_o[24] = (syndrome_o == 7'h5e) ^ data_i[24];
    data_o[25] = (syndrome_o == 7'h5f) ^ data_i[25];
    data_o[26] = (syndrome_o == 7'h61) ^ data_i[26];
    data_o[27] = (syndrome_o == 7'h62) ^ data_i[27];
    data_o[28] = (syndrome_o == 7'h63) ^ data_i[28];
    data_o[29] = (syndrome_o == 7'h64) ^ data_i[29];
    data_o[30] = (syndrome_o == 7'h65) ^ data_i[30];
    data_o[31] = (syndrome_o == 7'h66) ^ data_i[31];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[6];
    err_o[1] = |syndrome_o[5:0] & ~syndrome_o[6];
  end
endmodule : prim_secded_inv_hamming_39_32_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_39_32_enc (
  input        [31:0] data_i,
  output logic [38:0] data_o
);

  always_comb begin : p_encode
    data_o = 39'(data_i);
    data_o[32] = ^(data_o & 39'h0056AAAD5B);
    data_o[33] = ^(data_o & 39'h009B33366D);
    data_o[34] = ^(data_o & 39'h00E3C3C78E);
    data_o[35] = ^(data_o & 39'h0003FC07F0);
    data_o[36] = ^(data_o & 39'h0003FFF800);
    data_o[37] = ^(data_o & 39'h00FC000000);
    data_o[38] = ^(data_o & 39'h3FFFFFFFFF);
    data_o ^= 39'h2A00000000;
  end

endmodule : prim_secded_inv_hamming_39_32_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_72_64_dec (
  input        [71:0] data_i,
  output logic [63:0] data_o,
  output logic [7:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 72'hAA0000000000000000) & 72'h01AB55555556AAAD5B);
    syndrome_o[1] = ^((data_i ^ 72'hAA0000000000000000) & 72'h02CD9999999B33366D);
    syndrome_o[2] = ^((data_i ^ 72'hAA0000000000000000) & 72'h04F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^((data_i ^ 72'hAA0000000000000000) & 72'h0801FE01FE03FC07F0);
    syndrome_o[4] = ^((data_i ^ 72'hAA0000000000000000) & 72'h1001FFFE0003FFF800);
    syndrome_o[5] = ^((data_i ^ 72'hAA0000000000000000) & 72'h2001FFFFFFFC000000);
    syndrome_o[6] = ^((data_i ^ 72'hAA0000000000000000) & 72'h40FE00000000000000);
    syndrome_o[7] = ^((data_i ^ 72'hAA0000000000000000) & 72'hFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
  end
endmodule : prim_secded_inv_hamming_72_64_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_72_64_enc (
  input        [63:0] data_i,
  output logic [71:0] data_o
);

  always_comb begin : p_encode
    data_o = 72'(data_i);
    data_o[64] = ^(data_o & 72'h00AB55555556AAAD5B);
    data_o[65] = ^(data_o & 72'h00CD9999999B33366D);
    data_o[66] = ^(data_o & 72'h00F1E1E1E1E3C3C78E);
    data_o[67] = ^(data_o & 72'h0001FE01FE03FC07F0);
    data_o[68] = ^(data_o & 72'h0001FFFE0003FFF800);
    data_o[69] = ^(data_o & 72'h0001FFFFFFFC000000);
    data_o[70] = ^(data_o & 72'h00FE00000000000000);
    data_o[71] = ^(data_o & 72'h7FFFFFFFFFFFFFFFFF);
    data_o ^= 72'hAA0000000000000000;
  end

endmodule : prim_secded_inv_hamming_72_64_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED decoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_76_68_dec (
  input        [75:0] data_i,
  output logic [67:0] data_o,
  output logic [7:0] syndrome_o,
  output logic [1:0] err_o
);

  always_comb begin : p_encode
    // Syndrome calculation
    syndrome_o[0] = ^((data_i ^ 76'hAA00000000000000000) & 76'h01AAB55555556AAAD5B);
    syndrome_o[1] = ^((data_i ^ 76'hAA00000000000000000) & 76'h02CCD9999999B33366D);
    syndrome_o[2] = ^((data_i ^ 76'hAA00000000000000000) & 76'h040F1E1E1E1E3C3C78E);
    syndrome_o[3] = ^((data_i ^ 76'hAA00000000000000000) & 76'h08F01FE01FE03FC07F0);
    syndrome_o[4] = ^((data_i ^ 76'hAA00000000000000000) & 76'h10001FFFE0003FFF800);
    syndrome_o[5] = ^((data_i ^ 76'hAA00000000000000000) & 76'h20001FFFFFFFC000000);
    syndrome_o[6] = ^((data_i ^ 76'hAA00000000000000000) & 76'h40FFE00000000000000);
    syndrome_o[7] = ^((data_i ^ 76'hAA00000000000000000) & 76'hFFFFFFFFFFFFFFFFFFF);

    // Corrected output calculation
    data_o[0] = (syndrome_o == 8'h83) ^ data_i[0];
    data_o[1] = (syndrome_o == 8'h85) ^ data_i[1];
    data_o[2] = (syndrome_o == 8'h86) ^ data_i[2];
    data_o[3] = (syndrome_o == 8'h87) ^ data_i[3];
    data_o[4] = (syndrome_o == 8'h89) ^ data_i[4];
    data_o[5] = (syndrome_o == 8'h8a) ^ data_i[5];
    data_o[6] = (syndrome_o == 8'h8b) ^ data_i[6];
    data_o[7] = (syndrome_o == 8'h8c) ^ data_i[7];
    data_o[8] = (syndrome_o == 8'h8d) ^ data_i[8];
    data_o[9] = (syndrome_o == 8'h8e) ^ data_i[9];
    data_o[10] = (syndrome_o == 8'h8f) ^ data_i[10];
    data_o[11] = (syndrome_o == 8'h91) ^ data_i[11];
    data_o[12] = (syndrome_o == 8'h92) ^ data_i[12];
    data_o[13] = (syndrome_o == 8'h93) ^ data_i[13];
    data_o[14] = (syndrome_o == 8'h94) ^ data_i[14];
    data_o[15] = (syndrome_o == 8'h95) ^ data_i[15];
    data_o[16] = (syndrome_o == 8'h96) ^ data_i[16];
    data_o[17] = (syndrome_o == 8'h97) ^ data_i[17];
    data_o[18] = (syndrome_o == 8'h98) ^ data_i[18];
    data_o[19] = (syndrome_o == 8'h99) ^ data_i[19];
    data_o[20] = (syndrome_o == 8'h9a) ^ data_i[20];
    data_o[21] = (syndrome_o == 8'h9b) ^ data_i[21];
    data_o[22] = (syndrome_o == 8'h9c) ^ data_i[22];
    data_o[23] = (syndrome_o == 8'h9d) ^ data_i[23];
    data_o[24] = (syndrome_o == 8'h9e) ^ data_i[24];
    data_o[25] = (syndrome_o == 8'h9f) ^ data_i[25];
    data_o[26] = (syndrome_o == 8'ha1) ^ data_i[26];
    data_o[27] = (syndrome_o == 8'ha2) ^ data_i[27];
    data_o[28] = (syndrome_o == 8'ha3) ^ data_i[28];
    data_o[29] = (syndrome_o == 8'ha4) ^ data_i[29];
    data_o[30] = (syndrome_o == 8'ha5) ^ data_i[30];
    data_o[31] = (syndrome_o == 8'ha6) ^ data_i[31];
    data_o[32] = (syndrome_o == 8'ha7) ^ data_i[32];
    data_o[33] = (syndrome_o == 8'ha8) ^ data_i[33];
    data_o[34] = (syndrome_o == 8'ha9) ^ data_i[34];
    data_o[35] = (syndrome_o == 8'haa) ^ data_i[35];
    data_o[36] = (syndrome_o == 8'hab) ^ data_i[36];
    data_o[37] = (syndrome_o == 8'hac) ^ data_i[37];
    data_o[38] = (syndrome_o == 8'had) ^ data_i[38];
    data_o[39] = (syndrome_o == 8'hae) ^ data_i[39];
    data_o[40] = (syndrome_o == 8'haf) ^ data_i[40];
    data_o[41] = (syndrome_o == 8'hb0) ^ data_i[41];
    data_o[42] = (syndrome_o == 8'hb1) ^ data_i[42];
    data_o[43] = (syndrome_o == 8'hb2) ^ data_i[43];
    data_o[44] = (syndrome_o == 8'hb3) ^ data_i[44];
    data_o[45] = (syndrome_o == 8'hb4) ^ data_i[45];
    data_o[46] = (syndrome_o == 8'hb5) ^ data_i[46];
    data_o[47] = (syndrome_o == 8'hb6) ^ data_i[47];
    data_o[48] = (syndrome_o == 8'hb7) ^ data_i[48];
    data_o[49] = (syndrome_o == 8'hb8) ^ data_i[49];
    data_o[50] = (syndrome_o == 8'hb9) ^ data_i[50];
    data_o[51] = (syndrome_o == 8'hba) ^ data_i[51];
    data_o[52] = (syndrome_o == 8'hbb) ^ data_i[52];
    data_o[53] = (syndrome_o == 8'hbc) ^ data_i[53];
    data_o[54] = (syndrome_o == 8'hbd) ^ data_i[54];
    data_o[55] = (syndrome_o == 8'hbe) ^ data_i[55];
    data_o[56] = (syndrome_o == 8'hbf) ^ data_i[56];
    data_o[57] = (syndrome_o == 8'hc1) ^ data_i[57];
    data_o[58] = (syndrome_o == 8'hc2) ^ data_i[58];
    data_o[59] = (syndrome_o == 8'hc3) ^ data_i[59];
    data_o[60] = (syndrome_o == 8'hc4) ^ data_i[60];
    data_o[61] = (syndrome_o == 8'hc5) ^ data_i[61];
    data_o[62] = (syndrome_o == 8'hc6) ^ data_i[62];
    data_o[63] = (syndrome_o == 8'hc7) ^ data_i[63];
    data_o[64] = (syndrome_o == 8'hc8) ^ data_i[64];
    data_o[65] = (syndrome_o == 8'hc9) ^ data_i[65];
    data_o[66] = (syndrome_o == 8'hca) ^ data_i[66];
    data_o[67] = (syndrome_o == 8'hcb) ^ data_i[67];

    // err_o calc. bit0: single error, bit1: double error
    err_o[0] = syndrome_o[7];
    err_o[1] = |syndrome_o[6:0] & ~syndrome_o[7];
  end
endmodule : prim_secded_inv_hamming_76_68_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SECDED encoder generated by util/design/secded_gen.py

module prim_secded_inv_hamming_76_68_enc (
  input        [67:0] data_i,
  output logic [75:0] data_o
);

  always_comb begin : p_encode
    data_o = 76'(data_i);
    data_o[68] = ^(data_o & 76'h00AAB55555556AAAD5B);
    data_o[69] = ^(data_o & 76'h00CCD9999999B33366D);
    data_o[70] = ^(data_o & 76'h000F1E1E1E1E3C3C78E);
    data_o[71] = ^(data_o & 76'h00F01FE01FE03FC07F0);
    data_o[72] = ^(data_o & 76'h00001FFFE0003FFF800);
    data_o[73] = ^(data_o & 76'h00001FFFFFFFC000000);
    data_o[74] = ^(data_o & 76'h00FFE00000000000000);
    data_o[75] = ^(data_o & 76'h7FFFFFFFFFFFFFFFFFF);
    data_o ^= 76'hAA00000000000000000;
  end

endmodule : prim_secded_inv_hamming_76_68_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_and2

#(

  parameter int Width = 1

) (
  input        [Width-1:0] in0_i,
  input        [Width-1:0] in1_i,
  output logic [Width-1:0] out_o
);

  if (1) begin : gen_generic
    prim_generic_and2 #(
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_buf

#(

  parameter int Width = 1

) (
  input        [Width-1:0] in_i,
  output logic [Width-1:0] out_o
);

  if (1) begin : gen_generic
    prim_generic_buf #(
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_flop

#(

  parameter int               Width      = 1,
  parameter logic [Width-1:0] ResetValue = 0

) (
  input                    clk_i,
  input                    rst_ni,
  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_o
);

  if (1) begin : gen_generic
    prim_generic_flop #(
      .ResetValue(ResetValue),
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_xnor2

#(

  parameter int Width = 1

) (
  input        [Width-1:0] in0_i,
  input        [Width-1:0] in1_i,
  output logic [Width-1:0] out_o
);

  if (1) begin : gen_generic
    prim_generic_xnor2 #(
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_xor2

#(

  parameter int Width = 1

) (
  input        [Width-1:0] in0_i,
  input        [Width-1:0] in1_i,
  output logic [Width-1:0] out_o
);

  if (1) begin : gen_generic
    prim_generic_xor2 #(
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// N:1 fixed priority arbiter module (index 0 has highest prio)
//
// Verilog parameter
//   N:           Number of request ports
//   DW:          Data width
//   DataPort:    Set to 1 to enable the data port. Otherwise that port will be ignored.
//
// See also: prim_arbiter_ppc, prim_arbiter_tree

`include "prim_assert.sv"

module prim_arbiter_fixed #(
  parameter int N   = 8,
  parameter int DW  = 32,

  // Configurations
  // EnDataPort: {0, 1}, if 0, input data will be ignored
  parameter bit EnDataPort = 1,

  // Derived parameters
  localparam int IdxW = $clog2(N)
) (
  // used for assertions only
  input clk_i,
  input rst_ni,

  input        [ N-1:0]    req_i,
  input        [DW-1:0]    data_i [N],
  output logic [ N-1:0]    gnt_o,
  output logic [IdxW-1:0]  idx_o,

  output logic             valid_o,
  output logic [DW-1:0]    data_o,
  input                    ready_i
);

  `ASSERT_INIT(CheckNGreaterZero_A, N > 0)

  // this case is basically just a bypass
  if (N == 1) begin : gen_degenerate_case

    assign valid_o  = req_i[0];
    assign data_o   = data_i[0];
    assign gnt_o[0] = valid_o & ready_i;
    assign idx_o    = '0;

  end else begin : gen_normal_case

    // align to powers of 2 for simplicity
    // a full binary tree with N levels has 2**N + 2**N-1 nodes
    logic [2**(IdxW+1)-2:0]           req_tree;
    logic [2**(IdxW+1)-2:0]           gnt_tree;
    logic [2**(IdxW+1)-2:0][IdxW-1:0] idx_tree;
    logic [2**(IdxW+1)-2:0][DW-1:0]   data_tree;

    for (genvar level = 0; level < IdxW+1; level++) begin : gen_tree
      //
      // level+1   C0   C1   <- "Base1" points to the first node on "level+1",
      //            \  /         these nodes are the children of the nodes one level below
      // level       Pa      <- "Base0", points to the first node on "level",
      //                         these nodes are the parents of the nodes one level above
      //
      // hence we have the following indices for the Pa, C0, C1 nodes:
      // Pa = 2**level     - 1 + offset       = Base0 + offset
      // C0 = 2**(level+1) - 1 + 2*offset     = Base1 + 2*offset
      // C1 = 2**(level+1) - 1 + 2*offset + 1 = Base1 + 2*offset + 1
      //
      localparam int Base0 = (2**level)-1;
      localparam int Base1 = (2**(level+1))-1;

      for (genvar offset = 0; offset < 2**level; offset++) begin : gen_level
        localparam int Pa = Base0 + offset;
        localparam int C0 = Base1 + 2*offset;
        localparam int C1 = Base1 + 2*offset + 1;

        // this assigns the gated interrupt source signals, their
        // corresponding IDs and priorities to the tree leafs
        if (level == IdxW) begin : gen_leafs
          if (offset < N) begin : gen_assign
            // forward path
            assign req_tree[Pa]      = req_i[offset];
            assign idx_tree[Pa]      = offset;
            assign data_tree[Pa]     = data_i[offset];
            // backward (grant) path
            assign gnt_o[offset]     = gnt_tree[Pa];

          end else begin : gen_tie_off
            // forward path
            assign req_tree[Pa]  = '0;
            assign idx_tree[Pa]  = '0;
            assign data_tree[Pa] = '0;
            logic unused_sigs;
            assign unused_sigs = gnt_tree[Pa];
          end
        // this creates the node assignments
        end else begin : gen_nodes
          // forward path
          logic sel; // local helper variable
          always_comb begin : p_node
            // this always gives priority to the left child
            sel = ~req_tree[C0];
            // propagate requests
            req_tree[Pa]  = req_tree[C0] | req_tree[C1];
            // data and index muxes
            idx_tree[Pa]  = (sel) ? idx_tree[C1]  : idx_tree[C0];
            data_tree[Pa] = (sel) ? data_tree[C1] : data_tree[C0];
            // propagate the grants back to the input
            gnt_tree[C0] = gnt_tree[Pa] & ~sel;
            gnt_tree[C1] = gnt_tree[Pa] &  sel;
          end
        end
      end : gen_level
    end : gen_tree

    // the results can be found at the tree root
    if (EnDataPort) begin : gen_data_port
      assign data_o      = data_tree[0];
    end else begin : gen_no_dataport
      logic [DW-1:0] unused_data;
      assign unused_data = data_tree[0];
      assign data_o = '1;
    end

    assign idx_o       = idx_tree[0];
    assign valid_o     = req_tree[0];

    // this propagates a grant back to the input
    assign gnt_tree[0] = valid_o & ready_i;
  end

  ////////////////
  // assertions //
  ////////////////

  // KNOWN assertions on outputs, except for data as that may be partially X in simulation
  // e.g. when used on a BUS
  `ASSERT_KNOWN(ValidKnown_A, valid_o)
  `ASSERT_KNOWN(GrantKnown_A, gnt_o)
  `ASSERT_KNOWN(IdxKnown_A, idx_o)

  // Make sure no higher prio req is asserted
  `ASSERT(Priority_A, |req_i |-> req_i[idx_o] && (((N'(1'b1) << idx_o) - 1'b1) & req_i) == '0)

  // we can only grant one requestor at a time
  `ASSERT(CheckHotOne_A, $onehot0(gnt_o))
  // A grant implies that the sink is ready
  `ASSERT(GntImpliesReady_A, |gnt_o |-> ready_i)
  // A grant implies that the arbiter asserts valid as well
  `ASSERT(GntImpliesValid_A, |gnt_o |-> valid_o)
  // A request and a sink that is ready imply a grant
  `ASSERT(ReqAndReadyImplyGrant_A, |req_i && ready_i |-> |gnt_o)
  // A request and a sink that is ready imply a grant
  `ASSERT(ReqImpliesValid_A, |req_i |-> valid_o)
  // Both conditions above combined and reversed
  `ASSERT(ReadyAndValidImplyGrant_A, ready_i && valid_o |-> |gnt_o)
  // Both conditions above combined and reversed
  `ASSERT(NoReadyValidNoGrant_A, !(ready_i || valid_o) |-> gnt_o == 0)
  // check index / grant correspond
  `ASSERT(IndexIsCorrect_A, ready_i && valid_o |-> gnt_o[idx_o] && req_i[idx_o])

if (EnDataPort) begin: gen_data_port_assertion
  // data flow
  `ASSERT(DataFlow_A, ready_i && valid_o |-> data_o == data_i[idx_o])
end

endmodule : prim_arbiter_fixed


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// N:1 arbiter module
//
// Verilog parameter
//   N:           Number of request ports
//   DW:          Data width
//   DataPort:    Set to 1 to enable the data port. Otherwise that port will be ignored.
//
// This is the original implementation of the arbiter which relies on parallel prefix computing
// optimization to optimize the request / arbiter tree. Not all synthesis tools may support this.
//
// Note that the currently winning request is held if the data sink is not ready. This behavior is
// required by some interconnect protocols (AXI, TL). The module contains an assertion that checks
// this behavior.
//
// Also, this module contains a request stability assertion that checks that requests stay asserted
// until they have been served. This assertion can be gated by driving the req_chk_i low. This is
// a non-functional input and does not affect the designs behavior.
//
// See also: prim_arbiter_tree

`include "prim_assert.sv"

module prim_arbiter_ppc #(
  parameter int unsigned N  = 8,
  parameter int unsigned DW = 32,

  // Configurations
  // EnDataPort: {0, 1}, if 0, input data will be ignored
  parameter bit EnDataPort = 1,

  // Derived parameters
  // localparam int IdxW = $clog2(N)
  // localparam int IdxW = 1
  parameter int IdxW = 1
) (
  input clk_i,
  input rst_ni,

  input                    req_chk_i, // Used for gating assertions. Drive to 1 during normal
                                      // operation.
  input        [ N-1:0]    req_i,
  input        [DW-1:0]    data_i [N],
  output logic [ N-1:0]    gnt_o,
  output logic [IdxW-1:0]  idx_o,

  output logic             valid_o,
  output logic [DW-1:0]    data_o,
  input                    ready_i
);

  // req_chk_i is used for gating assertions only.
  logic unused_req_chk;
  assign unused_req_chk = req_chk_i;

  `ASSERT_INIT(CheckNGreaterZero_A, N > 0)

  // this case is basically just a bypass
  if (N == 1) begin : gen_degenerate_case

    assign valid_o  = req_i[0];
    assign data_o   = data_i[0];
    assign gnt_o[0] = valid_o & ready_i;
    assign idx_o    = '0;

  end else begin : gen_normal_case

    logic [N-1:0] masked_req;
    logic [N-1:0] ppc_out;
    logic [N-1:0] arb_req;
    logic [N-1:0] mask, mask_next;
    logic [N-1:0] winner;

    assign masked_req = mask & req_i;
    assign arb_req = (|masked_req) ? masked_req : req_i;

    // PPC
    //   Even below code looks O(n) but DC optimizes it to O(log(N))
    //   Using Parallel Prefix Computation
    always_comb begin
      ppc_out[0] = arb_req[0];
      for (int i = 1 ; i < N ; i++) begin
        ppc_out[i] = ppc_out[i-1] | arb_req[i];
      end
    end

    // Grant Generation: Leading-One detector
    assign winner = ppc_out ^ {ppc_out[N-2:0], 1'b0};
    assign gnt_o    = (ready_i) ? winner : '0;

    assign valid_o = |req_i;
    // Mask Generation
    assign mask_next = {ppc_out[N-2:0], 1'b0};
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        mask <= '0;
      end else if (valid_o && ready_i) begin
        // Latch only when requests accepted
        mask <= mask_next;
      end else if (valid_o && !ready_i) begin
        // Downstream isn't yet ready so, keep current request alive. (First come first serve)
        mask <= ppc_out;
      end
    end

    if (EnDataPort == 1) begin: gen_datapath
      always_comb begin
        data_o = '0;
        for (int i = 0 ; i < N ; i++) begin
          if (winner[i]) begin
            data_o = data_i[i];
          end
        end
      end
    end else begin: gen_nodatapath
      assign data_o = '1;
      // The following signal is used to avoid possible lint errors.
      logic [DW-1:0] unused_data [N];
      assign unused_data = data_i;
    end

    always_comb begin
      idx_o = '0;
      for (int unsigned i = 0 ; i < N ; i++) begin
        if (winner[i]) begin
          idx_o = i[IdxW-1:0];
        end
      end
    end
  end

  ////////////////
  // assertions //
  ////////////////

  // KNOWN assertions on outputs, except for data as that may be partially X in simulation
  // e.g. when used on a BUS
  `ASSERT_KNOWN(ValidKnown_A, valid_o)
  `ASSERT_KNOWN(GrantKnown_A, gnt_o)
  `ASSERT_KNOWN(IdxKnown_A, idx_o)

  // grant index shall be higher index than previous index, unless no higher requests exist.
  `ASSERT(RoundRobin_A,
      ##1 valid_o && ready_i && $past(ready_i) && $past(valid_o) &&
      |(req_i & ~((N'(1) << $past(idx_o)+1) - 1)) |->
      idx_o > $past(idx_o))
  // we can only grant one requestor at a time
  `ASSERT(CheckHotOne_A, $onehot0(gnt_o))
  // A grant implies that the sink is ready
  `ASSERT(GntImpliesReady_A, |gnt_o |-> ready_i)
  // A grant implies that the arbiter asserts valid as well
  `ASSERT(GntImpliesValid_A, |gnt_o |-> valid_o)
  // A request and a sink that is ready imply a grant
  `ASSERT(ReqAndReadyImplyGrant_A, |req_i && ready_i |-> |gnt_o)
  // A request and a sink that is ready imply a grant
  `ASSERT(ReqImpliesValid_A, |req_i |-> valid_o)
  // Both conditions above combined and reversed
  `ASSERT(ReadyAndValidImplyGrant_A, ready_i && valid_o |-> |gnt_o)
  // Both conditions above combined and reversed
  `ASSERT(NoReadyValidNoGrant_A, !(ready_i || valid_o) |-> gnt_o == 0)
  // check index / grant correspond
  `ASSERT(IndexIsCorrect_A, ready_i && valid_o |-> gnt_o[idx_o] && req_i[idx_o])

if (EnDataPort) begin: gen_data_port_assertion
  // data flow
  `ASSERT(DataFlow_A, ready_i && valid_o |-> data_o == data_i[idx_o])
end

  // requests must stay asserted until they have been granted
  `ASSUME(ReqStaysHighUntilGranted0_M, |req_i && !ready_i |=>
      (req_i & $past(req_i)) == $past(req_i), clk_i, !rst_ni || !req_chk_i)
  // check that the arbitration decision is held if the sink is not ready
  `ASSERT(LockArbDecision_A, |req_i && !ready_i |=> idx_o == $past(idx_o),
      clk_i, !rst_ni || !req_chk_i)

// FPV-only assertions with symbolic variables
`ifdef FPV_ON
  // symbolic variables
  int unsigned k;
  bit ReadyIsStable;
  bit ReqsAreStable;

  // constraints for symbolic variables
  `ASSUME(KStable_M, ##1 $stable(k))
  `ASSUME(KRange_M, k < N)
  // this is used enable checking for stable and unstable ready_i and req_i signals in the same run.
  // the symbolic variables act like a switch that the solver can trun on and off.
  `ASSUME(ReadyIsStable_M, ##1 $stable(ReadyIsStable))
  `ASSUME(ReqsAreStable_M, ##1 $stable(ReqsAreStable))
  `ASSUME(ReadyStable_M, ##1 !ReadyIsStable || $stable(ready_i))
  `ASSUME(ReqsStable_M, ##1 !ReqsAreStable || $stable(req_i))

  // A grant implies a request
  `ASSERT(GntImpliesReq_A, gnt_o[k] |-> req_i[k])

  // if request and ready are constantly held at 1, we should eventually get a grant
  `ASSERT(NoStarvation_A,
      ReqsAreStable && ReadyIsStable && ready_i && req_i[k] |->
      strong(##[0:$] gnt_o[k]))

  // if N requests are constantly asserted and ready is constant 1, each request must
  // be granted exactly once over a time window of N cycles for the arbiter to be fair.
  for (genvar n = 1; n <= N; n++) begin : gen_fairness
    integer gnt_cnt;
    `ASSERT(Fairness_A,
        ReqsAreStable && ReadyIsStable && ready_i && req_i[k] &&
        $countones(req_i) == n |->
        ##n gnt_cnt == $past(gnt_cnt, n) + 1)

    always_ff @(posedge clk_i or negedge rst_ni) begin : p_cnt
      if (!rst_ni) begin
        gnt_cnt <= 0;
      end else begin
        gnt_cnt <= gnt_cnt + gnt_o[k];
      end
    end
  end

  // requests must stay asserted until they have been granted
  `ASSUME(ReqStaysHighUntilGranted1_M, req_i[k] && !gnt_o[k] |=>
      req_i[k], clk_i, !rst_ni || !req_chk_i)
`endif

endmodule : prim_arbiter_ppc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// N:1 arbiter module
//
// Verilog parameter
//   N:           Number of request ports
//   DW:          Data width
//   DataPort:    Set to 1 to enable the data port. Otherwise that port will be ignored.
//
// This is a tree implementation of a round robin arbiter. It has the same behavior as the PPC
// implementation in prim_arbiter_ppc, and also uses a prefix summing approach to determine the next
// request to be granted. The main difference with respect to the PPC arbiter is that the leading 1
// detection and the prefix summation are performed with a binary tree instead of a sequential loop.
// Also, if the data port is enabled, the data is muxed based on the local arbitration decisions  at
// each node of the arbiter tree. This means that the data can propagate through the tree
// simultaneously with the requests, instead of waiting for the arbitration to determine the winner
// index first. As a result, this design has a shorter critical path than other implementations,
// leading to better ovberall timing.
//
// Note that the currently winning request is held if the data sink is not ready. This behavior is
// required by some interconnect protocols (AXI, TL). The module contains an assertion that checks
// this behavior.
//
// Also, this module contains a request stability assertion that checks that requests stay asserted
// until they have been served. This assertion can be gated by driving the req_chk_i low. This is
// a non-functional input and does not affect the designs behavior.
//
// See also: prim_arbiter_ppc

`include "prim_assert.sv"

module prim_arbiter_tree #(
  parameter int N   = 8,
  parameter int DW  = 32,

  // Configurations
  // EnDataPort: {0, 1}, if 0, input data will be ignored
  parameter bit EnDataPort = 1,

  // Derived parameters
  localparam int IdxW = $clog2(N)
) (
  input clk_i,
  input rst_ni,

  input                    req_chk_i, // Used for gating assertions. Drive to 1 during normal
                                      // operation.
  input        [ N-1:0]    req_i,
  input        [DW-1:0]    data_i [N],
  output logic [ N-1:0]    gnt_o,
  output logic [IdxW-1:0]  idx_o,

  output logic             valid_o,
  output logic [DW-1:0]    data_o,
  input                    ready_i
);

  // req_chk_i is used for gating assertions only.
  logic unused_req_chk;
  assign unused_req_chk = req_chk_i;

  `ASSERT_INIT(CheckNGreaterZero_A, N > 0)

  // this case is basically just a bypass
  if (N == 1) begin : gen_degenerate_case

    assign valid_o  = req_i[0];
    assign data_o   = data_i[0];
    assign gnt_o[0] = valid_o & ready_i;
    assign idx_o    = '0;

  end else begin : gen_normal_case

    // align to powers of 2 for simplicity
    // a full binary tree with N levels has 2**N + 2**N-1 nodes
    logic [2**(IdxW+1)-2:0]           req_tree;
    logic [2**(IdxW+1)-2:0]           prio_tree;
    logic [2**(IdxW+1)-2:0]           sel_tree;
    logic [2**(IdxW+1)-2:0]           mask_tree;
    logic [2**(IdxW+1)-2:0][IdxW-1:0] idx_tree;
    logic [2**(IdxW+1)-2:0][DW-1:0]   data_tree;
    logic [N-1:0]                     prio_mask_d, prio_mask_q;

    for (genvar level = 0; level < IdxW+1; level++) begin : gen_tree
      //
      // level+1   C0   C1   <- "Base1" points to the first node on "level+1",
      //            \  /         these nodes are the children of the nodes one level below
      // level       Pa      <- "Base0", points to the first node on "level",
      //                         these nodes are the parents of the nodes one level above
      //
      // hence we have the following indices for the Pa, C0, C1 nodes:
      // Pa = 2**level     - 1 + offset       = Base0 + offset
      // C0 = 2**(level+1) - 1 + 2*offset     = Base1 + 2*offset
      // C1 = 2**(level+1) - 1 + 2*offset + 1 = Base1 + 2*offset + 1
      //
      localparam int Base0 = (2**level)-1;
      localparam int Base1 = (2**(level+1))-1;

      for (genvar offset = 0; offset < 2**level; offset++) begin : gen_level
        localparam int Pa = Base0 + offset;
        localparam int C0 = Base1 + 2*offset;
        localparam int C1 = Base1 + 2*offset + 1;

        // this assigns the gated interrupt source signals, their
        // corresponding IDs and priorities to the tree leafs
        if (level == IdxW) begin : gen_leafs
          if (offset < N) begin : gen_assign
            // forward path (requests and data)
            // all requests inputs are assigned to the request tree
            assign req_tree[Pa]      = req_i[offset];
            // we basically split the incoming request vector into two halves with the following
            // priority assignment. the prio_mask_q register contains a prefix sum that has been
            // computed using the last winning index, and hence masks out all requests at offsets
            // lower or equal the previously granted index. hence, all higher indices are considered
            // first in the arbitration tree nodes below, before considering the lower indices.
            assign prio_tree[Pa]     = req_i[offset] & prio_mask_q[offset];
            // input for the index muxes (used to compute the winner index)
            assign idx_tree[Pa]      = offset;
            // input for the data muxes
            assign data_tree[Pa]     = data_i[offset];

            // backward path (grants and prefix sum)
            // grant if selected, ready and request asserted
            assign gnt_o[offset]       = req_i[offset] & sel_tree[Pa] & ready_i;
            // only update mask if there is a valid request
            assign prio_mask_d[offset] = (|req_i) ?
                                         mask_tree[Pa] | sel_tree[Pa] & ~ready_i :
                                         prio_mask_q[offset];
          end else begin : gen_tie_off
            // forward path
            assign req_tree[Pa]  = '0;
            assign prio_tree[Pa] = '0;
            assign idx_tree[Pa]  = '0;
            assign data_tree[Pa] = '0;
            logic unused_sigs;
            assign unused_sigs = ^{mask_tree[Pa],
                                   sel_tree[Pa]};
          end
        // this creates the node assignments
        end else begin : gen_nodes
          // local helper variable
          logic sel;

          // forward path (requests and data)
          // each node looks at its two children, and selects the one with higher priority
          assign sel = ~req_tree[C0] | ~prio_tree[C0] & prio_tree[C1];
          // propagate requests
          assign req_tree[Pa]  = req_tree[C0] | req_tree[C1];
          assign prio_tree[Pa] = prio_tree[C1] | prio_tree[C0];
          // data and index muxes
          // Note: these ternaries have triggered a synthesis bug in Vivado versions older
          // than 2020.2. If the problem resurfaces again, have a look at issue #1408.
          assign idx_tree[Pa]  = (sel) ? idx_tree[C1]  : idx_tree[C0];
          assign data_tree[Pa] = (sel) ? data_tree[C1] : data_tree[C0];

          // backward path (grants and prefix sum)
          // this propagates the selction index back and computes a hot one mask
          assign sel_tree[C0] = sel_tree[Pa] & ~sel;
          assign sel_tree[C1] = sel_tree[Pa] &  sel;
          // this performs a prefix sum for masking the input requests in the next cycle
          assign mask_tree[C0] = mask_tree[Pa];
          assign mask_tree[C1] = mask_tree[Pa] | sel_tree[C0];
        end
      end : gen_level
    end : gen_tree

    // the results can be found at the tree root
    if (EnDataPort) begin : gen_data_port
      assign data_o      = data_tree[0];
    end else begin : gen_no_dataport
      logic [DW-1:0] unused_data;
      assign unused_data = data_tree[0];
      assign data_o = '1;
    end

    // This index is unused.
    logic unused_prio_tree;
    assign unused_prio_tree = prio_tree[0];

    assign idx_o       = idx_tree[0];
    assign valid_o     = req_tree[0];

    // the select tree computes a hot one signal that indicates which request is currently selected
    assign sel_tree[0] = 1'b1;
    // the mask tree is basically a prefix sum of the hot one select signal computed above
    assign mask_tree[0] = 1'b0;

    always_ff @(posedge clk_i or negedge rst_ni) begin : p_mask_reg
      if (!rst_ni) begin
        prio_mask_q <= '0;
      end else begin
        prio_mask_q <= prio_mask_d;
      end
    end
  end

  ////////////////
  // assertions //
  ////////////////

  // KNOWN assertions on outputs, except for data as that may be partially X in simulation
  // e.g. when used on a BUS
  `ASSERT_KNOWN(ValidKnown_A, valid_o)
  `ASSERT_KNOWN(GrantKnown_A, gnt_o)
  `ASSERT_KNOWN(IdxKnown_A, idx_o)

  // grant index shall be higher index than previous index, unless no higher requests exist.
  `ASSERT(RoundRobin_A,
      ##1 valid_o && ready_i && $past(ready_i) && $past(valid_o) &&
      |(req_i & ~((N'(1) << $past(idx_o)+1) - 1)) |->
      idx_o > $past(idx_o))
  // we can only grant one requestor at a time
  `ASSERT(CheckHotOne_A, $onehot0(gnt_o))
  // A grant implies that the sink is ready
  `ASSERT(GntImpliesReady_A, |gnt_o |-> ready_i)
  // A grant implies that the arbiter asserts valid as well
  `ASSERT(GntImpliesValid_A, |gnt_o |-> valid_o)
  // A request and a sink that is ready imply a grant
  `ASSERT(ReqAndReadyImplyGrant_A, |req_i && ready_i |-> |gnt_o)
  // A request and a sink that is ready imply a grant
  `ASSERT(ReqImpliesValid_A, |req_i |-> valid_o)
  // Both conditions above combined and reversed
  `ASSERT(ReadyAndValidImplyGrant_A, ready_i && valid_o |-> |gnt_o)
  // Both conditions above combined and reversed
  `ASSERT(NoReadyValidNoGrant_A, !(ready_i || valid_o) |-> gnt_o == 0)
  // check index / grant correspond
  `ASSERT(IndexIsCorrect_A, ready_i && valid_o |-> gnt_o[idx_o] && req_i[idx_o])

if (EnDataPort) begin: gen_data_port_assertion
  // data flow
  `ASSERT(DataFlow_A, ready_i && valid_o |-> data_o == data_i[idx_o])
end

  // requests must stay asserted until they have been granted
  `ASSUME(ReqStaysHighUntilGranted0_M, |req_i && !ready_i |=>
      (req_i & $past(req_i)) == $past(req_i), clk_i, !rst_ni || !req_chk_i)
  // check that the arbitration decision is held if the sink is not ready
  `ASSERT(LockArbDecision_A, |req_i && !ready_i |=> idx_o == $past(idx_o),
      clk_i, !rst_ni || !req_chk_i)

// FPV-only assertions with symbolic variables
`ifdef FPV_ON
  // symbolic variables
  int unsigned k;
  bit ReadyIsStable;
  bit ReqsAreStable;

  // constraints for symbolic variables
  `ASSUME(KStable_M, ##1 $stable(k))
  `ASSUME(KRange_M, k < N)
  // this is used enable checking for stable and unstable ready_i and req_i signals in the same run.
  // the symbolic variables act like a switch that the solver can trun on and off.
  `ASSUME(ReadyIsStable_M, ##1 $stable(ReadyIsStable))
  `ASSUME(ReqsAreStable_M, ##1 $stable(ReqsAreStable))
  `ASSUME(ReadyStable_M, ##1 !ReadyIsStable || $stable(ready_i))
  `ASSUME(ReqsStable_M, ##1 !ReqsAreStable || $stable(req_i))

  // A grant implies a request
  `ASSERT(GntImpliesReq_A, gnt_o[k] |-> req_i[k])

  // if request and ready are constantly held at 1, we should eventually get a grant
  `ASSERT(NoStarvation_A,
      ReqsAreStable && ReadyIsStable && ready_i && req_i[k] |->
      strong(##[0:$] gnt_o[k]))

  // if N requests are constantly asserted and ready is constant 1, each request must
  // be granted exactly once over a time window of N cycles for the arbiter to be fair.
  for (genvar n = 1; n <= N; n++) begin : gen_fairness
    integer gnt_cnt;
    `ASSERT(Fairness_A,
        ReqsAreStable && ReadyIsStable && ready_i && req_i[k] &&
        $countones(req_i) == n |->
        ##n gnt_cnt == $past(gnt_cnt, n) + 1)

    always_ff @(posedge clk_i or negedge rst_ni) begin : p_cnt
      if (!rst_ni) begin
        gnt_cnt <= 0;
      end else begin
        gnt_cnt <= gnt_cnt + gnt_o[k];
      end
    end
  end

  // requests must stay asserted until they have been granted
  `ASSUME(ReqStaysHighUntilGranted1_M, req_i[k] && !gnt_o[k] |=>
      req_i[k], clk_i, !rst_ni || !req_chk_i)
`endif

endmodule : prim_arbiter_tree


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This is a wrapper module that instantiates two prim_aribter_tree modules.
// The reason for two is similar to modules such as prim_count/prim_lfsr where
// we use spatial redundancy to ensure the arbitration results are not altered.
//
// Note there are limits to this check, as the inputs to the duplicated arbiter
// is still a single lane. So an upstream attack can defeat this module.  The
// duplication merely protects against attacks directly on the arbiter.

`include "prim_assert.sv"

module prim_arbiter_tree_dup #(
  parameter int N   = 8,
  parameter int DW  = 32,

  // Configurations
  // EnDataPort: {0, 1}, if 0, input data will be ignored
  parameter bit EnDataPort = 1,

  // if arbiter has fixed priority
  parameter bit FixedArb = 0,

  // Derived parameters
  localparam int IdxW = $clog2(N)
) (
  input clk_i,
  input rst_ni,

  input                    req_chk_i, // Used for gating assertions. Drive to 1 during normal
                                      // operation.
  input        [ N-1:0]    req_i,
  input        [DW-1:0]    data_i [N],
  output logic [ N-1:0]    gnt_o,
  output logic [IdxW-1:0]  idx_o,

  output logic             valid_o,
  output logic [DW-1:0]    data_o,
  input                    ready_i,
  output logic             err_o
);

  localparam int ArbInstances = 2;

  //typedef struct packed {
  //  logic [N-1:0] req;
  //  logic [N-1:0][DW-1:0] data;
  //} arb_inputs_t;

  typedef struct packed {
    logic valid;
    logic [N-1:0] gnt;
    logic [IdxW-1:0] idx;
    logic [DW-1:0] data;
  } arb_outputs_t;

  // buffer up the inputs separately for each instance
  //arb_inputs_t arb_in;
  //arb_inputs_t [ArbInstances-1:0] arb_input_buf;
  arb_outputs_t [ArbInstances-1:0] arb_output_buf;

  for (genvar i = 0; i < ArbInstances; i++) begin : gen_input_bufs
    logic [N-1:0] req_buf;
    prim_buf #(
      .Width(N)
    ) u_req_buf (
      .in_i(req_i),
      .out_o(req_buf)
    );

    logic [DW-1:0] data_buf [N];
    for (genvar j = 0; j < N; j++) begin : gen_data_bufs
      prim_buf #(
        .Width(DW)
      ) u_dat_buf (
        .in_i(data_i[j]),
        .out_o(data_buf[j])
      );
    end

    if (FixedArb) begin : gen_fixed_arbiter
      prim_arbiter_fixed  #(
        .N(N),
        .DW(DW),
        .EnDataPort(EnDataPort)
      ) u_arb (
        .clk_i,
        .rst_ni,
        .req_i(req_buf),
        .data_i(data_buf),
        .gnt_o(arb_output_buf[i].gnt),
        .idx_o(arb_output_buf[i].idx),
        .valid_o(arb_output_buf[i].valid),
        .data_o(arb_output_buf[i].data),
        .ready_i
      );
      logic unused_req_chk;
      assign unused_req_chk = req_chk_i;

    end else begin : gen_rr_arbiter
      prim_arbiter_tree #(
        .N(N),
        .DW(DW),
        .EnDataPort(EnDataPort)
      ) u_arb (
        .clk_i,
        .rst_ni,
        .req_chk_i,
        .req_i(req_buf),
        .data_i(data_buf),
        .gnt_o(arb_output_buf[i].gnt),
        .idx_o(arb_output_buf[i].idx),
        .valid_o(arb_output_buf[i].valid),
        .data_o(arb_output_buf[i].data),
        .ready_i
      );
    end
  end

  // the last buffered position is sent out
  assign gnt_o = arb_output_buf[ArbInstances-1].gnt;
  assign idx_o = arb_output_buf[ArbInstances-1].idx;
  assign valid_o = arb_output_buf[ArbInstances-1].valid;
  assign data_o = arb_output_buf[ArbInstances-1].data;

  // Check the last buffer index against all other instances
  logic [ArbInstances-2:0] output_delta;

  for (genvar i = 0; i < ArbInstances-1; i++) begin : gen_checks
    assign output_delta[i] = arb_output_buf[ArbInstances-1] != arb_output_buf[i];
  end

  logic err_d, err_q;
  // There is an error if anything ever disagrees
  assign err_d = |output_delta;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else begin
      err_q <= err_d | err_q;
    end
  end

  assign err_o = err_q;

endmodule // prim_arbiter_tree


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This module should be instantiated within flops of CDC synchronization primitives,
// and allows DV to model real CDC delays within simulations, especially useful at the chip level
// or in IPs that communicate across clock domains.
//
// The instrumentation is very simple: when this is enabled the input into the first
// synchronizer flop has a mux where the select is randomly set. One of the mux inputs is the input
// of this module, and the other is the output of the first flop: selecting the latter models the
// effect of the first flop missing the input transition.
//
// Notice the delay should cause the input to be skipped by at most a single cycle. As a perhaps
// unnecessary precaution, the select will only be allowed to be random when the input changes.

module prim_cdc_rand_delay #(
    parameter int DataWidth = 1,
    parameter bit Enable = 1
) (
    input logic                   clk_i,
    input logic                   rst_ni,
    input logic [DataWidth-1:0]   prev_data_i,
    input logic [DataWidth-1:0]   src_data_i,
    output logic [DataWidth-1:0]  dst_data_o
);
`ifdef SIMULATION
  if (Enable) begin : gen_enable

    // This controls dst_data_o: any bit with its data_sel set uses prev_data_i, others use
    // src_data_i.
    bit [DataWidth-1:0] data_sel;
    bit                 cdc_instrumentation_enabled;

    function automatic bit [DataWidth-1:0] fast_randomize();
      bit [DataWidth-1:0] data;
      if (DataWidth <= 32) begin
        data = $urandom();
      end else begin
        if (!std::randomize(data)) $fatal(1, "%t: [%m] Failed to randomize data", $time);
      end
      return data;
    endfunction

    initial begin
      void'($value$plusargs("cdc_instrumentation_enabled=%d", cdc_instrumentation_enabled));
      data_sel = '0;
    end

    // Set data_sel at random combinationally when the input changes.
    always @(src_data_i) begin
      data_sel = cdc_instrumentation_enabled ? fast_randomize() : 0;
    end

    // Clear data_del on any cycle start.
    always @(posedge clk_i or negedge rst_ni) begin
      data_sel <= 0;
    end

    always_comb dst_data_o = (prev_data_i & data_sel) | (src_data_i & ~data_sel);
  end else begin : gen_no_enable
    assign dst_data_o = src_data_i;
  end
`else  // SIMULATION
    assign dst_data_o = src_data_i;
`endif  // SIMULATION
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This is a simple data diffusion primitive that is constructed in a similar fashion
// as the PRESENT cipher (i.e. it uses a substitution/permutation network). Note however
// that this is **not** cryptographically secure. The main purpose of this primitive is to
// provide a cheap diffusion mechanism for arbitrarily sized vectors.
//
// See also: prim_prince, prim_present, prim_cipher_pkg

module prim_subst_perm #(
  parameter int DataWidth = 64,
  parameter int NumRounds = 31,
  parameter bit Decrypt   = 0    // 0: encrypt, 1: decrypt
) (
  input        [DataWidth-1:0] data_i,
  input        [DataWidth-1:0] key_i,
  output logic [DataWidth-1:0] data_o
);

  //////////////
  // datapath //
  //////////////

  // The "split_var" hint that we pass to verilator here tells it to schedule the different parts of
  // data_state separately. This avoids an UNOPTFLAT error where it would otherwise see a dependency
  // chain
  //
  //    data_state -> data_state_sbox -> data_state
  //
  logic [NumRounds:0][DataWidth-1:0] data_state /* verilator split_var */;

  // initialize
  assign data_state[0] = data_i;

  for (genvar r = 0; r < NumRounds; r++) begin : gen_round
    logic [DataWidth-1:0] data_state_sbox, data_state_flipped;
    ////////////////////////////////
    // decryption pass, performs inverse permutation and sbox
    if (Decrypt) begin : gen_dec
      always_comb begin : p_dec
        data_state_sbox = data_state[r] ^ key_i;
        // Reverse odd/even grouping
        data_state_flipped = data_state_sbox;
        for (int k = 0; k < DataWidth/2; k++) begin
          data_state_flipped[k * 2]     = data_state_sbox[k];
          data_state_flipped[k * 2 + 1] = data_state_sbox[k + DataWidth/2];
        end
        // Flip vector
        for (int k = 0; k < DataWidth; k++) begin
          data_state_sbox[DataWidth - 1 - k] = data_state_flipped[k];
        end
        // Inverse SBox layer
        for (int k = 0; k < DataWidth/4; k++) begin
          data_state_sbox[k*4 +: 4] = prim_cipher_pkg::PRESENT_SBOX4_INV[data_state_sbox[k*4 +: 4]];
        end
        data_state[r + 1] = data_state_sbox;
      end
    ////////////////////////////////
    // encryption pass
    end else begin : gen_enc
      always_comb begin : p_enc
        data_state_sbox = data_state[r] ^ key_i;
        // This SBox layer is aligned to nibbles, so the uppermost bits may not be affected by this.
        // However, the permutation below ensures that these bits get shuffled to a different
        // position when performing multiple rounds.
        for (int k = 0; k < DataWidth/4; k++) begin
          data_state_sbox[k*4 +: 4] = prim_cipher_pkg::PRESENT_SBOX4[data_state_sbox[k*4 +: 4]];
        end
        // Flip the vector to move the MSB positions into the LSB positions
        for (int k = 0; k < DataWidth; k++) begin
          data_state_flipped[DataWidth - 1 - k] = data_state_sbox[k];
        end
        // Regroup bits such that all even indices are stacked up first, followed by all odd
        // indices. Note that if the Width is odd, this is still ok, since
        // the uppermost bit just stays in place in that case.
        data_state_sbox = data_state_flipped;
        for (int k = 0; k < DataWidth/2; k++) begin
          data_state_sbox[k]               = data_state_flipped[k * 2];
          data_state_sbox[k + DataWidth/2] = data_state_flipped[k * 2 + 1];
        end
        data_state[r + 1] = data_state_sbox;
      end
    end // gen_enc
    ////////////////////////////////
  end // gen_round

  // finalize
  assign data_o = data_state[NumRounds] ^ key_i;

endmodule : prim_subst_perm


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module is an implementation of the encryption pass of the 64bit PRESENT
// block cipher. It is a fully unrolled combinational implementation that
// supports both key sizes specified in the paper (80bit and 128bit). Further,
// the number of rounds is fully configurable, and the primitive supports a
// 32bit block cipher flavor which is not specified in the original paper. It
// should be noted, however, that the 32bit version is **not** secure and must
// not be used in a setting where cryptographic cipher strength is required. The
// 32bit variant is only intended to be used as a lightweight data scrambling
// device.
//
// See also: prim_prince, prim_cipher_pkg
//
// References: - https://en.wikipedia.org/wiki/PRESENT
//             - https://en.wikipedia.org/wiki/Prince_(cipher)
//             - http://www.lightweightcrypto.org/present/present_ches2007.pdf
//             - https://eprint.iacr.org/2012/529.pdf
//             - https://csrc.nist.gov/csrc/media/events/lightweight-cryptography-workshop-2015/
//               documents/papers/session7-maene-paper.pdf

`include "prim_assert.sv"
module prim_present #(
  parameter int DataWidth = 64,  // {32, 64}
  parameter int KeyWidth  = 128, // {64, 80, 128}
  // Number of rounds to perform in total (>0)
  parameter int NumRounds = 31,
  // Number of physically instantiated PRESENT rounds.
  // This can be used to construct e.g. an iterative
  // full-round implementation that only has one physical
  // round instance by setting NumRounds = 31 and NumPhysRounds = 1.
  // Note that NumPhysRounds needs to divide NumRounds.
  parameter int NumPhysRounds = NumRounds,
  // Note that the decryption pass needs a modified key,
  // to be calculated by performing NumRounds key updates
  parameter bit Decrypt   = 0    // 0: encrypt, 1: decrypt
) (
  input        [DataWidth-1:0] data_i,
  input        [KeyWidth-1:0]  key_i,
  // Starting round index for keyschedule [1 ... 31].
  // Set this to 5'd1 for a fully unrolled encryption, and 5'd31 for a fully unrolled decryption.
  input        [4:0]           idx_i,
  output logic [DataWidth-1:0] data_o,
  output logic [KeyWidth-1:0]  key_o,
  // Next round index for keyschedule
  // (Enc: idx_i + NumPhysRounds, Dec: idx_i - NumPhysRounds)
  // Can be ignored for a fully unrolled implementation.
  output logic [4:0]           idx_o
);

  //////////////
  // datapath //
  //////////////

  logic [NumPhysRounds:0][DataWidth-1:0] data_state;
  logic [NumPhysRounds:0][KeyWidth-1:0]  round_key;
  logic [NumPhysRounds:0][4:0]           round_idx;

  // initialize
  assign data_state[0] = data_i;
  assign round_key[0]  = key_i;
  assign round_idx[0]  = idx_i;

  for (genvar k = 0; k < NumPhysRounds; k++) begin : gen_round
    logic [DataWidth-1:0] data_state_xor, data_state_sbox;
    // cipher layers
    assign data_state_xor  = data_state[k] ^ round_key[k][KeyWidth-1 : KeyWidth-DataWidth];
    ////////////////////////////////
    // decryption pass, performs inverse permutation, sbox and keyschedule
    if (Decrypt) begin : gen_dec
      // Decrement round count.
      assign round_idx[k+1] = round_idx[k] - 1'b1;
      // original 64bit variant
      if (DataWidth == 64) begin : gen_d64
        assign data_state_sbox = prim_cipher_pkg::perm_64bit(data_state_xor,
                                                             prim_cipher_pkg::PRESENT_PERM64_INV);
        assign data_state[k+1] = prim_cipher_pkg::sbox4_64bit(data_state_sbox,
                                                              prim_cipher_pkg::PRESENT_SBOX4_INV);
      // reduced 32bit variant
      end else begin : gen_d32
        assign data_state_sbox = prim_cipher_pkg::perm_32bit(data_state_xor,
                                                             prim_cipher_pkg::PRESENT_PERM32_INV);
        assign data_state[k+1] = prim_cipher_pkg::sbox4_32bit(data_state_sbox,
                                                              prim_cipher_pkg::PRESENT_SBOX4_INV);
      end
      // update round key, count goes from 1 to 31 (max)
      // original 128bit key variant
      if (KeyWidth == 128) begin : gen_k128
        assign round_key[k+1]  = prim_cipher_pkg::present_inv_update_key128(round_key[k],
                                                                            round_idx[k]);
      // original 80bit key variant
      end else if (KeyWidth == 80) begin : gen_k80
        assign round_key[k+1]  = prim_cipher_pkg::present_inv_update_key80(round_key[k],
                                                                           round_idx[k]);
      // reduced 64bit key variant
      end else begin : gen_k64
        assign round_key[k+1]  = prim_cipher_pkg::present_inv_update_key64(round_key[k],
                                                                           round_idx[k]);
      end
    ////////////////////////////////
    // encryption pass
    end else begin : gen_enc
      // Increment round count.
      assign round_idx[k+1] = round_idx[k] + 1'b1;
      // original 64bit variant
      if (DataWidth == 64) begin : gen_d64
        assign data_state_sbox = prim_cipher_pkg::sbox4_64bit(data_state_xor,
                                                              prim_cipher_pkg::PRESENT_SBOX4);
        assign data_state[k+1] = prim_cipher_pkg::perm_64bit(data_state_sbox,
                                                             prim_cipher_pkg::PRESENT_PERM64);
      // reduced 32bit variant
      end else begin : gen_d32
        assign data_state_sbox = prim_cipher_pkg::sbox4_32bit(data_state_xor,
                                                              prim_cipher_pkg::PRESENT_SBOX4);
        assign data_state[k+1] = prim_cipher_pkg::perm_32bit(data_state_sbox,
                                                             prim_cipher_pkg::PRESENT_PERM32);
      end
      // update round key, count goes from 1 to 31 (max)
      // original 128bit key variant
      if (KeyWidth == 128) begin : gen_k128
        assign round_key[k+1]  = prim_cipher_pkg::present_update_key128(round_key[k], round_idx[k]);
      // original 80bit key variant
      end else if (KeyWidth == 80) begin : gen_k80
        assign round_key[k+1]  = prim_cipher_pkg::present_update_key80(round_key[k], round_idx[k]);
      // reduced 64bit key variant
      end else begin : gen_k64
        assign round_key[k+1]  = prim_cipher_pkg::present_update_key64(round_key[k], round_idx[k]);
      end
    end // gen_enc
    ////////////////////////////////
  end // gen_round

  // This only needs to be applied after the last round.
  // Note that for a full-round implementation the output index
  // will be 0 for enc/dec for the last round (either due to wraparound or subtraction).
  localparam int LastRoundIdx = (Decrypt != 0 || NumRounds == 31) ? 0 : NumRounds+1;
  assign data_o = (int'(idx_o) == LastRoundIdx) ?
      data_state[NumPhysRounds] ^
      round_key[NumPhysRounds][KeyWidth-1 : KeyWidth-DataWidth] :
      data_state[NumPhysRounds];

  assign key_o  = round_key[NumPhysRounds];
  assign idx_o  = round_idx[NumPhysRounds];

  ////////////////
  // assertions //
  ////////////////

  `ASSERT_INIT(SupportedWidths_A, (DataWidth == 64 && KeyWidth inside {80, 128}) ||
                                  (DataWidth == 32 && KeyWidth == 64))
  `ASSERT_INIT(SupportedNumRounds_A, NumRounds > 0 && NumRounds <= 31)
  `ASSERT_INIT(SupportedNumPhysRounds0_A, NumPhysRounds > 0 && NumPhysRounds <= NumRounds)
  // Currently we do not support other arrangements
  `ASSERT_INIT(SupportedNumPhysRounds1_A, (NumRounds % NumPhysRounds) == 0)

endmodule : prim_present


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module is an implementation of the 64bit PRINCE block cipher. It is a fully unrolled
// combinational implementation with configurable number of rounds. Optionally, registers for the
// data and key states can be enabled, if this is required. Due to the reflective construction of
// this cipher, the same circuit can be used for encryption and decryption, as described below.
// Further, the primitive supports a 32bit block cipher flavor which is not specified in the
// original paper. It should be noted, however, that the 32bit version is **not** secure and must
// not be used in a setting where cryptographic cipher strength is required. The 32bit variant is
// only intended to be used as a lightweight data scrambling device.
//
// See also: prim_present, prim_cipher_pkg
//
// References: - https://en.wikipedia.org/wiki/PRESENT
//             - https://en.wikipedia.org/wiki/Prince_(cipher)
//             - http://www.lightweightcrypto.org/present/present_ches2007.pdf
//             - https://csrc.nist.gov/csrc/media/events/lightweight-cryptography-workshop-2015/
//               documents/papers/session7-maene-paper.pdf
//             - https://eprint.iacr.org/2012/529.pdf
//             - https://eprint.iacr.org/2015/372.pdf
//             - https://eprint.iacr.org/2014/656.pdf

`include "prim_assert.sv"
module prim_prince #(
  parameter int DataWidth     = 64,
  parameter int KeyWidth      = 128,
  // The construction is reflective. Total number of rounds is 2*NumRoundsHalf + 2
  parameter int NumRoundsHalf = 5,
  // This primitive uses the new key schedule proposed in https://eprint.iacr.org/2014/656.pdf
  // Setting this parameter to 1 falls back to the original key schedule.
  parameter bit UseOldKeySched = 1'b0,
  // This instantiates a data register halfway in the primitive.
  parameter bit HalfwayDataReg = 1'b0,
  // This instantiates a key register halfway in the primitive.
  parameter bit HalfwayKeyReg = 1'b0
) (
  input                        clk_i,
  input                        rst_ni,

  input                        valid_i,
  input        [DataWidth-1:0] data_i,
  input        [KeyWidth-1:0]  key_i,
  input                        dec_i,   // set to 1 for decryption
  output logic                 valid_o,
  output logic [DataWidth-1:0] data_o
);

  ///////////////////
  // key expansion //
  ///////////////////

  logic [DataWidth-1:0] k0, k0_prime_d, k1_d, k0_new_d, k0_prime_q, k1_q, k0_new_q;
  always_comb begin : p_key_expansion
    k0         = key_i[2*DataWidth-1 : DataWidth];
    k0_prime_d = {k0[0], k0[DataWidth-1:2], k0[DataWidth-1] ^ k0[1]};
    k1_d       = key_i[DataWidth-1:0];

    // modify key for decryption
    if (dec_i) begin
      k0          = k0_prime_d;
      k0_prime_d  = key_i[2*DataWidth-1 : DataWidth];
      k1_d       ^= prim_cipher_pkg::PRINCE_ALPHA_CONST[DataWidth-1:0];
    end
  end

  if (UseOldKeySched) begin : gen_legacy_keyschedule
    // In this case we constantly use k1.
    assign k0_new_d = k1_d;
  end else begin : gen_new_keyschedule
    // Imroved keyschedule proposed by https://eprint.iacr.org/2014/656.pdf
    // In this case we alternate between k1 and k0.
    always_comb begin : p_new_keyschedule_k0_alpha
      k0_new_d = key_i[2*DataWidth-1 : DataWidth];
      // We need to apply the alpha constant here as well, just as for k1 in decryption mode.
      if (dec_i) begin
        k0_new_d ^= prim_cipher_pkg::PRINCE_ALPHA_CONST[DataWidth-1:0];
      end
    end
  end

  if (HalfwayKeyReg) begin : gen_key_reg
    always_ff @(posedge clk_i or negedge rst_ni) begin : p_key_reg
      if (!rst_ni) begin
        k1_q       <= '0;
        k0_prime_q <= '0;
        k0_new_q   <= '0;
      end else begin
        if (valid_i) begin
          k1_q       <= k1_d;
          k0_prime_q <= k0_prime_d;
          k0_new_q   <= k0_new_d;
        end
      end
    end
  end else begin : gen_no_key_reg
    // just pass the key through in this case
    assign k1_q       = k1_d;
    assign k0_prime_q = k0_prime_d;
    assign k0_new_q   = k0_new_d;
  end

  //////////////
  // datapath //
  //////////////

  // State variable for holding the rounds
  logic [NumRoundsHalf:0][DataWidth-1:0] data_state_lo;
  logic [NumRoundsHalf:0][DataWidth-1:0] data_state_hi;

  // pre-round XOR
  always_comb begin : p_pre_round_xor
    data_state_lo[0] = data_i ^ k0;
    data_state_lo[0] ^= k1_d;
    data_state_lo[0] ^= prim_cipher_pkg::PRINCE_ROUND_CONST[0][DataWidth-1:0];
  end

  // forward pass
  for (genvar k = 1; k <= NumRoundsHalf; k++) begin : gen_fwd_pass
    logic [DataWidth-1:0] data_state_round;
    if (DataWidth == 64) begin : gen_fwd_d64
      always_comb begin : p_fwd_d64
        data_state_round = prim_cipher_pkg::sbox4_64bit(data_state_lo[k-1],
            prim_cipher_pkg::PRINCE_SBOX4);
        data_state_round = prim_cipher_pkg::prince_mult_prime_64bit(data_state_round);
        data_state_round = prim_cipher_pkg::prince_shiftrows_64bit(data_state_round,
            prim_cipher_pkg::PRINCE_SHIFT_ROWS64);
      end
    end else begin : gen_fwd_d32
      always_comb begin : p_fwd_d32
        data_state_round = prim_cipher_pkg::sbox4_32bit(data_state_lo[k-1],
            prim_cipher_pkg::PRINCE_SBOX4);
        data_state_round = prim_cipher_pkg::prince_mult_prime_32bit(data_state_round);
        data_state_round = prim_cipher_pkg::prince_shiftrows_32bit(data_state_round,
            prim_cipher_pkg::PRINCE_SHIFT_ROWS64);
      end
    end
    logic [DataWidth-1:0] data_state_xor;
    assign data_state_xor = data_state_round ^
                            prim_cipher_pkg::PRINCE_ROUND_CONST[k][DataWidth-1:0];
    // improved keyschedule proposed by https://eprint.iacr.org/2014/656.pdf
    if (k % 2 == 1) begin : gen_fwd_key_odd
      assign data_state_lo[k]  = data_state_xor ^ k0_new_d;
    end else begin : gen_fwd_key_even
      assign data_state_lo[k]  = data_state_xor ^ k1_d;
    end
  end

  // middle part
  logic [DataWidth-1:0] data_state_middle_d, data_state_middle_q, data_state_middle;
  if (DataWidth == 64) begin : gen_middle_d64
    always_comb begin : p_middle_d64
      data_state_middle_d = prim_cipher_pkg::sbox4_64bit(data_state_lo[NumRoundsHalf],
          prim_cipher_pkg::PRINCE_SBOX4);
      data_state_middle = prim_cipher_pkg::prince_mult_prime_64bit(data_state_middle_q);
      data_state_middle = prim_cipher_pkg::sbox4_64bit(data_state_middle,
          prim_cipher_pkg::PRINCE_SBOX4_INV);
    end
  end else begin : gen_middle_d32
    always_comb begin : p_middle_d32
      data_state_middle_d = prim_cipher_pkg::sbox4_32bit(data_state_middle[NumRoundsHalf],
          prim_cipher_pkg::PRINCE_SBOX4);
      data_state_middle = prim_cipher_pkg::prince_mult_prime_32bit(data_state_middle_q);
      data_state_middle = prim_cipher_pkg::sbox4_32bit(data_state_middle,
          prim_cipher_pkg::PRINCE_SBOX4_INV);
    end
  end

  if (HalfwayDataReg) begin : gen_data_reg
    logic valid_q;
    always_ff @(posedge clk_i or negedge rst_ni) begin : p_data_reg
      if (!rst_ni) begin
        valid_q <= 1'b0;
        data_state_middle_q <= '0;
      end else begin
        valid_q <= valid_i;
        if (valid_i) begin
          data_state_middle_q <= data_state_middle_d;
        end
      end
    end
    assign valid_o = valid_q;
  end else begin : gen_no_data_reg
    // just pass data through in this case
    assign data_state_middle_q = data_state_middle_d;
    assign valid_o = valid_i;
  end

  assign data_state_hi[0] = data_state_middle;

  // backward pass
  for (genvar k = 1; k <= NumRoundsHalf; k++) begin : gen_bwd_pass
    logic [DataWidth-1:0] data_state_xor0, data_state_xor1;
    // improved keyschedule proposed by https://eprint.iacr.org/2014/656.pdf
    if ((NumRoundsHalf + k + 1) % 2 == 1) begin : gen_bkwd_key_odd
      assign data_state_xor0 = data_state_hi[k-1] ^ k0_new_q;
    end else begin : gen_bkwd_key_even
      assign data_state_xor0 = data_state_hi[k-1] ^ k1_q;
    end
    // the construction is reflective, hence the subtraction with NumRoundsHalf
    assign data_state_xor1 = data_state_xor0 ^
                             prim_cipher_pkg::PRINCE_ROUND_CONST[10-NumRoundsHalf+k][DataWidth-1:0];

    logic [DataWidth-1:0] data_state_bwd;
    if (DataWidth == 64) begin : gen_bwd_d64
      always_comb begin : p_bwd_d64
        data_state_bwd = prim_cipher_pkg::prince_shiftrows_64bit(data_state_xor1,
            prim_cipher_pkg::PRINCE_SHIFT_ROWS64_INV);
        data_state_bwd = prim_cipher_pkg::prince_mult_prime_64bit(data_state_bwd);
        data_state_hi[k] = prim_cipher_pkg::sbox4_64bit(data_state_bwd,
            prim_cipher_pkg::PRINCE_SBOX4_INV);
      end
    end else begin : gen_bwd_d32
      always_comb begin : p_bwd_d32
        data_state_bwd = prim_cipher_pkg::prince_shiftrows_32bit(data_state_xor1,
            prim_cipher_pkg::PRINCE_SHIFT_ROWS64_INV);
        data_state_bwd = prim_cipher_pkg::prince_mult_prime_32bit(data_state_bwd);
        data_state_hi[k] = prim_cipher_pkg::sbox4_32bit(data_state_bwd,
            prim_cipher_pkg::PRINCE_SBOX4_INV);
      end
    end
  end

  // post-rounds
  always_comb begin : p_post_round_xor
    data_o  = data_state_hi[NumRoundsHalf] ^
              prim_cipher_pkg::PRINCE_ROUND_CONST[11][DataWidth-1:0];
    data_o ^= k1_q;
    data_o ^= k0_prime_q;
  end

  ////////////////
  // assertions //
  ////////////////

  `ASSERT_INIT(SupportedWidths_A, (DataWidth == 64 && KeyWidth == 128) ||
                                  (DataWidth == 32 && KeyWidth == 64))
  `ASSERT_INIT(SupportedNumRounds_A, NumRoundsHalf > 0 && NumRoundsHalf < 6)


endmodule : prim_prince


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Hardened counter primitive:
//
// This internally uses a cross counter scheme with primary and a secondary counter, where the
// secondary counter counts in reverse direction. The sum of both counters must remain constant and
// equal to 2**Width-1 or otherwise an err_o will be asserted.
//
// This counter supports a generic clear / set / increment / decrement interface:
//
// clr_i: This clears the primary counter to ResetValue and adjusts the secondary counter to match
//        (i.e. 2**Width-1-ResetValue). Clear has priority over set, increment and decrement.
// set_i: This sets the primary counter to set_cnt_i and adjusts the secondary counter to match
//        (i.e. 2**Width-1-set_cnt_i). Set has priority over increment and decrement.
// incr_en_i: Increments the primary counter by step_i, and decrements the secondary by step_i.
// decr_en_i: Decrements the primary counter by step_i, and increments the secondary by step_i.
//
// Note that if both incr_en_i and decr_en_i are asserted at the same time, the counter remains
// unchanged. The counter is also protected against under- and overflows.

`include "prim_assert.sv"

module prim_count #(
  parameter int Width = 2,
  // Can be used to reset the counter to a different value than 0, for example when
  // the counter is used as a down-counter.
  parameter logic [Width-1:0] ResetValue = '0,
  // This should only be disabled in special circumstances, for example
  // in non-comportable IPs where an error does not trigger an alert.
  parameter bit EnableAlertTriggerSVA = 1
) (
  input clk_i,
  input rst_ni,
  input clr_i,
  input set_i,
  input [Width-1:0] set_cnt_i,         // Set value for the counter.
  input incr_en_i,
  input decr_en_i,
  input [Width-1:0] step_i,            // Increment/decrement step when enabled.
  output logic [Width-1:0] cnt_o,      // Current counter state
  output logic [Width-1:0] cnt_next_o, // Next counter state
  output logic err_o
);

  ///////////////////
  // Counter logic //
  ///////////////////

  // Reset Values for primary and secondary counters.
  localparam int NumCnt = 2;
  localparam logic [NumCnt-1:0][Width-1:0] ResetValues = {{Width{1'b1}} - ResetValue, // secondary
                                                          ResetValue};                // primary

  logic [NumCnt-1:0][Width-1:0] cnt_d, cnt_q, fpv_force;

`ifndef FPV_SEC_CM_ON
  // This becomes a free variable in FPV.
  assign fpv_force = '0;
`endif

  for (genvar k = 0; k < NumCnt; k++) begin : gen_cnts
    // Note that increments / decrements are reversed for the secondary counter.
    logic incr_en, decr_en;
    logic [Width-1:0] set_val;
    if (k == 0) begin : gen_up_cnt
      assign incr_en = incr_en_i;
      assign decr_en = decr_en_i;
      assign set_val = set_cnt_i;
    end else begin : gen_dn_cnt
      assign incr_en = decr_en_i;
      assign decr_en = incr_en_i;
      // The secondary value needs to be adjusted accordingly.
      assign set_val = {Width{1'b1}} - set_cnt_i;
    end

    // Main counter logic
    logic [Width:0] ext_cnt;
    assign ext_cnt = (decr_en) ? {1'b0, cnt_q[k]} - {1'b0, step_i} :
                     (incr_en) ? {1'b0, cnt_q[k]} + {1'b0, step_i} : {1'b0, cnt_q[k]};

    // Saturation logic
    logic uflow, oflow;
    assign oflow = incr_en && ext_cnt[Width];
    assign uflow = decr_en && ext_cnt[Width];
    logic [Width-1:0] cnt_sat;
    assign cnt_sat = (uflow) ? '0            :
                     (oflow) ? {Width{1'b1}} : ext_cnt[Width-1:0];

    // Clock gate flops when in saturation, and do not
    // count if both incr_en and decr_en are asserted.
    logic cnt_en;
    assign cnt_en = (incr_en ^ decr_en) &&
                    ((incr_en && !(&cnt_q[k])) ||
                    (decr_en && !(cnt_q[k] == '0)));

    // Counter muxes
    assign cnt_d[k] = (clr_i)  ? ResetValues[k] :
                      (set_i)  ? set_val        :
                      (cnt_en) ? cnt_sat        : cnt_q[k];

    logic [Width-1:0] cnt_unforced_q;
    prim_flop #(
      .Width(Width),
      .ResetValue(ResetValues[k])
    ) u_cnt_flop (
      .clk_i,
      .rst_ni,
      .d_i(cnt_d[k]),
      .q_o(cnt_unforced_q)
    );

    // fpv_force is only used during FPV.
    assign cnt_q[k] = fpv_force[k] + cnt_unforced_q;
  end

  // The sum of both counters must always equal the counter maximum.
  logic [Width:0] sum;
  assign sum = (cnt_q[0] + cnt_q[1]);
  assign err_o = (sum != {1'b0, {Width{1'b1}}});

  // Output count values
  assign cnt_o      = cnt_q[0];
  assign cnt_next_o = cnt_d[0];

  ////////////////
  // Assertions //
  ////////////////
`ifdef INC_ASSERT
  //VCS coverage off
  // pragma coverage off

  // We need to disable most assertions in that case using a helper signal.
  // We can't rely on err_o since some error patterns cannot be detected (e.g. all error
  // patterns that still fullfill the sum constraint).
  logic fpv_err_present;
  assign fpv_err_present = |fpv_force;

  // Helper functions for assertions.
  function automatic logic signed [Width+1:0] max(logic signed [Width+1:0] a,
                                                  logic signed [Width+1:0] b);
    return (a > b) ? a : b;
  endfunction

  function automatic logic signed [Width+1:0] min(logic signed [Width+1:0] a,
                                                  logic signed [Width+1:0] b);
    return (a < b) ? a : b;
  endfunction
  //VCS coverage on
  // pragma coverage on

  // Cnt next
  `ASSERT(CntNext_A,
      rst_ni
      |=>
      cnt_o == $past(cnt_next_o),
      clk_i, err_o || fpv_err_present || !rst_ni)

  // Clear
  `ASSERT(ClrFwd_A,
      rst_ni && clr_i
      |=>
      (cnt_o == ResetValue) &&
      (cnt_q[1] == ({Width{1'b1}} - ResetValue)),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(ClrBkwd_A,
      rst_ni && !(incr_en_i || decr_en_i || set_i) ##1
      $changed(cnt_o) && $changed(cnt_q[1])
      |->
      $past(clr_i),
      clk_i, err_o || fpv_err_present || !rst_ni)

  // Set
  `ASSERT(SetFwd_A,
      rst_ni && set_i && !clr_i
      |=>
      (cnt_o == $past(set_cnt_i)) &&
      (cnt_q[1] == ({Width{1'b1}} - $past(set_cnt_i))),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(SetBkwd_A,
      rst_ni && !(incr_en_i || decr_en_i || clr_i) ##1
      $changed(cnt_o) && $changed(cnt_q[1])
      |->
      $past(set_i),
      clk_i, err_o || fpv_err_present || !rst_ni)

  // Do not count if both increment and decrement are asserted.
  `ASSERT(IncrDecrUpDnCnt_A,
      rst_ni && incr_en_i && decr_en_i && !(clr_i || set_i)
      |=>
      $stable(cnt_o) && $stable(cnt_q[1]),
      clk_i, err_o || fpv_err_present || !rst_ni)

  // Up counter
  `ASSERT(IncrUpCnt_A,
      rst_ni && incr_en_i && !(clr_i || set_i || decr_en_i)
      |=>
      cnt_o == min($past(cnt_o) + $past({2'b0, step_i}), {2'b0, {Width{1'b1}}}),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(IncrDnCnt_A,
      rst_ni && incr_en_i && !(clr_i || set_i || decr_en_i)
      |=>
      cnt_q[1] == max($past(signed'({2'b0, cnt_q[1]})) - $past({2'b0, step_i}), '0),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(UpCntIncrStable_A,
      incr_en_i && !(clr_i || set_i || decr_en_i) &&
      cnt_o == {Width{1'b1}}
      |=>
      $stable(cnt_o),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(UpCntDecrStable_A,
      decr_en_i && !(clr_i || set_i || incr_en_i) &&
      cnt_o == '0
      |=>
      $stable(cnt_o),
      clk_i, err_o || fpv_err_present || !rst_ni)

  // Down counter
  `ASSERT(DecrUpCnt_A,
      rst_ni && decr_en_i && !(clr_i || set_i || incr_en_i)
      |=>
      cnt_o == max($past(signed'({2'b0, cnt_o})) - $past({2'b0, step_i}), '0),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(DecrDnCnt_A,
      rst_ni && decr_en_i && !(clr_i || set_i || incr_en_i)
      |=>
      cnt_q[1] == min($past(cnt_q[1]) + $past({2'b0, step_i}), {2'b0, {Width{1'b1}}}),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(DnCntIncrStable_A,
      rst_ni && incr_en_i && !(clr_i || set_i || decr_en_i) &&
      cnt_q[1] == '0
      |=>
      $stable(cnt_q[1]),
      clk_i, err_o || fpv_err_present || !rst_ni)
  `ASSERT(DnCntDecrStable_A,
      rst_ni && decr_en_i && !(clr_i || set_i || incr_en_i) &&
      cnt_q[1] == {Width{1'b1}}
      |=>
      $stable(cnt_q[1]),
      clk_i, err_o || fpv_err_present || !rst_ni)

  // Error
  `ASSERT(CntErrForward_A,
      (cnt_q[1] + cnt_q[0]) != {Width{1'b1}}
      |->
      err_o)
  `ASSERT(CntErrBackward_A,
      err_o
      |->
      (cnt_q[1] + cnt_q[0]) != {Width{1'b1}})

  // This logic that will be assign to one, when user adds macro
  // ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT to check the error with alert, in case that prim_count
  // is used in design without adding this assertion check.
  logic unused_assert_connected;

  `ASSERT_INIT_NET(AssertConnected_A, unused_assert_connected === 1'b1 || !EnableAlertTriggerSVA)
`endif

endmodule // prim_count


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_clock_mux2 #(
  parameter bit NoFpgaBufG = 1'b0 // this parameter serves no function in the generic model
) (
  input        clk0_i,
  input        clk1_i,
  input        sel_i,
  output logic clk_o
);

  // We model the mux with logic operations for GTECH runs.
  assign clk_o = (sel_i & clk1_i) | (~sel_i & clk0_i);

  // make sure sel is never X (including during reset)
  // need to use ##1 as this could break with inverted clocks that
  // start with a rising edge at the beginning of the simulation.
  `ASSERT(selKnown0, ##1 !$isunknown(sel_i), clk0_i, 0)
  `ASSERT(selKnown1, ##1 !$isunknown(sel_i), clk1_i, 0)

endmodule : prim_generic_clock_mux2


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Generic, technology independent pad wrapper. This is NOT synthesizable!


`include "prim_assert.sv"

module prim_generic_pad_wrapper
  import prim_pad_wrapper_pkg::*;
#(
  // These parameters are ignored in this model.
  parameter pad_type_e PadType = BidirStd,
  parameter scan_role_e ScanRole = NoScan
) (
  // This is only used for scanmode (not used in generic models)
  input              clk_scan_i,
  input              scanmode_i,
  // Power sequencing signals (not used in generic models)
  input pad_pok_t    pok_i,
  // Main Pad signals
  inout wire         inout_io, // bidirectional pad
  output logic       in_o,     // input data
  output logic       in_raw_o, // uninverted output data
  input              ie_i,     // input enable
  input              out_i,    // output data
  input              oe_i,     // output enable
  input pad_attr_t   attr_i    // additional pad attributes
);

  // analog pads cannot have a scan role.
  `ASSERT_INIT(AnalogNoScan_A, PadType != AnalogIn0 || ScanRole == NoScan)

  //VCS coverage off
  // pragma coverage off
  // not all signals are used here.
  logic unused_sigs;
  assign unused_sigs = ^{attr_i.slew_rate,
                         attr_i.drive_strength[3:1],
                         attr_i.od_en,
                         attr_i.schmitt_en,
                         attr_i.keep_en,
                         scanmode_i,
                         pok_i};
  //VCS coverage on
  // pragma coverage on

  if (PadType == InputStd) begin : gen_input_only
    //VCS coverage off
    // pragma coverage off
    logic unused_in_sigs;
    assign unused_in_sigs = ^{out_i,
                              oe_i,
                              attr_i.virt_od_en,
                              attr_i.drive_strength};
    //VCS coverage on
    // pragma coverage on

    assign in_raw_o = (ie_i) ? inout_io  : 1'bz;
    // input inversion
    assign in_o = attr_i.invert ^ in_raw_o;

  // pulls are not supported by verilator
  `ifndef VERILATOR
    // pullup / pulldown termination
    assign (weak0, weak1) inout_io = attr_i.pull_en ? attr_i.pull_select : 1'bz;
  `endif
  end else if (PadType == BidirTol ||
               PadType == DualBidirTol ||
               PadType == BidirOd ||
               PadType == BidirStd) begin : gen_bidir

    assign in_raw_o = (ie_i) ? inout_io  : 1'bz;
    // input inversion
    assign in_o = attr_i.invert ^ in_raw_o;

    // virtual open drain emulation
    logic oe, out;
    assign out = out_i ^ attr_i.invert;
    assign oe  = oe_i & ((attr_i.virt_od_en & ~out) | ~attr_i.virt_od_en);

  // drive strength attributes are not supported by verilator
  `ifdef VERILATOR
    assign inout_io = (oe)   ? out : 1'bz;
  `else
    // different driver types
    assign (strong0, strong1) inout_io = (oe && attr_i.drive_strength[0]) ? out : 1'bz;
    assign (pull0, pull1)     inout_io = (oe && !attr_i.drive_strength[0]) ? out : 1'bz;
    // pullup / pulldown termination
    assign (weak0, weak1)     inout_io = attr_i.pull_en ? attr_i.pull_select : 1'bz;
  `endif
  end else if (PadType == AnalogIn0 || PadType == AnalogIn1) begin : gen_analog

    //VCS coverage off
    // pragma coverage off
    logic unused_ana_sigs;
    assign unused_ana_sigs = ^{attr_i, out_i, oe_i, ie_i};
    //VCS coverage on
    // pragma coverage on

    assign inout_io = 1'bz; // explicitly make this tristate to avoid lint errors.
    assign in_o = inout_io;
    assign in_raw_o = inout_io;

  end else begin : gen_invalid_config
    // this should throw link warnings in elaboration
    assert_static_in_generate_config_not_available
        assert_static_in_generate_config_not_available();
  end

endmodule : prim_generic_pad_wrapper


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Synchronous single-port SRAM model

`include "prim_assert.sv"

module prim_generic_ram_1p import prim_ram_1p_pkg::*; #(
  parameter  int Width           = 32, // bit
  parameter  int Depth           = 128,
  parameter  int DataBitsPerMask = 1, // Number of data bits per bit of write mask
  parameter      MemInitFile     = "", // VMEM file to initialize the memory with

  localparam int Aw              = $clog2(Depth)  // derived parameter
) (
  input  logic             clk_i,

  input  logic             req_i,
  input  logic             write_i,
  input  logic [Aw-1:0]    addr_i,
  input  logic [Width-1:0] wdata_i,
  input  logic [Width-1:0] wmask_i,
  output logic [Width-1:0] rdata_o, // Read data. Data is returned one cycle after req_i is high.
  input ram_1p_cfg_t       cfg_i
);

// For certain synthesis experiments we compile the design with generic models to get an unmapped
// netlist (GTECH). In these synthesis experiments, we typically black-box the memory models since
// these are going to be simulated using plain RTL models in netlist simulations. This can be done
// by analyzing and elaborating the design, and then removing the memory submodules before writing
// out the verilog netlist. However, memory arrays can take a long time to elaborate, and in case
// of dual port rams they can even trigger elab errors due to multiple processes writing to the
// same memory variable concurrently. To this end, we exclude the entire logic in this module in
// these runs with the following macro.
`ifndef SYNTHESIS_MEMORY_BLACK_BOXING

  // Width must be fully divisible by DataBitsPerMask
  `ASSERT_INIT(DataBitsPerMaskCheck_A, (Width % DataBitsPerMask) == 0)

  logic unused_cfg;
  assign unused_cfg = ^cfg_i;

  // Width of internal write mask. Note wmask_i input into the module is always assumed
  // to be the full bit mask
  localparam int MaskWidth = Width / DataBitsPerMask;

  logic [Width-1:0]     mem [Depth];
  logic [MaskWidth-1:0] wmask;

  for (genvar k = 0; k < MaskWidth; k++) begin : gen_wmask
    assign wmask[k] = &wmask_i[k*DataBitsPerMask +: DataBitsPerMask];

    // Ensure that all mask bits within a group have the same value for a write
    `ASSERT(MaskCheck_A, req_i && write_i |->
        wmask_i[k*DataBitsPerMask +: DataBitsPerMask] inside {{DataBitsPerMask{1'b1}}, '0},
        clk_i, '0)
  end

  // using always instead of always_ff to avoid 'ICPD  - illegal combination of drivers' error
  // thrown when using $readmemh system task to backdoor load an image
  // always @(posedge clk_i) begin
  //   if (req_i) begin
  //     if (write_i) begin
  //       for (int i=0; i < MaskWidth; i = i + 1) begin
  //         if (wmask[i]) begin
  //           mem[addr_i][i*DataBitsPerMask +: DataBitsPerMask] <=
  //             wdata_i[i*DataBitsPerMask +: DataBitsPerMask];
  //         end
  //       end
  //     end else begin
  //       rdata_o <= mem[addr_i];
  //     end
  //   end
  // end

// Conditional instantiation based on MaskWidth
generate
  if (MaskWidth == 1) begin : gen_array_1024x39
    sram_array_1p1024x39m39 sram_imem (
      .clk_i(clk_i),
      .req_i(req_i),
      .write_i(write_i),
      .addr_i(addr_i),
      .wdata_i(wdata_i),
      .wmask_i(wmask),
      .rdata_o(rdata_o)
    );
  end else begin : gen_array_128x312
    sram_array_1p128x312m39 sram_dmem (
      .clk_i(clk_i),
      .req_i(req_i),
      .write_i(write_i),
      .addr_i(addr_i),
      .wdata_i(wdata_i),
      .wmask_i(wmask),
      .rdata_o(rdata_o)
    );
  end
endgenerate

  `include "prim_util_memload.svh"
`endif
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_rom import prim_rom_pkg::*; #(
  parameter  int Width       = 32,
  parameter  int Depth       = 2048, // 8kB default
  parameter      MemInitFile = "", // VMEM file to initialize the memory with

  localparam int Aw          = $clog2(Depth)
) (
  input  logic             clk_i,
  input  logic             req_i,
  input  logic [Aw-1:0]    addr_i,
  output logic [Width-1:0] rdata_o,
  input rom_cfg_t          cfg_i
);

  logic unused_cfg;
  assign unused_cfg = ^cfg_i;

  logic [Width-1:0] mem [Depth];

  always_ff @(posedge clk_i) begin
    if (req_i) begin
      rdata_o <= mem[addr_i];
    end
  end

  `include "prim_util_memload.svh"

  ////////////////
  // ASSERTIONS //
  ////////////////

  // Control Signals should never be X
  `ASSERT(noXOnCsI, !$isunknown(req_i), clk_i, '0)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module implements different LFSR types:
//
// 0) Galois XOR type LFSR ([1], internal XOR gates, very fast).
//    Parameterizable width from 4 to 64 bits.
//    Coefficients obtained from [2].
//
// 1) Fibonacci XNOR type LFSR, parameterizable from 3 to 168 bits.
//    Coefficients obtained from [3].
//
// All flavors have an additional entropy input and lockup protection, which
// reseeds the state once it has accidentally fallen into the all-zero (XOR) or
// all-one (XNOR) state. Further, an external seed can be loaded into the LFSR
// state at runtime. If that seed is all-zero (XOR case) or all-one (XNOR case),
// the state will be reseeded in the next cycle using the lockup protection mechanism.
// Note that the external seed input takes precedence over internal state updates.
//
// All polynomials up to 34 bit in length have been verified in simulation.
//
// Refs: [1] https://en.wikipedia.org/wiki/Linear-feedback_shift_register
//       [2] https://users.ece.cmu.edu/~koopman/lfsr/
//       [3] https://www.xilinx.com/support/documentation/application_notes/xapp052.pdf

`include "prim_assert.sv"

module prim_lfsr #(
  // Lfsr Type, can be FIB_XNOR or GAL_XOR
  parameter                    LfsrType     = "GAL_XOR",
  // Lfsr width
  parameter int unsigned       LfsrDw       = 32,
  // Derived parameter, do not override
  localparam int unsigned      LfsrIdxDw    = $clog2(LfsrDw),
  // Width of the entropy input to be XOR'd into state (lfsr_q[EntropyDw-1:0])
  parameter int unsigned       EntropyDw    =  8,
  // Width of output tap (from lfsr_q[StateOutDw-1:0])
  parameter int unsigned       StateOutDw   =  8,
  // Lfsr reset state, must be nonzero!
  parameter logic [LfsrDw-1:0] DefaultSeed  = LfsrDw'(1),
  // Custom polynomial coeffs
  parameter logic [LfsrDw-1:0] CustomCoeffs = '0,
  // If StatePermEn is set to 1, the custom permutation specified via StatePerm is applied to the
  // state output, in order to break linear shifting patterns of the LFSR. Note that this
  // permutation represents a way of customizing the LFSR via a random netlist constant. This is
  // different from the NonLinearOut feature below which just transforms the output non-linearly
  // with a fixed function. In most cases, designers should consider enabling StatePermEn as it
  // comes basically "for free" in terms of area and timing impact. NonLinearOut on the other hand
  // has area and timing implications and designers should consider whether the use of that feature
  // is justified.
  parameter bit                StatePermEn  = 1'b0,
  parameter logic [LfsrDw-1:0][LfsrIdxDw-1:0] StatePerm = '0,
  // Enable this for DV, disable this for long LFSRs in FPV
  parameter bit                MaxLenSVA    = 1'b1,
  // Can be disabled in cases where seed and entropy
  // inputs are unused in order to not distort coverage
  // (the SVA will be unreachable in such cases)
  parameter bit                LockupSVA    = 1'b1,
  parameter bit                ExtSeedSVA   = 1'b1,
  // Introduce non-linearity to lfsr output. Note, unlike StatePermEn, this feature is not "for
  // free". Please double check that this feature is indeed required. Also note that this feature
  // is only available for LFSRs that have a power-of-two width greater or equal 16bit.
  parameter bit                NonLinearOut = 1'b0
) (
  input                         clk_i,
  input                         rst_ni,
  input                         seed_en_i, // load external seed into the state (takes precedence)
  input        [LfsrDw-1:0]     seed_i,    // external seed input
  input                         lfsr_en_i, // enables the LFSR
  input        [EntropyDw-1:0]  entropy_i, // additional entropy to be XOR'ed into the state
  output logic [StateOutDw-1:0] state_o    // (partial) LFSR state output
);

  // automatically generated with util/design/get-lfsr-coeffs.py script
  localparam int unsigned GAL_XOR_LUT_OFF = 4;
  localparam logic [63:0] GAL_XOR_COEFFS [61] =
    '{ 64'h9,
       64'h12,
       64'h21,
       64'h41,
       64'h8E,
       64'h108,
       64'h204,
       64'h402,
       64'h829,
       64'h100D,
       64'h2015,
       64'h4001,
       64'h8016,
       64'h10004,
       64'h20013,
       64'h40013,
       64'h80004,
       64'h100002,
       64'h200001,
       64'h400010,
       64'h80000D,
       64'h1000004,
       64'h2000023,
       64'h4000013,
       64'h8000004,
       64'h10000002,
       64'h20000029,
       64'h40000004,
       64'h80000057,
       64'h100000029,
       64'h200000073,
       64'h400000002,
       64'h80000003B,
       64'h100000001F,
       64'h2000000031,
       64'h4000000008,
       64'h800000001C,
       64'h10000000004,
       64'h2000000001F,
       64'h4000000002C,
       64'h80000000032,
       64'h10000000000D,
       64'h200000000097,
       64'h400000000010,
       64'h80000000005B,
       64'h1000000000038,
       64'h200000000000E,
       64'h4000000000025,
       64'h8000000000004,
       64'h10000000000023,
       64'h2000000000003E,
       64'h40000000000023,
       64'h8000000000004A,
       64'h100000000000016,
       64'h200000000000031,
       64'h40000000000003D,
       64'h800000000000001,
       64'h1000000000000013,
       64'h2000000000000034,
       64'h4000000000000001,
       64'h800000000000000D };

  // automatically generated with get-lfsr-coeffs.py script
  localparam int unsigned FIB_XNOR_LUT_OFF = 3;
  localparam logic [167:0] FIB_XNOR_COEFFS [166] =
    '{ 168'h6,
       168'hC,
       168'h14,
       168'h30,
       168'h60,
       168'hB8,
       168'h110,
       168'h240,
       168'h500,
       168'h829,
       168'h100D,
       168'h2015,
       168'h6000,
       168'hD008,
       168'h12000,
       168'h20400,
       168'h40023,
       168'h90000,
       168'h140000,
       168'h300000,
       168'h420000,
       168'hE10000,
       168'h1200000,
       168'h2000023,
       168'h4000013,
       168'h9000000,
       168'h14000000,
       168'h20000029,
       168'h48000000,
       168'h80200003,
       168'h100080000,
       168'h204000003,
       168'h500000000,
       168'h801000000,
       168'h100000001F,
       168'h2000000031,
       168'h4400000000,
       168'hA000140000,
       168'h12000000000,
       168'h300000C0000,
       168'h63000000000,
       168'hC0000030000,
       168'h1B0000000000,
       168'h300003000000,
       168'h420000000000,
       168'hC00000180000,
       168'h1008000000000,
       168'h3000000C00000,
       168'h6000C00000000,
       168'h9000000000000,
       168'h18003000000000,
       168'h30000000030000,
       168'h40000040000000,
       168'hC0000600000000,
       168'h102000000000000,
       168'h200004000000000,
       168'h600003000000000,
       168'hC00000000000000,
       168'h1800300000000000,
       168'h3000000000000030,
       168'h6000000000000000,
       168'hD800000000000000,
       168'h10000400000000000,
       168'h30180000000000000,
       168'h60300000000000000,
       168'h80400000000000000,
       168'h140000028000000000,
       168'h300060000000000000,
       168'h410000000000000000,
       168'h820000000001040000,
       168'h1000000800000000000,
       168'h3000600000000000000,
       168'h6018000000000000000,
       168'hC000000018000000000,
       168'h18000000600000000000,
       168'h30000600000000000000,
       168'h40200000000000000000,
       168'hC0000000060000000000,
       168'h110000000000000000000,
       168'h240000000480000000000,
       168'h600000000003000000000,
       168'h800400000000000000000,
       168'h1800000300000000000000,
       168'h3003000000000000000000,
       168'h4002000000000000000000,
       168'hC000000000000000018000,
       168'h10000000004000000000000,
       168'h30000C00000000000000000,
       168'h600000000000000000000C0,
       168'hC00C0000000000000000000,
       168'h140000000000000000000000,
       168'h200001000000000000000000,
       168'h400800000000000000000000,
       168'hA00000000001400000000000,
       168'h1040000000000000000000000,
       168'h2004000000000000000000000,
       168'h5000000000028000000000000,
       168'h8000000004000000000000000,
       168'h18600000000000000000000000,
       168'h30000000000000000C00000000,
       168'h40200000000000000000000000,
       168'hC0300000000000000000000000,
       168'h100010000000000000000000000,
       168'h200040000000000000000000000,
       168'h5000000000000000A0000000000,
       168'h800000010000000000000000000,
       168'h1860000000000000000000000000,
       168'h3003000000000000000000000000,
       168'h4010000000000000000000000000,
       168'hA000000000140000000000000000,
       168'h10080000000000000000000000000,
       168'h30000000000000000000180000000,
       168'h60018000000000000000000000000,
       168'hC0000000000000000300000000000,
       168'h140005000000000000000000000000,
       168'h200000001000000000000000000000,
       168'h404000000000000000000000000000,
       168'h810000000000000000000000000102,
       168'h1000040000000000000000000000000,
       168'h3000000000000006000000000000000,
       168'h5000000000000000000000000000000,
       168'h8000000004000000000000000000000,
       168'h18000000000000000000000000030000,
       168'h30000000030000000000000000000000,
       168'h60000000000000000000000000000000,
       168'hA0000014000000000000000000000000,
       168'h108000000000000000000000000000000,
       168'h240000000000000000000000000000000,
       168'h600000000000C00000000000000000000,
       168'h800000040000000000000000000000000,
       168'h1800000000000300000000000000000000,
       168'h2000000000000010000000000000000000,
       168'h4008000000000000000000000000000000,
       168'hC000000000000000000000000000000600,
       168'h10000080000000000000000000000000000,
       168'h30600000000000000000000000000000000,
       168'h4A400000000000000000000000000000000,
       168'h80000004000000000000000000000000000,
       168'h180000003000000000000000000000000000,
       168'h200001000000000000000000000000000000,
       168'h600006000000000000000000000000000000,
       168'hC00000000000000006000000000000000000,
       168'h1000000000000100000000000000000000000,
       168'h3000000000000006000000000000000000000,
       168'h6000000003000000000000000000000000000,
       168'h8000001000000000000000000000000000000,
       168'h1800000000000000000000000000C000000000,
       168'h20000000000001000000000000000000000000,
       168'h48000000000000000000000000000000000000,
       168'hC0000000000000006000000000000000000000,
       168'h180000000000000000000000000000000000000,
       168'h280000000000000000000000000000005000000,
       168'h60000000C000000000000000000000000000000,
       168'hC00000000000000000000000000018000000000,
       168'h1800000600000000000000000000000000000000,
       168'h3000000C00000000000000000000000000000000,
       168'h4000000080000000000000000000000000000000,
       168'hC000300000000000000000000000000000000000,
       168'h10000400000000000000000000000000000000000,
       168'h30000000000000000000006000000000000000000,
       168'h600000000000000C0000000000000000000000000,
       168'hC0060000000000000000000000000000000000000,
       168'h180000006000000000000000000000000000000000,
       168'h3000000000C0000000000000000000000000000000,
       168'h410000000000000000000000000000000000000000,
       168'hA00140000000000000000000000000000000000000 };

  logic lockup;
  logic [LfsrDw-1:0] lfsr_d, lfsr_q;
  logic [LfsrDw-1:0] next_lfsr_state, coeffs;

  // Enable the randomization of DefaultSeed using DefaultSeedLocal in DV simulations.
  `ifdef SIMULATION
  `ifdef VERILATOR
      localparam logic [LfsrDw-1:0] DefaultSeedLocal = DefaultSeed;

  `else
    logic [LfsrDw-1:0] DefaultSeedLocal;
    logic prim_lfsr_use_default_seed;

    initial begin : p_randomize_default_seed
      if (!$value$plusargs("prim_lfsr_use_default_seed=%0d", prim_lfsr_use_default_seed)) begin
        // 30% of the time, use the DefaultSeed parameter; 70% of the time, randomize it.
        `ASSERT_I(UseDefaultSeedRandomizeCheck_A, std::randomize(prim_lfsr_use_default_seed) with {
                                                  prim_lfsr_use_default_seed dist {0:/7, 1:/3};})
      end
      if (prim_lfsr_use_default_seed) begin
        DefaultSeedLocal = DefaultSeed;
      end else begin
        // Randomize the DefaultSeedLocal ensuring its not all 0s or all 1s.
        `ASSERT_I(DefaultSeedLocalRandomizeCheck_A, std::randomize(DefaultSeedLocal) with {
                                                    !(DefaultSeedLocal inside {'0, '1});})
      end
      $display("%m: DefaultSeed = 0x%0h, DefaultSeedLocal = 0x%0h", DefaultSeed, DefaultSeedLocal);
    end
  `endif  // ifdef VERILATOR

  `else
    localparam logic [LfsrDw-1:0] DefaultSeedLocal = DefaultSeed;

  `endif  // ifdef SIMULATION

  ////////////////
  // Galois XOR //
  ////////////////
  if (64'(LfsrType) == 64'("GAL_XOR")) begin : gen_gal_xor

    // if custom polynomial is provided
    if (CustomCoeffs > 0) begin : gen_custom
      assign coeffs = CustomCoeffs[LfsrDw-1:0];
    end else begin : gen_lut
      assign coeffs = GAL_XOR_COEFFS[LfsrDw-GAL_XOR_LUT_OFF][LfsrDw-1:0];
      // check that the most significant bit of polynomial is 1
      `ASSERT_INIT(MinLfsrWidth_A, LfsrDw >= $low(GAL_XOR_COEFFS)+GAL_XOR_LUT_OFF)
      `ASSERT_INIT(MaxLfsrWidth_A, LfsrDw <= $high(GAL_XOR_COEFFS)+GAL_XOR_LUT_OFF)
    end

    // calculate next state using internal XOR feedback and entropy input
    assign next_lfsr_state = LfsrDw'(entropy_i) ^ ({LfsrDw{lfsr_q[0]}} & coeffs) ^ (lfsr_q >> 1);

    // lockup condition is all-zero
    assign lockup = ~(|lfsr_q);

    // check that seed is not all-zero
    `ASSERT_INIT(DefaultSeedNzCheck_A, |DefaultSeedLocal)


  ////////////////////
  // Fibonacci XNOR //
  ////////////////////
  end else if (64'(LfsrType) == "FIB_XNOR") begin : gen_fib_xnor

    // if custom polynomial is provided
    if (CustomCoeffs > 0) begin : gen_custom
      assign coeffs = CustomCoeffs[LfsrDw-1:0];
    end else begin : gen_lut
      assign coeffs = FIB_XNOR_COEFFS[LfsrDw-FIB_XNOR_LUT_OFF][LfsrDw-1:0];
      // check that the most significant bit of polynomial is 1
      `ASSERT_INIT(MinLfsrWidth_A, LfsrDw >= $low(FIB_XNOR_COEFFS)+FIB_XNOR_LUT_OFF)
      `ASSERT_INIT(MaxLfsrWidth_A, LfsrDw <= $high(FIB_XNOR_COEFFS)+FIB_XNOR_LUT_OFF)
    end

    // calculate next state using external XNOR feedback and entropy input
    assign next_lfsr_state = LfsrDw'(entropy_i) ^ {lfsr_q[LfsrDw-2:0], ~(^(lfsr_q & coeffs))};

    // lockup condition is all-ones
    assign lockup = &lfsr_q;

    // check that seed is not all-ones
    `ASSERT_INIT(DefaultSeedNzCheck_A, !(&DefaultSeedLocal))


  /////////////
  // Unknown //
  /////////////
  end else begin : gen_unknown_type
    assign coeffs = '0;
    assign next_lfsr_state = '0;
    assign lockup = 1'b0;
    `ASSERT_INIT(UnknownLfsrType_A, 0)
  end


  //////////////////
  // Shared logic //
  //////////////////

  assign lfsr_d = (seed_en_i)           ? seed_i          :
                  (lfsr_en_i && lockup) ? DefaultSeedLocal     :
                  (lfsr_en_i)           ? next_lfsr_state :
                                          lfsr_q;

  logic [LfsrDw-1:0] sbox_out;
  if (NonLinearOut) begin : gen_out_non_linear
    // The "aligned" permutation ensures that adjacent bits do not go into the same SBox. It is
    // different from the state permutation that can be specified via the StatePerm parameter. The
    // permutation taps out 4 SBox input bits at regular stride intervals. E.g., for a 16bit
    // vector, the input assignment looks as follows:
    //
    // SBox0: 0,  4,  8, 12
    // SBox1: 1,  5,  9, 13
    // SBox2: 2,  6, 10, 14
    // SBox3: 3,  7, 11, 15
    //
    // Note that this permutation can be produced by filling the input vector into matrix columns
    // and reading out the SBox inputs as matrix rows.
    localparam int NumSboxes = LfsrDw / 4;
    // Fill in the input vector in col-major order.
    logic [3:0][NumSboxes-1:0][LfsrIdxDw-1:0] matrix_indices;
    for (genvar j = 0; j < LfsrDw; j++) begin : gen_input_idx_map
      assign matrix_indices[j / NumSboxes][j % NumSboxes] = j;
    end
    // Due to the LFSR shifting pattern, the above permutation has the property that the output of
    // SBox(n) is going to be equal to SBox(n+1) in the subsequent cycle (unless the LFSR polynomial
    // modifies some of the associated shifted bits via an XOR tap).
    // We therefore tweak this permutation by rotating and reversing some of the assignment matrix
    // columns. The rotation and reversion operations have been chosen such that this
    // generalizes to all power of two widths supported by the LFSR primitive. For 16bit, this
    // looks as follows:
    //
    // SBox0: 0,  6, 11, 14
    // SBox1: 1,  7, 10, 13
    // SBox2: 2,  4,  9, 12
    // SBox3: 3,  5,  8, 15
    //
    // This can be achieved by:
    //   1) down rotating the second column by NumSboxes/2
    //   2) reversing the third column
    //   3) down rotating the fourth column by 1 and reversing it
    //
    logic [3:0][NumSboxes-1:0][LfsrIdxDw-1:0] matrix_rotrev_indices;
    typedef logic [NumSboxes-1:0][LfsrIdxDw-1:0] matrix_col_t;

    // left-rotates a matrix column by the shift amount
    function automatic matrix_col_t lrotcol(matrix_col_t col, integer shift);
      matrix_col_t out;
      for (int k = 0; k < NumSboxes; k++) begin
        out[(k + shift) % NumSboxes] = col[k];
      end
      return out;
    endfunction : lrotcol

    // reverses a matrix column
    function automatic matrix_col_t revcol(logic [NumSboxes-1:0][LfsrIdxDw-1:0] col);
      return {<<LfsrIdxDw{col}};
    endfunction : revcol

    // Reverses a matrix column
    //zdr
    // function automatic matrix_col_t revcol(matrix_col_t col);
    //   matrix_col_t reversed_col;
    //   // Iterate over each row
    //   for (int row = 0; row < NumSboxes; row++) begin
    //     // Iterate over each bit within the row and reverse the bits
    //     for (int j = 0; j < LfsrIdxDw; j++) begin
    //       reversed_col[row][j] = col[row][LfsrIdxDw-1-j];
    //     end
    //   end
    //   return reversed_col;
    // endfunction : revcol

    always_comb begin : p_rotrev
      matrix_rotrev_indices[0] = matrix_indices[0];
      matrix_rotrev_indices[1] = lrotcol(matrix_indices[1], NumSboxes/2);
      matrix_rotrev_indices[2] = revcol(matrix_indices[2]);
      matrix_rotrev_indices[3] = revcol(lrotcol(matrix_indices[3], 1));
    end

    // Read out the matrix rows and linearize.
    logic [LfsrDw-1:0][LfsrIdxDw-1:0] sbox_in_indices;
    for (genvar k = 0; k < LfsrDw; k++) begin : gen_reverse_upper
      assign sbox_in_indices[k] = matrix_rotrev_indices[k % 4][k / 4];
    end

`ifndef SYNTHESIS
      // Check that the permutation is indeed a permutation.
      logic [LfsrDw-1:0] sbox_perm_test;
      always_comb begin : p_perm_check
        sbox_perm_test = '0;
        for (int k = 0; k < LfsrDw; k++) begin
          sbox_perm_test[sbox_in_indices[k]] = 1'b1;
        end
      end
      // All bit positions must be marked with 1.
      `ASSERT(SboxPermutationCheck_A, &sbox_perm_test)
`endif

`ifdef FPV_ON
      // Verify that the permutation indeed breaks linear shifting patterns of 4bit input groups.
      // The symbolic variables let the FPV tool select all sbox index combinations and linear shift
      // offsets.
      int shift;
      int unsigned sk, sj;
      `ASSUME(SjSkRange_M, (sj < NumSboxes) && (sk < NumSboxes))
      `ASSUME(SjSkDifferent_M, sj != sk)
      `ASSUME(SjSkStable_M, ##1 $stable(sj) && $stable(sk) && $stable(shift))
      `ASSERT(SboxInputIndexGroupIsUnique_A,
          !((((sbox_in_indices[sj * 4 + 0] + shift) % LfsrDw) == sbox_in_indices[sk * 4 + 0]) &&
            (((sbox_in_indices[sj * 4 + 1] + shift) % LfsrDw) == sbox_in_indices[sk * 4 + 1]) &&
            (((sbox_in_indices[sj * 4 + 2] + shift) % LfsrDw) == sbox_in_indices[sk * 4 + 2]) &&
            (((sbox_in_indices[sj * 4 + 3] + shift) % LfsrDw) == sbox_in_indices[sk * 4 + 3])))

      // this checks that the permutations does not preserve neighboring bit positions.
      // i.e. no two neighboring bits are mapped to neighboring bit positions.
      int y;
      int unsigned ik;
      `ASSUME(IkYRange_M, (ik < LfsrDw) && (y == 1 || y == -1))
      `ASSUME(IkStable_M, ##1 $stable(ik) && $stable(y))
      `ASSERT(IndicesNotAdjacent_A, (sbox_in_indices[ik] - sbox_in_indices[(ik + y) % LfsrDw]) != 1)
`endif

    // Use the permutation indices to create the SBox layer
    for (genvar k = 0; k < NumSboxes; k++) begin : gen_sboxes
      logic [3:0] sbox_in;
      assign sbox_in = {lfsr_q[sbox_in_indices[k*4 + 3]],
                        lfsr_q[sbox_in_indices[k*4 + 2]],
                        lfsr_q[sbox_in_indices[k*4 + 1]],
                        lfsr_q[sbox_in_indices[k*4 + 0]]};
      assign sbox_out[k*4 +: 4] = prim_cipher_pkg::PRINCE_SBOX4[sbox_in];
    end
  end else begin : gen_out_passthru
    assign sbox_out = lfsr_q;
  end

  // Random output permutation, defined at compile time
  if (StatePermEn) begin : gen_state_perm

    for (genvar k = 0; k < StateOutDw; k++) begin : gen_perm_loop
      assign state_o[k] = sbox_out[StatePerm[k]];
    end

    // if lfsr width is greater than the output, then by definition
    // not every bit will be picked
    if (LfsrDw > StateOutDw) begin : gen_tieoff_unused
      logic unused_sbox_out;
      assign unused_sbox_out = ^sbox_out;
    end

  end else begin : gen_no_state_perm
    assign state_o = StateOutDw'(sbox_out);
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_reg
    if (!rst_ni) begin
      lfsr_q <= DefaultSeedLocal;
    end else begin
      lfsr_q <= lfsr_d;
    end
  end


  ///////////////////////
  // shared assertions //
  ///////////////////////

  `ASSERT_KNOWN(DataKnownO_A, state_o)

// the code below is not meant to be synthesized,
// but it is intended to be used in simulation and FPV
`ifndef SYNTHESIS
  function automatic logic [LfsrDw-1:0] compute_next_state(logic [LfsrDw-1:0]    lfsrcoeffs,
                                                           logic [EntropyDw-1:0] entropy,
                                                           logic [LfsrDw-1:0]    current_state);
    logic state0;
    logic [LfsrDw-1:0] next_state;

    next_state = current_state;

    // Galois XOR
    if (64'(LfsrType) == 64'("GAL_XOR")) begin
      if (next_state == 0) begin
        next_state = DefaultSeedLocal;
      end else begin
        state0 = next_state[0];
        next_state = next_state >> 1;
        if (state0) next_state ^= lfsrcoeffs;
        next_state ^= LfsrDw'(entropy);
      end
    // Fibonacci XNOR
    end else if (64'(LfsrType) == "FIB_XNOR") begin
      if (&next_state) begin
        next_state = DefaultSeedLocal;
      end else begin
        state0 = ~(^(next_state & lfsrcoeffs));
        next_state = next_state << 1;
        next_state[0] = state0;
        next_state ^= LfsrDw'(entropy);
      end
    end else begin
      $error("unknown lfsr type");
    end

    return next_state;
  endfunction : compute_next_state

  // check whether next state is computed correctly
  // we shift the assertion by one clock cycle (##1) in order to avoid
  // erroneous SVA triggers right after reset deassertion in cases where
  // the precondition is true throughout the reset.
  // this can happen since the disable_iff evaluates using unsampled values,
  // meaning that the assertion may already read rst_ni == 1 on an active
  // clock edge while the flops in the design have not yet changed state.
  `ASSERT(NextStateCheck_A, ##1 lfsr_en_i && !seed_en_i |=> lfsr_q ==
      compute_next_state(coeffs, $past(entropy_i), $past(lfsr_q)))

  // Only check this if enabled.
  if (StatePermEn) begin : gen_perm_check
    // Check that the supplied permutation is valid.
    logic [LfsrDw-1:0] lfsr_perm_test;
    initial begin : p_perm_check
      lfsr_perm_test = '0;
      for (int k = 0; k < LfsrDw; k++) begin
        lfsr_perm_test[StatePerm[k]] = 1'b1;
      end
      // All bit positions must be marked with 1.
      `ASSERT_I(PermutationCheck_A, &lfsr_perm_test)
    end
  end

`endif

  `ASSERT_INIT(InputWidth_A, LfsrDw >= EntropyDw)
  `ASSERT_INIT(OutputWidth_A, LfsrDw >= StateOutDw)

  // MSB must be one in any case
  `ASSERT(CoeffCheck_A, coeffs[LfsrDw-1])

  // output check
  `ASSERT_KNOWN(OutputKnown_A, state_o)
  if (!StatePermEn && !NonLinearOut) begin : gen_output_sva
    `ASSERT(OutputCheck_A, state_o == StateOutDw'(lfsr_q))
  end
  // if no external input changes the lfsr state, a lockup must not occur (by design)
  //`ASSERT(NoLockups_A, (!entropy_i) && (!seed_en_i) |=> !lockup, clk_i, !rst_ni)
  `ASSERT(NoLockups_A, lfsr_en_i && !entropy_i && !seed_en_i |=> !lockup)

  // this can be disabled if unused in order to not distort coverage
  if (ExtSeedSVA) begin : gen_ext_seed_sva
    // check that external seed is correctly loaded into the state
    // rst_ni is used directly as part of the pre-condition since the usage of rst_ni
    // in disable_iff is unsampled.  See #1985 for more details
    `ASSERT(ExtDefaultSeedInputCheck_A, (seed_en_i && rst_ni) |=> lfsr_q == $past(seed_i))
  end

  // if the external seed mechanism is not used,
  // there is theoretically no way we end up in a lockup condition
  // in order to not distort coverage, this SVA can be disabled in such cases
  if (LockupSVA) begin : gen_lockup_mechanism_sva
    // check that a stuck LFSR is correctly reseeded
    `ASSERT(LfsrLockupCheck_A, lfsr_en_i && lockup && !seed_en_i |=> !lockup)
  end

  // If non-linear output requested, the LFSR width must be a power of 2 and greater than 16.
  if(NonLinearOut) begin : gen_nonlinear_align_check_sva
    `ASSERT_INIT(SboxByteAlign_A, 2**$clog2(LfsrDw) == LfsrDw && LfsrDw >= 16)
  end

  if (MaxLenSVA) begin : gen_max_len_sva
`ifndef SYNTHESIS
    // the code below is a workaround to enable long sequences to be checked.
    // some simulators do not support SVA sequences longer than 2**32-1.
    logic [LfsrDw-1:0] cnt_d, cnt_q;
    logic perturbed_d, perturbed_q;
    logic [LfsrDw-1:0] cmp_val;

    assign cmp_val = {{(LfsrDw-1){1'b1}}, 1'b0}; // 2**LfsrDw-2
    assign cnt_d = (lfsr_en_i && lockup)             ? '0           :
                   (lfsr_en_i && (cnt_q == cmp_val)) ? '0           :
                   (lfsr_en_i)                       ? cnt_q + 1'b1 :
                                                       cnt_q;

    assign perturbed_d = perturbed_q | (|entropy_i) | seed_en_i;

    always_ff @(posedge clk_i or negedge rst_ni) begin : p_max_len
      if (!rst_ni) begin
        cnt_q       <= '0;
        perturbed_q <= 1'b0;
      end else begin
        cnt_q       <= cnt_d;
        perturbed_q <= perturbed_d;
      end
    end

    `ASSERT(MaximalLengthCheck0_A, cnt_q == 0 |-> lfsr_q == DefaultSeedLocal,
        clk_i, !rst_ni || perturbed_q)
    `ASSERT(MaximalLengthCheck1_A, cnt_q != 0 |-> lfsr_q != DefaultSeedLocal,
        clk_i, !rst_ni || perturbed_q)
`endif
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// The module implements a binary tree to find the maximal entry. the solution
// has O(N) area and O(log(N)) delay complexity, and thus scales well with
// many input sources.
//
// Note that only input values marked as "valid" are respected in the maximum computation.
// If there are multiple valid inputs with the same value, the tree will always select the input
// with the smallest index.
//
// If none of the input values are valid, the output index will be 0 and the output value will
// be equal to the input value at index 0.


`include "prim_assert.sv"

module prim_max_tree #(
  parameter int NumSrc = 32,
  parameter int Width = 8,
  // Derived parameters
  localparam int SrcWidth = $clog2(NumSrc)
) (
  // The module is combinational - the clock and reset are only used for assertions.
  input                         clk_i,
  input                         rst_ni,
  input [NumSrc-1:0][Width-1:0] values_i,    // Input values
  input [NumSrc-1:0]            valid_i,     // Input valid bits
  output logic [Width-1:0]      max_value_o, // Maximum value
  output logic [SrcWidth-1:0]   max_idx_o,   // Index of the maximum value
  output logic                  max_valid_o  // Whether any of the inputs is valid
);

  ///////////////////////
  // Binary tree logic //
  ///////////////////////

  // This only works with 2 or more sources.
  `ASSERT_INIT(NumSources_A, NumSrc >= 2)

  // Align to powers of 2 for simplicity.
  // A full binary tree with N levels has 2**N + 2**N-1 nodes.
  localparam int NumLevels = $clog2(NumSrc);
  logic [2**(NumLevels+1)-2:0]               vld_tree;
  logic [2**(NumLevels+1)-2:0][SrcWidth-1:0] idx_tree;
  logic [2**(NumLevels+1)-2:0][Width-1:0]    max_tree;

  for (genvar level = 0; level < NumLevels+1; level++) begin : gen_tree
    //
    // level+1   C0   C1   <- "Base1" points to the first node on "level+1",
    //            \  /         these nodes are the children of the nodes one level below
    // level       Pa      <- "Base0", points to the first node on "level",
    //                         these nodes are the parents of the nodes one level above
    //
    // hence we have the following indices for the paPa, C0, C1 nodes:
    // Pa = 2**level     - 1 + offset       = Base0 + offset
    // C0 = 2**(level+1) - 1 + 2*offset     = Base1 + 2*offset
    // C1 = 2**(level+1) - 1 + 2*offset + 1 = Base1 + 2*offset + 1
    //
    localparam int Base0 = (2**level)-1;
    localparam int Base1 = (2**(level+1))-1;

    for (genvar offset = 0; offset < 2**level; offset++) begin : gen_level
      localparam int Pa = Base0 + offset;
      localparam int C0 = Base1 + 2*offset;
      localparam int C1 = Base1 + 2*offset + 1;

      // This assigns the input values, their corresponding IDs and valid signals to the tree leafs.
      if (level == NumLevels) begin : gen_leafs
        if (offset < NumSrc) begin : gen_assign
          assign vld_tree[Pa] = valid_i[offset];
          assign idx_tree[Pa] = offset;
          assign max_tree[Pa] = values_i[offset];
        end else begin : gen_tie_off
          assign vld_tree[Pa] = '0;
          assign idx_tree[Pa] = '0;
          assign max_tree[Pa] = '0;
        end
      // This creates the node assignments.
      end else begin : gen_nodes
        logic sel; // Local helper variable
        // In case only one of the parents is valid, forward that one
        // In case both parents are valid, forward the one with higher value
        assign sel = (~vld_tree[C0] & vld_tree[C1]) |
                     (vld_tree[C0] & vld_tree[C1] & logic'(max_tree[C1] > max_tree[C0]));
        // Forwarding muxes
        // Note: these ternaries have triggered a synthesis bug in Vivado versions older
        // than 2020.2. If the problem resurfaces again, have a look at issue #1408.
        assign vld_tree[Pa] = (sel) ? vld_tree[C1] : vld_tree[C0];
        assign idx_tree[Pa] = (sel) ? idx_tree[C1] : idx_tree[C0];
        assign max_tree[Pa] = (sel) ? max_tree[C1] : max_tree[C0];
      end
    end : gen_level
  end : gen_tree


  // The results can be found at the tree root
  assign max_valid_o = vld_tree[0];
  assign max_idx_o   = idx_tree[0];
  assign max_value_o = max_tree[0];

  ////////////////
  // Assertions //
  ////////////////

`ifdef INC_ASSERT
  //VCS coverage off
  // pragma coverage off

  // Helper functions for assertions below.
  function automatic logic [Width-1:0] max_value (input logic [NumSrc-1:0][Width-1:0] values_i,
                                                  input logic [NumSrc-1:0]            valid_i);
    logic [Width-1:0] value = '0;
    for (int k = 0; k < NumSrc; k++) begin
      if (valid_i[k] && values_i[k] > value) begin
        value = values_i[k];
      end
    end
    return value;
  endfunction : max_value

  function automatic logic [SrcWidth-1:0] max_idx (input logic [NumSrc-1:0][Width-1:0] values_i,
                                                   input logic [NumSrc-1:0]            valid_i);
    logic [Width-1:0] value = '0;
    logic [SrcWidth-1:0] idx = '0;
    for (int k = NumSrc-1; k >= 0; k--) begin
      if (valid_i[k] && values_i[k] >= value) begin
        value = values_i[k];
        idx = k;
      end
    end
    return idx;
  endfunction : max_idx

  logic [Width-1:0] max_value_exp;
  logic [SrcWidth-1:0] max_idx_exp;
  assign max_value_exp = max_value(values_i, valid_i);
  assign max_idx_exp = max_idx(values_i, valid_i);
  //VCS coverage on
  // pragma coverage on

  // TODO(10588): Below syntax is not supported in xcelium, track xcelium cases #46591452.
  // `ASSERT(ValidInImpliesValidOut_A, |valid_i <-> max_valid_o)
  `ASSERT(ValidInImpliesValidOut_A, |valid_i === max_valid_o)
  `ASSERT(MaxComputation_A, max_valid_o |-> max_value_o == max_value_exp)
  `ASSERT(MaxComputationInvalid_A, !max_valid_o |-> max_value_o == values_i[0])
  `ASSERT(MaxIndexComputation_A, max_valid_o |-> max_idx_o == max_idx_exp)
  `ASSERT(MaxIndexComputationInvalid_A, !max_valid_o |-> max_idx_o == '0)
`endif

endmodule : prim_max_tree


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Extend the output with the msb of the input

`include "prim_assert.sv"

module prim_msb_extend # (
  parameter int InWidth = 2,
  parameter int OutWidth = 2
) (
  input [InWidth-1:0] in_i,
  output [OutWidth-1:0] out_o
);

  `ASSERT_INIT(WidthCheck_A, OutWidth >= InWidth)

  localparam int WidthDiff = OutWidth - InWidth;

  if (WidthDiff == 0) begin : gen_feedthru
    assign out_o = in_i;
  end else begin : gen_tieoff
    assign out_o = {{WidthDiff{in_i[InWidth-1]}}, in_i};
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Domain-Oriented Masking GF(2) Multiplier with 2-shares
// ref: Higher-Order Side-Channel Protected Implementations of Keccak
//     https://eprint.iacr.org/2017/395.pdf
//
// q0 = a0 & b0 + (a0 & b1 + z)
// q1 = a1 & b1 + (a1 & b0 + z)
// () ==> registered
//
// all input should be stable for two clocks
// as the output is valid after a clock
// For z, it can use other slice from the state
// as it is fairly random w.r.t the current inputs.

// General formula of Q in the paper
// Qi = t{i,i} + Sig(j>i,d)(t{i,j}+Z{i+j*(j-1)/2}) + Sig(j<i,d)(t{i,j}+Z{j+i*(i-1)/2})
// for d=1 (NumShare 2 for first order protection)
// Q0 = t{0,0} + Sig(j>0,1)(t{0,j}+Z{j(j-1)/2}) + Sig(j<0,d)(..)
//    = a0&b0  + (a0&b1 + z0                    + 0)
// Q1 = t{1,1} + sig(j>1,1)(...) + sig(j<1,1)(t{1,j} + Z{j})
//    = a1&b1  + (0              + a1&b0 + z0)

`include "prim_assert.sv"

module prim_dom_and_2share #(
  parameter int DW = 64, // Input width
  parameter bit Pipeline = 1'b0 // Enable full pipelining
) (
  input clk_i,
  input rst_ni,

  input [DW-1:0] a0_i, // share0 of a
  input [DW-1:0] a1_i, // share1 of a
  input [DW-1:0] b0_i, // share0 of b
  input [DW-1:0] b1_i, // share1 of b
  input          z_valid_i, // random number input validity
  input [DW-1:0] z_i,  // random number

  output logic [DW-1:0] q0_o, // share0 of q
  output logic [DW-1:0] q1_o, // share1 of q
  output logic [DW-1:0] prd_o // pseudo-random data for other instances
);

  logic [DW-1:0] t0_d, t0_q, t1_d, t1_q;
  logic [DW-1:0] t_a0b0, t_a1b1;
  logic [DW-1:0] t_a0b0_d, t_a1b1_d;
  logic [DW-1:0] t_a0b1, t_a1b0;

  /////////////////
  // Calculation //
  /////////////////
  // Inner-domain terms
  assign t_a0b0_d = a0_i & b0_i;
  assign t_a1b1_d = a1_i & b1_i;

  // Cross-domain terms
  assign t_a0b1 = a0_i & b1_i;
  assign t_a1b0 = a1_i & b0_i;

  ///////////////
  // Resharing //
  ///////////////
  // Resharing of cross-domain terms

  // Preserve the logic sequence for XOR not to proceed cross-domain AND.
  prim_xor2 #(
    .Width ( DW*2 )
  ) u_prim_xor_t01 (
    .in0_i ( {t_a0b1, t_a1b0} ),
    .in1_i ( {z_i,    z_i}    ),
    .out_o ( {t0_d,   t1_d}   )
  );

  // Register stage
  prim_flop_en #(
    .Width      ( DW*2 ),
    .ResetValue ( '0   )
  ) u_prim_flop_t01 (
    .clk_i  ( clk_i        ),
    .rst_ni ( rst_ni       ),
    .en_i   ( z_valid_i    ),
    .d_i    ( {t0_d, t1_d} ),
    .q_o    ( {t0_q, t1_q} )
  );

  /////////////////////////
  // Optional Pipelining //
  /////////////////////////

  if (Pipeline == 1'b1) begin : gen_inner_domain_regs
    // Add pipeline registers on inner-domain terms prior to integration. This allows accepting new
    // input data every clock cycle and prevents SCA leakage occurring due to the integration of
    // reshared cross-domain terms with inner-domain terms derived from different input data.

    logic [DW-1:0] t_a0b0_q, t_a1b1_q;
    prim_flop_en #(
      .Width      ( DW*2 ),
      .ResetValue ( '0   )
    ) u_prim_flop_tab01 (
      .clk_i  ( clk_i                ),
      .rst_ni ( rst_ni               ),
      .en_i   ( z_valid_i            ),
      .d_i    ( {t_a0b0_d, t_a1b1_d} ),
      .q_o    ( {t_a0b0_q, t_a1b1_q} )
    );

    assign t_a0b0 = t_a0b0_q;
    assign t_a1b1 = t_a1b1_q;

  end else begin : gen_no_inner_domain_regs
    // Do not add the optional pipeline registers on the inner-domain terms. This allows to save
    // some area in case the multiplier does not need to accept new data in every cycle. However,
    // this can cause SCA leakage as during the clock cycle in which new data arrives, the new
    // inner-domain terms are integrated with the previous, reshared cross-domain terms.

    assign t_a0b0 = t_a0b0_d;
    assign t_a1b1 = t_a1b1_d;
  end

  /////////////////
  // Integration //
  /////////////////

  // Preserve the logic sequence for XOR not to proceed the inner-domain AND.
  prim_xor2 #(
    .Width ( DW*2 )
  ) u_prim_xor_q01 (
    .in0_i ( {t_a0b0, t_a1b1} ),
    .in1_i ( {t0_q,   t1_q}   ),
    .out_o ( {q0_o,   q1_o}   )
  );

  // Use intermediate results for remasking computations in another instance in the following
  // clock cycle. Use one share only. Directly use output of flops updating with z_valid_i.
  // t1_q is obtained by remasking t_a1b0 with z_i. Since z_i is uniformly distributed and
  // independent of a1/b0_i, t1_q is also uniformly distributed and independent of a1/b0_i.
  // For details, see Lemma 1 in Canright, "A very compact 'perfectly masked' S-box for AES
  // (corrected)" available at https://eprint.iacr.org/2009/011.pdf
  assign prd_o = t1_q;

  // DOM AND should be same as unmasked computation
  // The correct test sequence will be:
  //   1. inputs are changed
  //   2. check if z_valid_i,
  //   3. at the next cycle, inputs are still stable (assumption) - only in case Pipeline = 0
  //   4. and results Q == A & B (assertion)

  // To speed up the FPV process, random value is ready in less than or
  // equal to two cycles.
  `ASSUME_FPV(RandomReadyInShortTime_A,
    $changed(a0_i) || $changed(a1_i) || $changed(b0_i) || $changed(b1_i)
      |-> ##[0:2] z_valid_i,
    clk_i, !rst_ni)

  if (Pipeline == 0) begin: g_assert_stable
    // If Pipeline is not set, the computation takes two cycles without flop
    // crossing the domain. In this case, the signal should be stable for at
    // least two cycles.
    `ASSUME(StableTwoCycles_M,
      ($changed(a0_i)  || $changed(a1_i) || $changed(b0_i) || $changed(b1_i))
        ##[0:$] z_valid_i |=>
        $stable(a0_i) && $stable(a1_i) && $stable(b0_i) && $stable(b1_i))
  end

  `ASSERT(UnmaskedAndMatched_A,
    z_valid_i |=> (q0_o ^ q1_o) ==
      (($past(a0_i) ^ $past(a1_i)) & ($past(b0_i) ^ $past(b1_i))),
    clk_i, !rst_ni)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_sec_anchor_buf #(
  parameter int Width = 1
) (
  input        [Width-1:0] in_i,
  output logic [Width-1:0] out_o
);

  prim_buf #(
    .Width(Width)
  ) u_secure_anchor_buf (
    .in_i,
    .out_o
  );

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_sec_anchor_flop #(
  parameter int               Width      = 1,
  parameter logic [Width-1:0] ResetValue = 0
) (
  input                    clk_i,
  input                    rst_ni,
  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_o
);

  prim_flop #(
    .Width(Width),
    .ResetValue(ResetValue)
  ) u_secure_anchor_flop (
    .clk_i,
    .rst_ni,
    .d_i,
    .q_o
  );

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_sparse_fsm_flop #(
  parameter int               Width      = 1,
  parameter type              StateEnumT = logic [Width-1:0],
  parameter logic [Width-1:0] ResetValue = '0,
  // This should only be disabled in special circumstances, for example
  // in non-comportable IPs where an error does not trigger an alert.
  parameter bit               EnableAlertTriggerSVA = 1
`ifdef SIMULATION
  ,
  // In case this parameter is set to a non-empty string, the
  // prim_sparse_fsm_flop_if will also force the signal with this name
  // in the parent module that instantiates prim_sparse_fsm_flop.
  parameter string            CustomForceName = ""
`endif
) (
  input             clk_i,
  input             rst_ni,
  input  StateEnumT state_i,
  output StateEnumT state_o
);

  logic unused_err_o;

  logic [Width-1:0] state_raw;
  prim_flop #(
    .Width(Width),
    .ResetValue(ResetValue)
  ) u_state_flop (
    .clk_i,
    .rst_ni,
    .d_i(state_i),
    .q_o(state_raw)
  );
  assign state_o = StateEnumT'(state_raw);

  `ifdef INC_ASSERT
  assign unused_err_o = is_undefined_state(state_o);

  function automatic logic is_undefined_state(StateEnumT sig);
    // This is written with a vector in order to make it amenable to x-prop analysis.
    logic is_defined = 1'b0;
    for (int i = 0, StateEnumT t = t.first(); i < t.num(); i += 1, t = t.next()) begin
      is_defined |= (sig === t);
    end
    return ~is_defined;
  endfunction

  `else
    assign unused_err_o = 1'b0;
  `endif

  // If ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT is declared, the unused_assert_connected signal will
  // be set to 1 and the below check will pass.
  // If the assertion is not declared however, the statement below will fail.
  `ifdef INC_ASSERT
  logic unused_assert_connected;

  `ASSERT_INIT_NET(AssertConnected_A, unused_assert_connected === 1'b1 || !EnableAlertTriggerSVA)
  `endif

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package prim_subreg_pkg;

  // Register access specifier
  typedef enum logic [2:0] {
    SwAccessRW  = 3'd0, // Read-write
    SwAccessRO  = 3'd1, // Read-only
    SwAccessWO  = 3'd2, // Write-only
    SwAccessW1C = 3'd3, // Write 1 to clear
    SwAccessW1S = 3'd4, // Write 1 to set
    SwAccessW0C = 3'd5, // Write 0 to clear
    SwAccessRC  = 3'd6  // Read to clear. Do not use, only exists for compatibility.
  } sw_access_e;
endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Component handling register CDC
//
// Currently, this module only works correctly when paired with tlul_adapter_reg.
// This is because tlul_adapter_reg does not emit a new transaction to the same
// register if it discovers it is currently busy. Please see the BusySrcReqChk_A
// assertion below for more details.
//
// If in the future this assumption changes, we can modify this module easily to
// support the new behavior.

`include "prim_assert.sv"

module prim_reg_cdc #(
  parameter int DataWidth = 32,
  parameter logic [DataWidth-1:0] ResetVal = 32'h0,
  parameter logic [DataWidth-1:0] BitMask = 32'hFFFFFFFF,
  // whether this instance needs to support independent hardware writes
  parameter bit DstWrReq = 0
) (
  input clk_src_i,
  input rst_src_ni,
  input clk_dst_i,
  input rst_dst_ni,
  input src_regwen_i,
  input src_we_i,
  input src_re_i,
  input [DataWidth-1:0] src_wd_i,
  output logic src_busy_o,
  output logic [DataWidth-1:0] src_qs_o,
  input  [DataWidth-1:0] dst_ds_i,
  input  [DataWidth-1:0] dst_qs_i,
  input  dst_update_i,
  output logic dst_we_o,
  output logic dst_re_o,
  output logic dst_regwen_o,
  output logic [DataWidth-1:0] dst_wd_o
);

  ////////////////////////////
  // Source domain
  ////////////////////////////
  localparam int TxnWidth = 3;

  logic src_ack;
  logic src_busy_q;
  logic [DataWidth-1:0] src_q;
  logic [TxnWidth-1:0] txn_bits_q;
  logic src_req;

  assign src_req = src_we_i | src_re_i;

  // busy indication back-pressures upstream if the register is accessed
  // again.  The busy indication is also used as a "commit" indication for
  // resolving software and hardware write conflicts
  always_ff @(posedge clk_src_i or negedge rst_src_ni) begin
    if (!rst_src_ni) begin
      src_busy_q <= '0;
    end else if (src_req) begin
      src_busy_q <= 1'b1;
    end else if (src_ack) begin
      src_busy_q <= 1'b0;
    end
  end

  // A src_ack should only be sent if there was a src_req.
  // src_busy_q asserts whenever there is a src_req.  By association,
  // whenever src_ack is seen, then src_busy must be high.
  `ASSERT(SrcAckBusyChk_A, src_ack |-> src_busy_q, clk_src_i, !rst_src_ni)

  assign src_busy_o = src_busy_q;

  // src_q acts as both the write holding register and the software read back
  // register.
  // When software performs a write, the write data is captured in src_q for
  // CDC purposes.  When not performing a write, the src_q reflects the most recent
  // hardware value. For registes with no hardware access, this is simply the
  // the value programmed by software (or in the case R1C, W1C etc) the value after
  // the operation. For registers with hardware access, this reflects a potentially
  // delayed version of the real value, as the software facing updates lag real
  // time updates.
  //
  // To resolve software and hardware conflicts, the process is as follows:
  // When software issues a write, this module asserts "busy".  While busy,
  // src_q does not take on destination value updates.  Since the
  // logic has committed to updating based on software command, there is an irreversible
  // window from which hardware writes are ignored.  Once the busy window completes,
  // the cdc portion then begins sampling once more.
  //
  // This is consistent with prim_subreg_arb where during software / hardware conflicts,
  // software is always prioritized.  The main difference is the conflict resolution window
  // is now larger instead of just one destination clock cycle.

  logic busy;
  assign busy = src_busy_q & !src_ack;

  // This is the current destination value
  logic [DataWidth-1:0] dst_qs;
  logic src_update;
  always_ff @(posedge clk_src_i or negedge rst_src_ni) begin
    if (!rst_src_ni) begin
      src_q <= ResetVal;
      txn_bits_q <= '0;
    end else if (src_req) begin
      // See assertion below
      // At the beginning of a software initiated transaction, the following
      // values are captured in the src_q/txn_bits_q flops to ensure they cannot
      // change for the duration of the synchronization operation.
      src_q <= src_wd_i & BitMask;
      txn_bits_q <= {src_we_i, src_re_i, src_regwen_i};
    end else if (src_busy_q && src_ack || src_update && !busy) begin
      // sample data whenever a busy transaction finishes OR
      // when an update pulse is seen.
      // TODO: We should add a cover group to test different sync timings
      // between src_ack and src_update. Ie, there can be 3 scearios:
      // 1. update one cycle before ack
      // 2. ack one cycle before update
      // 3. update / ack on the same cycle
      // During all 3 cases the read data should be correct
      src_q <= dst_qs;
      txn_bits_q <= '0;
    end
  end

  // The current design (tlul_adapter_reg) does not spit out a request if the destination it chooses
  // (decoded from address) is busy. So this creates a situation in the current design where
  // src_req_i and busy can never be high at the same time.
  // While the code above could be coded directly to be expressed as `src_req & !busy`, which makes
  // the intent clearer, it ends up causing coverage holes from the tool's perspective since that
  // condition cannot be met.
  // Thus we add an assertion here to ensure the condition is always satisfied.
  `ASSERT(BusySrcReqChk_A, busy |-> !src_req, clk_src_i, !rst_src_ni)

  // reserved bits are not used
  logic unused_wd;
  assign unused_wd = ^src_wd_i;

  // src_q is always updated in the clk_src domain.
  // when performing an update to the destination domain, it is guaranteed
  // to not change by protocol.
  assign src_qs_o = src_q;
  assign dst_wd_o = src_q;

  ////////////////////////////
  // CDC handling
  ////////////////////////////

  logic dst_req_from_src;
  logic dst_req;


  // the software transaction is pulse synced across the domain.
  // the prim_reg_cdc_arb module handles conflicts with ongoing hardware updates.
  prim_pulse_sync u_src_to_dst_req (
    .clk_src_i,
    .rst_src_ni,
    .clk_dst_i,
    .rst_dst_ni,
    .src_pulse_i(src_req),
    .dst_pulse_o(dst_req_from_src)
  );

  prim_reg_cdc_arb #(
    .DataWidth(DataWidth),
    .ResetVal(ResetVal),
    .DstWrReq(DstWrReq)
  ) u_arb (
    .clk_src_i,
    .rst_src_ni,
    .clk_dst_i,
    .rst_dst_ni,
    .src_ack_o(src_ack),
    .src_update_o(src_update),
    .dst_req_i(dst_req_from_src),
    .dst_req_o(dst_req),
    .dst_update_i,
    .dst_ds_i,
    .dst_qs_i,
    .dst_qs_o(dst_qs)
  );


  // Each is valid only when destination request pulse is high
  assign {dst_we_o, dst_re_o, dst_regwen_o} = txn_bits_q & {TxnWidth{dst_req}};

  `ASSERT_KNOWN(SrcBusyKnown_A, src_busy_o, clk_src_i, !rst_src_ni)
  `ASSERT_KNOWN(DstReqKnown_A, dst_req, clk_dst_i, !rst_dst_ni)

  // If busy goes high, we must eventually see an ack
  `ifdef FPV_ON
    `ASSERT(HungHandShake_A, $rose(src_req) |-> strong(##[0:$] src_ack), clk_src_i, !rst_src_ni)
    // TODO: #14913 check if we can add additional sim assertions.
  `endif
endmodule // prim_subreg_cdc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Component handling register CDC

`include "prim_assert.sv"

// There are three handling scenarios.
// 1. The register can only be updated by software.
// 2. The register can be updated by both software and hardware.
// 3. The register can only be updated by hardware.
//
// For the first scenario, hardware updates are completely ignored.
// The software facing register (`src_q` in prim_reg_cdc) simply reflects
// the value affected by software.  Since there is no possibility the
// register value can change otherwise, there is no need to sample or
// do any other coordination between the two domains. In this case,
// we use the gen_passthru block below.
//
// For the second scenario, one of 4 things can happen:
// 1. A software update without conflict
// 2. A hardware update without conflict
// 3. A software update is initiated when a hardware update is in-flight
// 4. A hardware update is initiated when a software update is in-flight
//
// For the first case, it behaves similarly to the gen_passthru scenario.
//
// For the second case, the hardware update indication and update value are
// captured, and the intent to change is synchronized back to the software
// domain. While this happens, other hardware updates are ignored. Any hardware
// change during the update is then detected as a difference between the
// transit register `dst_qs_o` and the current hardware register value `dst_qs_i`.
// When this change is observed after the current handshake completes, another
// handshake event is generated to bring the latest hardware value over to the
// software domain.
//
// For the third case, if a hardware update event is already in progress, the
// software event is held and not acknowledged.  Once the hardware event completes,
// then the software event proceeds through its normal updating process.
//
// For the forth case, if a hardware update event is received while a software
// update is in progress, the hardware update is ignored, and the logic behaves
// similarly to the second case. Specifically, after the software update completes,
// a delta is observed between the transit register and the current hardware value,
// and a new handshake event is generated.
//
// The third scenario can be folded into the second scenario. The only difference
// is that of the 4 cases identified, only case 2 can happen since there is never a
// software initiated update.

module prim_reg_cdc_arb #(
  parameter int DataWidth = 32,
  parameter logic [DataWidth-1:0] ResetVal = 32'h0,
  parameter bit DstWrReq = 0
) (
  input clk_src_i,
  input rst_src_ni,
  input clk_dst_i,
  input rst_dst_ni,
  // destination side acknowledging a software transaction
  output logic src_ack_o,
  // destination side requesting a source side update after
  // after hw update
  output logic src_update_o,
  // input request from prim_reg_cdc
  input dst_req_i,
  // output request to prim_subreg
  output logic dst_req_o,
  input dst_update_i,
  // ds allows us to sample the destination domain register
  // one cycle earlier instead of waiting for it to be reflected
  // in the qs.
  // This is important because a general use case is that interrupts
  // are captured alongside payloads from the destination domain into
  // the source domain. If we rely on `qs` only, then it is very likely
  // that the software observed value will be behind the interrupt
  // assertion.  If the destination clock is very slow, this can seem
  // an error on the part of the hardware.
  input [DataWidth-1:0] dst_ds_i,
  input [DataWidth-1:0] dst_qs_i,
  output logic [DataWidth-1:0] dst_qs_o
);

  typedef enum logic {
    SelSwReq,
    SelHwReq
  } req_sel_e;

  typedef enum logic [1:0] {
    StIdle,
    StWait
  } state_e;


  // Only honor the incoming destinate update request if the incoming
  // value is actually different from what is already completed in the
  // handshake
  logic dst_update;
  assign dst_update = dst_update_i & (dst_qs_o != dst_ds_i);

  if (DstWrReq) begin : gen_wr_req
    logic dst_lat_q;
    logic dst_lat_d;
    logic dst_update_req;
    logic dst_update_ack;
    req_sel_e id_q;

    state_e state_q, state_d;
    // Make sure to indent the following later
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        state_q <= StIdle;
      end else begin
        state_q <= state_d;
      end
    end

    logic busy;
    logic dst_req_q, dst_req;
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        dst_req_q <= '0;
      end else if (dst_req_q && dst_lat_d) begin
        // if request is held, when the transaction starts,
        // automatically clear.
        // dst_lat_d is safe to used here because dst_req_q, if set,
        // always has priority over other hardware based events.
        dst_req_q <= '0;
      end else if (dst_req_i && !dst_req_q && busy) begin
        // if destination request arrives when a handshake event
        // is already ongoing, hold on to request and send later
        dst_req_q <= 1'b1;
      end
    end
    assign dst_req = dst_req_q | dst_req_i;

    // Hold data at the beginning of a transaction
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        dst_qs_o <= ResetVal;
      end else if (dst_lat_d) begin
        dst_qs_o <= dst_ds_i;
      end else if (dst_lat_q) begin
        dst_qs_o <= dst_qs_i;
      end
    end

    // Which type of transaction is being ack'd back?
    // 0 - software initiated request
    // 1 - hardware initiated request
    // The id information is used by prim_reg_cdc to disambiguate
    // simultaneous updates from software and hardware.
    // See scenario 2 case 3 for an example of how this is handled.
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        id_q <= SelSwReq;
      end else if (dst_update_req && dst_update_ack) begin
        id_q <= SelSwReq;
      end else if (dst_req && dst_lat_d) begin
        id_q <= SelSwReq;
      end else if (!dst_req && dst_lat_d) begin
        id_q <= SelHwReq;
      end else if (dst_lat_q) begin
        id_q <= SelHwReq;
      end
    end

    // if a destination update is received when the system is idle and there is no
    // software side request, hw update must be selected.
    `ASSERT(DstUpdateReqCheck_A, ##1 dst_update & !dst_req & !busy |=> id_q == SelHwReq,
      clk_dst_i, !rst_dst_ni)

    // if hw select was chosen, then it must be the case there was a destination update
    // indication or there was a difference between the transit register and the
    // latest incoming value.
    `ASSERT(HwIdSelCheck_A, $rose(id_q == SelHwReq) |-> $past(dst_update_i, 1) ||
      $past(dst_lat_q, 1),
      clk_dst_i, !rst_dst_ni)


    // send out prim_subreg request only when proceeding
    // with software request
    assign dst_req_o = ~busy & dst_req;

    logic dst_hold_req;
    always_comb begin
      state_d = state_q;
      dst_hold_req = '0;

      // depending on when the request is received, we
      // may latch d or q.
      dst_lat_q = '0;
      dst_lat_d = '0;

      busy = 1'b1;

      unique case (state_q)
        StIdle: begin
          busy = '0;
          if (dst_req) begin
            // there's a software issued request for change
            state_d = StWait;
            dst_lat_d = 1'b1;
          end else if (dst_update) begin
            state_d = StWait;
            dst_lat_d = 1'b1;
          end else if (dst_qs_o != dst_qs_i) begin
            // there's a direct destination update
            // that was blocked by an ongoing transaction
            state_d = StWait;
            dst_lat_q = 1'b1;
          end
        end

        StWait: begin
          dst_hold_req = 1'b1;
          if (dst_update_ack) begin
            state_d = StIdle;
          end
        end

        default: begin
          state_d = StIdle;
        end
      endcase // unique case (state_q)
    end // always_comb

    assign dst_update_req = dst_hold_req | dst_lat_d | dst_lat_q;
    logic src_req;
    prim_sync_reqack u_dst_update_sync (
      .clk_src_i(clk_dst_i),
      .rst_src_ni(rst_dst_ni),
      .clk_dst_i(clk_src_i),
      .rst_dst_ni(rst_src_ni),
      .req_chk_i(1'b1),
      .src_req_i(dst_update_req),
      .src_ack_o(dst_update_ack),
      .dst_req_o(src_req),
      // immediate ack
      .dst_ack_i(src_req)
    );

    assign src_ack_o = src_req & (id_q == SelSwReq);
    assign src_update_o = src_req & (id_q == SelHwReq);

    // once hardware makes an update request, we must eventually see an update pulse
    `ifdef FPV_ON
      `ASSERT(ReqTimeout_A, $rose(id_q == SelHwReq) |-> s_eventually(src_update_o),
              clk_src_i, !rst_src_ni)
      // TODO: #14913 check if we can add additional sim assertions.
    `endif

    `ifdef FPV_ON
      //VCS coverage off
      // pragma coverage off

      logic async_flag;
      always_ff @(posedge clk_dst_i or negedge rst_dst_ni or posedge src_update_o) begin
        if (!rst_dst_ni) begin
          async_flag <= '0;
        end else if (src_update_o) begin
          async_flag <= '0;
        end else if (dst_update && !dst_req_o && !busy) begin
          async_flag <= 1'b1;
        end
      end

      //VCS coverage on
      // pragma coverage on

      // once hardware makes an update request, we must eventually see an update pulse
      // TODO: #14913 check if we can add additional sim assertions.
      `ASSERT(UpdateTimeout_A, $rose(async_flag) |-> s_eventually(src_update_o),
              clk_src_i, !rst_src_ni)
    `endif

  end else begin : gen_passthru
    // when there is no possibility of conflicting HW transactions,
    // we can assume that dst_qs_i will only ever take on the value
    // that is directly related to the transaction. As a result,
    // there is no need to latch further, and the end destination
    // can in fact be used as the holding register.
    assign dst_qs_o = dst_qs_i;
    assign dst_req_o = dst_req_i;

    // since there are no hw transactions, src_update_o is always '0
    assign src_update_o = '0;

    prim_pulse_sync u_dst_to_src_ack (
      .clk_src_i(clk_dst_i),
      .rst_src_ni(rst_dst_ni),
      .clk_dst_i(clk_src_i),
      .rst_dst_ni(rst_src_ni),
      .src_pulse_i(dst_req_i),
      .dst_pulse_o(src_ack_o)
    );

    logic unused_sigs;
    assign unused_sigs = |{dst_ds_i, dst_update};
  end



endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register slice conforming to Comportibility guide.

module prim_subreg
  import prim_subreg_pkg::*;
#(
  parameter int            DW       = 32,
  parameter sw_access_e    SwAccess = SwAccessRW,
  parameter logic [DW-1:0] RESVAL   = '0    // reset value
) (
  input clk_i,
  input rst_ni,

  // From SW: valid for RW, WO, W1C, W1S, W0C, RC
  // In case of RC, Top connects Read Pulse to we
  input          we,
  input [DW-1:0] wd,

  // From HW: valid for HRW, HWO
  input          de,
  input [DW-1:0] d,

  // output to HW and Reg Read
  output logic          qe,
  output logic [DW-1:0] q,

  // ds and qs have slightly different timing.
  // ds is the data that will be written into the flop,
  // while qs is the current flop value exposed to software.
  output logic [DW-1:0] ds,
  output logic [DW-1:0] qs
);

  logic          wr_en;
  logic [DW-1:0] wr_data;

  prim_subreg_arb #(
    .DW       ( DW       ),
    .SwAccess ( SwAccess )
  ) wr_en_data_arb (
    .we,
    .wd,
    .de,
    .d,
    .q,
    .wr_en,
    .wr_data
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      q <= RESVAL;
    end else if (wr_en) begin
      q <= wr_data;
    end
  end

  // feed back out for consolidation
  assign ds = wr_en ? wr_data : qs;
  assign qe = wr_en;
  assign qs = q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Write enable and data arbitration logic for register slice conforming to Comportibility guide.

module prim_subreg_arb
  import prim_subreg_pkg::*;
#(
  parameter int         DW       = 32,
  parameter sw_access_e SwAccess = SwAccessRW
) (
  // From SW: valid for RW, WO, W1C, W1S, W0C, RC.
  // In case of RC, top connects read pulse to we.
  input          we,
  input [DW-1:0] wd,

  // From HW: valid for HRW, HWO.
  input          de,
  input [DW-1:0] d,

  // From register: actual reg value.
  input [DW-1:0] q,

  // To register: actual write enable and write data.
  output logic          wr_en,
  output logic [DW-1:0] wr_data
);

  if (SwAccess inside {SwAccessRW, SwAccessWO}) begin : gen_w
    assign wr_en   = we | de;
    assign wr_data = (we == 1'b1) ? wd : d; // SW higher priority
    // Unused q - Prevent lint errors.
    logic [DW-1:0] unused_q;
    assign unused_q = q;
  end else if (SwAccess == SwAccessRO) begin : gen_ro
    assign wr_en   = de;
    assign wr_data = d;
    // Unused we, wd, q - Prevent lint errors.
    logic          unused_we;
    logic [DW-1:0] unused_wd;
    logic [DW-1:0] unused_q;
    assign unused_we = we;
    assign unused_wd = wd;
    assign unused_q  = q;
  end else if (SwAccess == SwAccessW1S) begin : gen_w1s
    // If SwAccess is W1S, then assume hw tries to clear.
    // So, give a chance HW to clear when SW tries to set.
    // If both try to set/clr at the same bit pos, SW wins.
    assign wr_en   = we | de;
    assign wr_data = (de ? d : q) | (we ? wd : '0);
  end else if (SwAccess == SwAccessW1C) begin : gen_w1c
    // If SwAccess is W1C, then assume hw tries to set.
    // So, give a chance HW to set when SW tries to clear.
    // If both try to set/clr at the same bit pos, SW wins.
    assign wr_en   = we | de;
    assign wr_data = (de ? d : q) & (we ? ~wd : '1);
  end else if (SwAccess == SwAccessW0C) begin : gen_w0c
    assign wr_en   = we | de;
    assign wr_data = (de ? d : q) & (we ? wd : '1);
  end else if (SwAccess == SwAccessRC) begin : gen_rc
    // This swtype is not recommended but exists for compatibility.
    // WARN: we signal is actually read signal not write enable.
    assign wr_en  = we | de;
    assign wr_data = (de ? d : q) & (we ? '0 : '1);
    // Unused wd - Prevent lint errors.
    logic [DW-1:0] unused_wd;
    assign unused_wd = wd;
  end else begin : gen_hw
    assign wr_en   = de;
    assign wr_data = d;
    // Unused we, wd, q - Prevent lint errors.
    logic          unused_we;
    logic [DW-1:0] unused_wd;
    logic [DW-1:0] unused_q;
    assign unused_we = we;
    assign unused_wd = wd;
    assign unused_q  = q;
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register slice conforming to Comportibility guide.

module prim_subreg_ext #(
  parameter int unsigned DW = 32
) (
  input          re,
  input          we,
  input [DW-1:0] wd,

  input [DW-1:0] d,

  // output to HW and Reg Read
  output logic          qe,
  output logic          qre,
  output logic [DW-1:0] q,
  output logic [DW-1:0] ds,
  output logic [DW-1:0] qs
);

  // for external registers, there is no difference
  // between qs and ds
  assign ds = d;
  assign qs = d;
  assign q = wd;
  assign qe = we;
  assign qre = re;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Shadowed register slice conforming to Comportibility guide.

`include "prim_assert.sv"

module prim_subreg_shadow
  import prim_subreg_pkg::*;
#(
  parameter int            DW       = 32,
  parameter sw_access_e    SwAccess = SwAccessRW,
  parameter logic [DW-1:0] RESVAL   = '0    // reset value
) (
  input clk_i,
  input rst_ni,
  input rst_shadowed_ni,

  // From SW: valid for RW, WO, W1C, W1S, W0C, RC.
  // SW reads clear phase unless SwAccess is RO.
  input          re,
  // In case of RC, top connects read pulse to we.
  input          we,
  input [DW-1:0] wd,

  // From HW: valid for HRW, HWO.
  input          de,
  input [DW-1:0] d,

  // Output to HW and Reg Read
  output logic          qe,
  output logic [DW-1:0] q,
  output logic [DW-1:0] ds,
  output logic [DW-1:0] qs,

  // Phase output to HW
  output logic phase,

  // Error conditions
  output logic err_update,
  output logic err_storage
);

  // Since the shadow register works with the 1's complement value,
  // we need to invert the polarity of the SW access if it is either "W1S" or "W0C".
  // W1C is forbidden since the W0S complement is not implemented.
  `ASSERT_INIT(CheckSwAccessIsLegal_A,
      SwAccess inside {SwAccessRW, SwAccessRO, SwAccessWO, SwAccessW1S, SwAccessW0C})
  localparam sw_access_e InvertedSwAccess = (SwAccess == SwAccessW1S) ? SwAccessW0C :
                                            (SwAccess == SwAccessW0C) ? SwAccessW1S : SwAccess;

  // For the staging register, we set the SwAccess to RW in case of W1S and W0C in
  // order to always capture the data value on the first write operation - no matter
  // whether the data value will actually have an effect. That way, we can still capture
  // inconsistent double writes which would otherwise be ignored due to the data value filtering
  // effect that W1S and W0C can have.
  localparam sw_access_e StagedSwAccess = (SwAccess == SwAccessW1S) ? SwAccessRW :
                                          (SwAccess == SwAccessW0C) ? SwAccessRW : SwAccess;

  // Subreg control signals
  logic          phase_clear;
  logic          phase_q;
  logic          staged_we, shadow_we, committed_we;
  logic          staged_de, shadow_de, committed_de;

  // Subreg status and data signals
  logic          committed_qe;
  logic [DW-1:0] staged_q,  shadow_q,  committed_q;
  logic [DW-1:0] committed_qs;

  // Effective write enable and write data signals.
  // These depend on we, de and wd, d, q as well as SwAccess.
  logic          wr_en;
  logic [DW-1:0] wr_data;

  prim_subreg_arb #(
    .DW       ( DW       ),
    .SwAccess ( SwAccess )
  ) wr_en_data_arb (
    .we      ( we      ),
    .wd      ( wd      ),
    .de      ( de      ),
    .d       ( d       ),
    .q       ( q       ),
    .wr_en   ( wr_en   ),
    .wr_data ( wr_data )
  );

  // Phase clearing:
  // - SW reads clear phase unless SwAccess is RO.
  // - In case of RO, SW should not interfere with update process.
  assign phase_clear = (SwAccess == SwAccessRO) ? 1'b0 : re;

  // Phase tracker:
  // - Reads from SW clear the phase back to 0.
  // - Writes have priority (can come from SW or HW).
  always_ff @(posedge clk_i or negedge rst_ni) begin : phase_reg
    if (!rst_ni) begin
      phase_q <= 1'b0;
    end else if (wr_en && !err_storage) begin
      phase_q <= ~phase_q;
    end else if (phase_clear || err_storage) begin
      phase_q <= 1'b0;
    end
  end

  // The staged register:
  // - Holds the 1's complement value.
  // - Written in Phase 0.
  // - Once storage error occurs, do not allow any further update until reset
  assign staged_we = we & ~phase_q & ~err_storage;
  assign staged_de = de & ~phase_q & ~err_storage;
  prim_subreg #(
    .DW       ( DW             ),
    .SwAccess ( StagedSwAccess ),
    .RESVAL   ( ~RESVAL        )
  ) staged_reg (
    .clk_i    ( clk_i     ),
    .rst_ni   ( rst_ni    ),
    .we       ( staged_we ),
    .wd       ( ~wr_data  ),
    .de       ( staged_de ),
    .d        ( ~d        ),
    .qe       (           ),
    .q        ( staged_q  ),
    .ds       (           ),
    .qs       (           )
  );

  // The shadow register:
  // - Holds the 1's complement value.
  // - Written in Phase 1.
  // - Writes are ignored in case of update errors.
  // - Gets the value from the staged register.
  // - Once storage error occurs, do not allow any further update until reset
  assign shadow_we = we & phase_q & ~err_update & ~err_storage;
  assign shadow_de = de & phase_q & ~err_update & ~err_storage;
  prim_subreg #(
    .DW       ( DW               ),
    .SwAccess ( InvertedSwAccess ),
    .RESVAL   ( ~RESVAL          )
  ) shadow_reg (
    .clk_i    ( clk_i           ),
    .rst_ni   ( rst_shadowed_ni ),
    .we       ( shadow_we       ),
    .wd       ( staged_q        ),
    .de       ( shadow_de       ),
    .d        ( staged_q        ),
    .qe       (                 ),
    .q        ( shadow_q        ),
    .ds       (                 ),
    .qs       (                 )
  );

  // The committed register:
  // - Written in Phase 1.
  // - Writes are ignored in case of update errors.
  assign committed_we = shadow_we;
  assign committed_de = shadow_de;
  prim_subreg #(
    .DW       ( DW       ),
    .SwAccess ( SwAccess ),
    .RESVAL   ( RESVAL   )
  ) committed_reg (
    .clk_i    ( clk_i        ),
    .rst_ni   ( rst_ni       ),
    .we       ( committed_we ),
    .wd       ( wr_data      ),
    .de       ( committed_de ),
    .d        ( d            ),
    .qe       ( committed_qe ),
    .q        ( committed_q  ),
    .ds       ( ds           ),
    .qs       ( committed_qs )
  );

  // Output phase for hwext.
  assign phase = phase_q;

  // Error detection - all bits must match.
  assign err_update  = (~staged_q != wr_data) ? phase_q & wr_en : 1'b0;
  assign err_storage = (~shadow_q != committed_q);

  // Remaining output assignments
  assign qe = committed_qe;
  assign q  = committed_q;
  assign qs = committed_qs;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Based on prim_max_tree, this module implements an explicit binary tree to find the
// sum of this inputs. The solution has O(N) area and O(log(N)) delay complexity, and
// thus scales well with many input sources.
//
// Note that only input values marked as "valid" are respected in the maximum computation.
// Invalid values are treated as 0.
//

`include "prim_assert.sv"

module prim_sum_tree #(
  parameter int NumSrc = 32,
  parameter int Width = 8
) (
  // The module is combinational - the clock and reset are only used for assertions.
  input                         clk_i,
  input                         rst_ni,
  input [NumSrc-1:0][Width-1:0] values_i,    // Input values
  input [NumSrc-1:0]            valid_i,     // Input valid bits
  output logic [Width-1:0]      sum_value_o, // Summation result
  output logic                  sum_valid_o  // Whether any of the inputs is valid
);

  ///////////////////////
  // Binary tree logic //
  ///////////////////////

  // This only works with 2 or more sources.
  `ASSERT_INIT(NumSources_A, NumSrc >= 2)

  // Align to powers of 2 for simplicity.
  // A full binary tree with N levels has 2**N + 2**N-1 nodes.
  localparam int NumLevels = $clog2(NumSrc);
  logic [2**(NumLevels+1)-2:0]               vld_tree;
  logic [2**(NumLevels+1)-2:0][Width-1:0]    sum_tree;

  for (genvar level = 0; level < NumLevels+1; level++) begin : gen_tree
    //
    // level+1   C0   C1   <- "Base1" points to the first node on "level+1",
    //            \  /         these nodes are the children of the nodes one level below
    // level       Pa      <- "Base0", points to the first node on "level",
    //                         these nodes are the parents of the nodes one level above
    //
    // hence we have the following indices for the paPa, C0, C1 nodes:
    // Pa = 2**level     - 1 + offset       = Base0 + offset
    // C0 = 2**(level+1) - 1 + 2*offset     = Base1 + 2*offset
    // C1 = 2**(level+1) - 1 + 2*offset + 1 = Base1 + 2*offset + 1
    //
    localparam int Base0 = (2**level)-1;
    localparam int Base1 = (2**(level+1))-1;

    for (genvar offset = 0; offset < 2**level; offset++) begin : gen_level
      localparam int Pa = Base0 + offset;
      localparam int C0 = Base1 + 2*offset;
      localparam int C1 = Base1 + 2*offset + 1;

      // This assigns the input values, their corresponding IDs and valid signals to the tree leafs.
      if (level == NumLevels) begin : gen_leafs
        if (offset < NumSrc) begin : gen_assign
          assign vld_tree[Pa] = valid_i[offset];
          assign sum_tree[Pa] = values_i[offset];
        end else begin : gen_tie_off
          assign vld_tree[Pa] = '0;
          assign sum_tree[Pa] = '0;
        end
      // This creates the node assignments.
      end else begin : gen_nodes
        logic [Width-1:0] node_sum; // Local helper variable
        // In case only one of the parents is valid, forward that one
        // In case both parents are valid, forward the one with higher value
        assign node_sum = (vld_tree[C0] & vld_tree[C1]) ? sum_tree[C1] + sum_tree[C0] :
                          (vld_tree[C0])                ? sum_tree[C0] :
                          (vld_tree[C1])                ? sum_tree[C1] :
                          {Width'(0)};

        // Forwarding muxes
        // Note: these ternaries have triggered a synthesis bug in Vivado versions older
        // than 2020.2. If the problem resurfaces again, have a look at issue #1408.
        assign vld_tree[Pa] = vld_tree[C1] | vld_tree[C0];
        assign sum_tree[Pa] = node_sum;
      end
    end : gen_level
  end : gen_tree


  // The results can be found at the tree root
  assign sum_valid_o = vld_tree[0];
  assign sum_value_o = sum_tree[0];

  ////////////////
  // Assertions //
  ////////////////

`ifdef INC_ASSERT
  //VCS coverage off
  // pragma coverage off

  // Helper functions for assertions below.
  function automatic logic [Width-1:0] sum_value (input logic [NumSrc-1:0][Width-1:0] values_i,
                                                  input logic [NumSrc-1:0]            valid_i);
    logic [Width-1:0] sum = '0;
    for (int k = 0; k < NumSrc; k++) begin
      if (valid_i[k]) begin
        sum += values_i[k];
      end
    end
    return sum;
  endfunction : sum_value

  logic [Width-1:0] sum_value_exp;
  assign sum_value_exp = sum_value(values_i, valid_i);
  //VCS coverage on
  // pragma coverage on

  `ASSERT(ValidInImpliesValidOut_A, |valid_i === sum_valid_o)
  `ASSERT(SumComputation_A, sum_valid_o |-> sum_value_o == sum_value_exp)
  `ASSERT(SumComputationInvalid_A, !sum_valid_o |-> sum_value_o == '0)
`endif

endmodule : prim_sum_tree


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0


/**
 * Utility functions
 */
package prim_util_pkg;
  /**
   * Math function: $clog2 as specified in Verilog-2005
   *
   * Do not use this function if $clog2() is available.
   *
   * clog2 =          0        for value == 0
   *         ceil(log2(value)) for value >= 1
   *
   * This implementation is a synthesizable variant of the $clog2 function as
   * specified in the Verilog-2005 standard (IEEE 1364-2005).
   *
   * To quote the standard:
   *   The system function $clog2 shall return the ceiling of the log
   *   base 2 of the argument (the log rounded up to an integer
   *   value). The argument can be an integer or an arbitrary sized
   *   vector value. The argument shall be treated as an unsigned
   *   value, and an argument value of 0 shall produce a result of 0.
   */
  function automatic integer _clog2(integer value);
    integer result;
    // Use an intermediate value to avoid assigning to an input port, which produces a warning in
    // Synopsys DC.
    integer v = value;
    v = v - 1;
    for (result = 0; v > 0; result++) begin
      v = v >> 1;
    end
    return result;
  endfunction


  /**
   * Math function: Number of bits needed to address |value| items.
   *
   *                  0        for value == 0
   * vbits =          1        for value == 1
   *         ceil(log2(value)) for value > 1
   *
   *
   * The primary use case for this function is the definition of registers/arrays
   * which are wide enough to contain |value| items.
   *
   * This function identical to $clog2() for all input values except the value 1;
   * it could be considered an "enhanced" $clog2() function.
   *
   *
   * Example 1:
   *   parameter Items = 1;
   *   localparam ItemsWidth = vbits(Items); // 1
   *   logic [ItemsWidth-1:0] item_register; // items_register is now [0:0]
   *
   * Example 2:
   *   parameter Items = 64;
   *   localparam ItemsWidth = vbits(Items); // 6
   *   logic [ItemsWidth-1:0] item_register; // items_register is now [5:0]
   *
   * Note: If you want to store the number "value" inside a register, you need
   * a register with size vbits(value + 1), since you also need to store
   * the number 0.
   *
   * Example 3:
   *   logic [vbits(64)-1:0]     store_64_logic_values; // width is [5:0]
   *   logic [vbits(64 + 1)-1:0] store_number_64;       // width is [6:0]
   */
  function automatic integer vbits(integer value);
`ifdef XCELIUM
    // The use of system functions was not allowed here in Verilog-2001, but is
    // valid since (System)Verilog-2005, which is also when $clog2() first
    // appeared.
    // Xcelium < 19.10 does not yet support the use of $clog2() here, fall back
    // to an implementation without a system function. Remove this workaround
    // if we require a newer Xcelium version.
    // See #2579 and #2597.
    return (value == 1) ? 1 : _clog2(value);
`else
    return (value == 1) ? 1 : $clog2(value);
`endif
  endfunction

`ifdef INC_ASSERT
  // Package-scoped variable to detect the end of simulation.
  //
  // Used only in DV simulations. The bit will be used by assertions in RTL to perform end-of-test
  // cleanup. It is set to 1 in `dv_test_status_pkg::dv_test_status()`, which is invoked right
  // before the simulation is terminated, to signal the status of the test.
  bit end_of_simulation;
`endif

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module implements XoShiRo256++ PRNG
//
// Additional Entropy input to XOR fresh entropy into the state.
// Lockup protection that reseeds the generator if it falls into the all-zero state.
//
// Refs: [1] D. Blackman and S. Vigna, Scrambled Linear Pseudorndom Number Generators
//           https://arxiv.org/pdf/1805.01407.pdf
//       [2] https://prng.di.unimi.it/
//       [3] https://en.wikipedia.org/wiki/Xorshift#xoshiro_and_xoroshiro

`include "prim_assert.sv"

module prim_xoshiro256pp #(
  // Output width, must be a multiple of 64
  parameter int unsigned       OutputDw       = 64,
  // PRNG reset state, must be nonzero!
  parameter logic [255:0]      DefaultSeed    = 256'(1'b1),

  parameter int unsigned NumStages = OutputDw / 64 // derived parameter
) (
  input  logic                  clk_i,
  input  logic                  rst_ni,
  input  logic                  seed_en_i,    // load external seed into the state
  input  logic [255:0]          seed_i,       // external seed input
  input  logic                  xoshiro_en_i, // enables the PRNG
  input  logic [255:0]          entropy_i,    // additional entropy to be XOR'ed into the state
  output logic [OutputDw-1:0]   data_o,       // PRNG output
  output logic                  all_zero_o   // alert signal indicates the all-zero state
);

  logic [255:0] unrolled_state [NumStages+1];
  logic [63:0] mid [NumStages];

  logic lockup;
  logic [255:0] xoshiro_d, xoshiro_q, next_xoshiro_state;

  function automatic logic [255:0] state_update (input logic [255:0] data_in);
    logic [63:0] a_in, b_in, c_in, d_in;
    logic [63:0] a_out, b_out, c_out, d_out;
    a_in = data_in[255:192];
    b_in = data_in[191:128];
    c_in = data_in[127:64];
    d_in = data_in[63:0];
    a_out = a_in ^ b_in ^ d_in;
    b_out = a_in ^ b_in ^ c_in;
    c_out = a_in ^ (b_in << 17) ^ c_in;
    d_out = {d_in[18:0], d_in[63:19]} ^ {b_in[18:0], b_in[63:19]};
    return {a_out, b_out, c_out, d_out};
  endfunction: state_update

  assign unrolled_state[0] = xoshiro_q;

  for (genvar k = 0; k < NumStages; k++) begin : gen_state_functions
    // State update function
    assign unrolled_state[k+1] = state_update(unrolled_state[k]);
    // State output function
    assign mid[k] = unrolled_state[k][255:192] + unrolled_state[k][63:0];
    assign data_o[(k+1)*64-1:k*64] = {mid[k][40:0], mid[k][63:41]} + unrolled_state[k][255:192];
  end

  assign next_xoshiro_state = entropy_i ^ unrolled_state[NumStages];
  assign xoshiro_d = (seed_en_i)              ? seed_i             :
                     (xoshiro_en_i && lockup) ? DefaultSeed        :
                     (xoshiro_en_i)           ? next_xoshiro_state : xoshiro_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_reg_state
    if (!rst_ni) begin
      xoshiro_q <= DefaultSeed;
    end else begin
      xoshiro_q <= xoshiro_d;
    end
  end

  // lockup condition is all-zero
  assign lockup = ~(|xoshiro_q);

  // Indicate that the state is all zeros.
  assign all_zero_o = lockup;

  // check that seed is not all-zero
  `ASSERT_INIT(DefaultSeedNzCheck_A, |DefaultSeed)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package lc_ctrl_reg_pkg;

  // Param list
  parameter int SiliconCreatorIdWidth = 16;
  parameter int ProductIdWidth = 16;
  parameter int RevisionIdWidth = 8;
  parameter int NumTokenWords = 4;
  parameter int CsrLcStateWidth = 30;
  parameter int CsrLcCountWidth = 5;
  parameter int CsrLcIdStateWidth = 32;
  parameter int CsrOtpTestCtrlWidth = 32;
  parameter int CsrOtpTestStatusWidth = 32;
  parameter int NumDeviceIdWords = 8;
  parameter int NumManufStateWords = 8;
  parameter int NumAlerts = 3;

  // Address widths within the block
  parameter int BlockAw = 8;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } fatal_prog_error;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_state_error;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_bus_integ_error;
  } lc_ctrl_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic [7:0]  q;
    logic        qe;
  } lc_ctrl_reg2hw_claim_transition_if_reg_t;

  typedef struct packed {
    logic        q;
    logic        qe;
  } lc_ctrl_reg2hw_transition_cmd_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } ext_clock_en;
    struct packed {
      logic        q;
      logic        qe;
    } volatile_raw_unlock;
  } lc_ctrl_reg2hw_transition_ctrl_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } lc_ctrl_reg2hw_transition_token_mreg_t;

  typedef struct packed {
    logic [29:0] q;
    logic        qe;
  } lc_ctrl_reg2hw_transition_target_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } lc_ctrl_reg2hw_otp_vendor_test_ctrl_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } initialized;
    struct packed {
      logic        d;
    } ready;
    struct packed {
      logic        d;
    } ext_clock_switched;
    struct packed {
      logic        d;
    } transition_successful;
    struct packed {
      logic        d;
    } transition_count_error;
    struct packed {
      logic        d;
    } transition_error;
    struct packed {
      logic        d;
    } token_error;
    struct packed {
      logic        d;
    } flash_rma_error;
    struct packed {
      logic        d;
    } otp_error;
    struct packed {
      logic        d;
    } state_error;
    struct packed {
      logic        d;
    } bus_integ_error;
    struct packed {
      logic        d;
    } otp_partition_error;
  } lc_ctrl_hw2reg_status_reg_t;

  typedef struct packed {
    logic [7:0]  d;
  } lc_ctrl_hw2reg_claim_transition_if_reg_t;

  typedef struct packed {
    logic        d;
  } lc_ctrl_hw2reg_transition_regwen_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } ext_clock_en;
    struct packed {
      logic        d;
    } volatile_raw_unlock;
  } lc_ctrl_hw2reg_transition_ctrl_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } lc_ctrl_hw2reg_transition_token_mreg_t;

  typedef struct packed {
    logic [29:0] d;
  } lc_ctrl_hw2reg_transition_target_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } lc_ctrl_hw2reg_otp_vendor_test_ctrl_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } lc_ctrl_hw2reg_otp_vendor_test_status_reg_t;

  typedef struct packed {
    logic [29:0] d;
  } lc_ctrl_hw2reg_lc_state_reg_t;

  typedef struct packed {
    logic [4:0]  d;
  } lc_ctrl_hw2reg_lc_transition_cnt_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } lc_ctrl_hw2reg_lc_id_state_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } product_id;
    struct packed {
      logic [15:0] d;
    } silicon_creator_id;
  } lc_ctrl_hw2reg_hw_revision0_reg_t;

  typedef struct packed {
    struct packed {
      logic [7:0]  d;
    } revision_id;
    struct packed {
      logic [23:0] d;
    } reserved;
  } lc_ctrl_hw2reg_hw_revision1_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } lc_ctrl_hw2reg_device_id_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } lc_ctrl_hw2reg_manuf_state_mreg_t;

  // Register -> HW type
  typedef struct packed {
    lc_ctrl_reg2hw_alert_test_reg_t alert_test; // [216:211]
    lc_ctrl_reg2hw_claim_transition_if_reg_t claim_transition_if; // [210:202]
    lc_ctrl_reg2hw_transition_cmd_reg_t transition_cmd; // [201:200]
    lc_ctrl_reg2hw_transition_ctrl_reg_t transition_ctrl; // [199:196]
    lc_ctrl_reg2hw_transition_token_mreg_t [3:0] transition_token; // [195:64]
    lc_ctrl_reg2hw_transition_target_reg_t transition_target; // [63:33]
    lc_ctrl_reg2hw_otp_vendor_test_ctrl_reg_t otp_vendor_test_ctrl; // [32:0]
  } lc_ctrl_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    lc_ctrl_hw2reg_status_reg_t status; // [887:876]
    lc_ctrl_hw2reg_claim_transition_if_reg_t claim_transition_if; // [875:868]
    lc_ctrl_hw2reg_transition_regwen_reg_t transition_regwen; // [867:867]
    lc_ctrl_hw2reg_transition_ctrl_reg_t transition_ctrl; // [866:865]
    lc_ctrl_hw2reg_transition_token_mreg_t [3:0] transition_token; // [864:737]
    lc_ctrl_hw2reg_transition_target_reg_t transition_target; // [736:707]
    lc_ctrl_hw2reg_otp_vendor_test_ctrl_reg_t otp_vendor_test_ctrl; // [706:675]
    lc_ctrl_hw2reg_otp_vendor_test_status_reg_t otp_vendor_test_status; // [674:643]
    lc_ctrl_hw2reg_lc_state_reg_t lc_state; // [642:613]
    lc_ctrl_hw2reg_lc_transition_cnt_reg_t lc_transition_cnt; // [612:608]
    lc_ctrl_hw2reg_lc_id_state_reg_t lc_id_state; // [607:576]
    lc_ctrl_hw2reg_hw_revision0_reg_t hw_revision0; // [575:544]
    lc_ctrl_hw2reg_hw_revision1_reg_t hw_revision1; // [543:512]
    lc_ctrl_hw2reg_device_id_mreg_t [7:0] device_id; // [511:256]
    lc_ctrl_hw2reg_manuf_state_mreg_t [7:0] manuf_state; // [255:0]
  } lc_ctrl_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] LC_CTRL_ALERT_TEST_OFFSET = 8'h 0;
  parameter logic [BlockAw-1:0] LC_CTRL_STATUS_OFFSET = 8'h 4;
  parameter logic [BlockAw-1:0] LC_CTRL_CLAIM_TRANSITION_IF_REGWEN_OFFSET = 8'h 8;
  parameter logic [BlockAw-1:0] LC_CTRL_CLAIM_TRANSITION_IF_OFFSET = 8'h c;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_REGWEN_OFFSET = 8'h 10;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_CMD_OFFSET = 8'h 14;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_CTRL_OFFSET = 8'h 18;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_TOKEN_0_OFFSET = 8'h 1c;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_TOKEN_1_OFFSET = 8'h 20;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_TOKEN_2_OFFSET = 8'h 24;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_TOKEN_3_OFFSET = 8'h 28;
  parameter logic [BlockAw-1:0] LC_CTRL_TRANSITION_TARGET_OFFSET = 8'h 2c;
  parameter logic [BlockAw-1:0] LC_CTRL_OTP_VENDOR_TEST_CTRL_OFFSET = 8'h 30;
  parameter logic [BlockAw-1:0] LC_CTRL_OTP_VENDOR_TEST_STATUS_OFFSET = 8'h 34;
  parameter logic [BlockAw-1:0] LC_CTRL_LC_STATE_OFFSET = 8'h 38;
  parameter logic [BlockAw-1:0] LC_CTRL_LC_TRANSITION_CNT_OFFSET = 8'h 3c;
  parameter logic [BlockAw-1:0] LC_CTRL_LC_ID_STATE_OFFSET = 8'h 40;
  parameter logic [BlockAw-1:0] LC_CTRL_HW_REVISION0_OFFSET = 8'h 44;
  parameter logic [BlockAw-1:0] LC_CTRL_HW_REVISION1_OFFSET = 8'h 48;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_0_OFFSET = 8'h 4c;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_1_OFFSET = 8'h 50;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_2_OFFSET = 8'h 54;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_3_OFFSET = 8'h 58;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_4_OFFSET = 8'h 5c;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_5_OFFSET = 8'h 60;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_6_OFFSET = 8'h 64;
  parameter logic [BlockAw-1:0] LC_CTRL_DEVICE_ID_7_OFFSET = 8'h 68;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_0_OFFSET = 8'h 6c;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_1_OFFSET = 8'h 70;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_2_OFFSET = 8'h 74;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_3_OFFSET = 8'h 78;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_4_OFFSET = 8'h 7c;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_5_OFFSET = 8'h 80;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_6_OFFSET = 8'h 84;
  parameter logic [BlockAw-1:0] LC_CTRL_MANUF_STATE_7_OFFSET = 8'h 88;

  // Reset values for hwext registers and their fields
  parameter logic [2:0] LC_CTRL_ALERT_TEST_RESVAL = 3'h 0;
  parameter logic [0:0] LC_CTRL_ALERT_TEST_FATAL_PROG_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] LC_CTRL_ALERT_TEST_FATAL_STATE_ERROR_RESVAL = 1'h 0;
  parameter logic [0:0] LC_CTRL_ALERT_TEST_FATAL_BUS_INTEG_ERROR_RESVAL = 1'h 0;
  parameter logic [11:0] LC_CTRL_STATUS_RESVAL = 12'h 0;
  parameter logic [7:0] LC_CTRL_CLAIM_TRANSITION_IF_RESVAL = 8'h 69;
  parameter logic [7:0] LC_CTRL_CLAIM_TRANSITION_IF_MUTEX_RESVAL = 8'h 69;
  parameter logic [0:0] LC_CTRL_TRANSITION_REGWEN_RESVAL = 1'h 0;
  parameter logic [0:0] LC_CTRL_TRANSITION_REGWEN_TRANSITION_REGWEN_RESVAL = 1'h 0;
  parameter logic [0:0] LC_CTRL_TRANSITION_CMD_RESVAL = 1'h 0;
  parameter logic [1:0] LC_CTRL_TRANSITION_CTRL_RESVAL = 2'h 0;
  parameter logic [31:0] LC_CTRL_TRANSITION_TOKEN_0_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_TRANSITION_TOKEN_1_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_TRANSITION_TOKEN_2_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_TRANSITION_TOKEN_3_RESVAL = 32'h 0;
  parameter logic [29:0] LC_CTRL_TRANSITION_TARGET_RESVAL = 30'h 0;
  parameter logic [31:0] LC_CTRL_OTP_VENDOR_TEST_CTRL_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_OTP_VENDOR_TEST_STATUS_RESVAL = 32'h 0;
  parameter logic [29:0] LC_CTRL_LC_STATE_RESVAL = 30'h 0;
  parameter logic [4:0] LC_CTRL_LC_TRANSITION_CNT_RESVAL = 5'h 0;
  parameter logic [31:0] LC_CTRL_LC_ID_STATE_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_HW_REVISION0_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_HW_REVISION1_RESVAL = 32'h 0;
  parameter logic [23:0] LC_CTRL_HW_REVISION1_RESERVED_RESVAL = 24'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_0_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_1_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_2_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_3_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_4_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_5_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_6_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_DEVICE_ID_7_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_0_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_1_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_2_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_3_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_4_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_5_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_6_RESVAL = 32'h 0;
  parameter logic [31:0] LC_CTRL_MANUF_STATE_7_RESVAL = 32'h 0;

  // Register index
  typedef enum int {
    LC_CTRL_ALERT_TEST,
    LC_CTRL_STATUS,
    LC_CTRL_CLAIM_TRANSITION_IF_REGWEN,
    LC_CTRL_CLAIM_TRANSITION_IF,
    LC_CTRL_TRANSITION_REGWEN,
    LC_CTRL_TRANSITION_CMD,
    LC_CTRL_TRANSITION_CTRL,
    LC_CTRL_TRANSITION_TOKEN_0,
    LC_CTRL_TRANSITION_TOKEN_1,
    LC_CTRL_TRANSITION_TOKEN_2,
    LC_CTRL_TRANSITION_TOKEN_3,
    LC_CTRL_TRANSITION_TARGET,
    LC_CTRL_OTP_VENDOR_TEST_CTRL,
    LC_CTRL_OTP_VENDOR_TEST_STATUS,
    LC_CTRL_LC_STATE,
    LC_CTRL_LC_TRANSITION_CNT,
    LC_CTRL_LC_ID_STATE,
    LC_CTRL_HW_REVISION0,
    LC_CTRL_HW_REVISION1,
    LC_CTRL_DEVICE_ID_0,
    LC_CTRL_DEVICE_ID_1,
    LC_CTRL_DEVICE_ID_2,
    LC_CTRL_DEVICE_ID_3,
    LC_CTRL_DEVICE_ID_4,
    LC_CTRL_DEVICE_ID_5,
    LC_CTRL_DEVICE_ID_6,
    LC_CTRL_DEVICE_ID_7,
    LC_CTRL_MANUF_STATE_0,
    LC_CTRL_MANUF_STATE_1,
    LC_CTRL_MANUF_STATE_2,
    LC_CTRL_MANUF_STATE_3,
    LC_CTRL_MANUF_STATE_4,
    LC_CTRL_MANUF_STATE_5,
    LC_CTRL_MANUF_STATE_6,
    LC_CTRL_MANUF_STATE_7
  } lc_ctrl_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] LC_CTRL_PERMIT [35] = '{
    4'b 0001, // index[ 0] LC_CTRL_ALERT_TEST
    4'b 0011, // index[ 1] LC_CTRL_STATUS
    4'b 0001, // index[ 2] LC_CTRL_CLAIM_TRANSITION_IF_REGWEN
    4'b 0001, // index[ 3] LC_CTRL_CLAIM_TRANSITION_IF
    4'b 0001, // index[ 4] LC_CTRL_TRANSITION_REGWEN
    4'b 0001, // index[ 5] LC_CTRL_TRANSITION_CMD
    4'b 0001, // index[ 6] LC_CTRL_TRANSITION_CTRL
    4'b 1111, // index[ 7] LC_CTRL_TRANSITION_TOKEN_0
    4'b 1111, // index[ 8] LC_CTRL_TRANSITION_TOKEN_1
    4'b 1111, // index[ 9] LC_CTRL_TRANSITION_TOKEN_2
    4'b 1111, // index[10] LC_CTRL_TRANSITION_TOKEN_3
    4'b 1111, // index[11] LC_CTRL_TRANSITION_TARGET
    4'b 1111, // index[12] LC_CTRL_OTP_VENDOR_TEST_CTRL
    4'b 1111, // index[13] LC_CTRL_OTP_VENDOR_TEST_STATUS
    4'b 1111, // index[14] LC_CTRL_LC_STATE
    4'b 0001, // index[15] LC_CTRL_LC_TRANSITION_CNT
    4'b 1111, // index[16] LC_CTRL_LC_ID_STATE
    4'b 1111, // index[17] LC_CTRL_HW_REVISION0
    4'b 1111, // index[18] LC_CTRL_HW_REVISION1
    4'b 1111, // index[19] LC_CTRL_DEVICE_ID_0
    4'b 1111, // index[20] LC_CTRL_DEVICE_ID_1
    4'b 1111, // index[21] LC_CTRL_DEVICE_ID_2
    4'b 1111, // index[22] LC_CTRL_DEVICE_ID_3
    4'b 1111, // index[23] LC_CTRL_DEVICE_ID_4
    4'b 1111, // index[24] LC_CTRL_DEVICE_ID_5
    4'b 1111, // index[25] LC_CTRL_DEVICE_ID_6
    4'b 1111, // index[26] LC_CTRL_DEVICE_ID_7
    4'b 1111, // index[27] LC_CTRL_MANUF_STATE_0
    4'b 1111, // index[28] LC_CTRL_MANUF_STATE_1
    4'b 1111, // index[29] LC_CTRL_MANUF_STATE_2
    4'b 1111, // index[30] LC_CTRL_MANUF_STATE_3
    4'b 1111, // index[31] LC_CTRL_MANUF_STATE_4
    4'b 1111, // index[32] LC_CTRL_MANUF_STATE_5
    4'b 1111, // index[33] LC_CTRL_MANUF_STATE_6
    4'b 1111  // index[34] LC_CTRL_MANUF_STATE_7
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Life cycle state encoding definition.
//
// DO NOT EDIT THIS FILE DIRECTLY.
// It has been generated with
// $ ./util/design/gen-lc-state-enc.py --seed 10167336684108184581
//
package lc_ctrl_state_pkg;

  import prim_util_pkg::vbits;

  ///////////////////////////////
  // General size declarations //
  ///////////////////////////////

  parameter int LcValueWidth = 16;

  parameter int NumLcStateValues = 20;
  parameter int LcStateWidth = NumLcStateValues * LcValueWidth;
  parameter int NumLcStates = 21;
  parameter int DecLcStateWidth = vbits(NumLcStates);
  // Redundant version used in the CSRs.
  parameter int DecLcStateNumRep = 32/DecLcStateWidth;
  parameter int ExtDecLcStateWidth = DecLcStateNumRep*DecLcStateWidth;

  parameter int NumLcCountValues = 24;
  parameter int LcCountWidth = NumLcCountValues * LcValueWidth;
  parameter int NumLcCountStates = 25;
  parameter int DecLcCountWidth = vbits(NumLcCountStates);

  // This state is not stored in OTP, but inferred from the locked
  // status of the secret partitions. Hence, only the decoded ID state
  // is declared here for exposure through the CSR interface.
  parameter int NumLcIdStates = 2;
  parameter int DecLcIdStateWidth = vbits(NumLcIdStates+1);
  // Redundant version used in the CSRs.
  parameter int DecLcIdStateNumRep = 32/DecLcIdStateWidth;
  parameter int ExtDecLcIdStateWidth = DecLcIdStateNumRep*DecLcIdStateWidth;

  /////////////////////////////////////////////
  // Life cycle manufacturing state encoding //
  /////////////////////////////////////////////

  // These values have been generated such that they are incrementally writeable with respect
  // to the ECC polynomial specified. The values are used to define the life cycle manufacturing
  // state and transition counter encoding in lc_ctrl_pkg.sv.
  //
  // The values are unique and have the following statistics (considering all 16
  // data and 6 ECC bits):
  //
  // - Minimum Hamming weight: 6
  // - Maximum Hamming weight: 16
  // - Minimum Hamming distance from any other value: 6
  // - Maximum Hamming distance from any other value: 20
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: --
  //  6: ||| (5.90%)
  //  7: --
  //  8: |||||||||| (16.14%)
  //  9: --
  // 10: |||||||||||||||||||| (30.15%)
  // 11: --
  // 12: |||||||||||||||||| (28.45%)
  // 13: --
  // 14: |||||||||| (15.10%)
  // 15: --
  // 16: || (3.87%)
  // 17: --
  // 18:  (0.37%)
  // 19: --
  // 20:  (0.03%)
  // 21: --
  // 22: --
  //
  //
  // Note that the ECC bits are not defined in this package as they will be calculated by
  // the OTP ECC logic at runtime.

  // SEC_CM: MANUF.STATE.SPARSE
  // The A/B values are used for the encoded LC state.
  parameter logic [15:0] A0 = 16'b0001011010010010; // ECC: 6'b110011
  parameter logic [15:0] B0 = 16'b1001111111110010; // ECC: 6'b111011

  parameter logic [15:0] A1 = 16'b1011000000101110; // ECC: 6'b011010
  parameter logic [15:0] B1 = 16'b1011010000111111; // ECC: 6'b111111

  parameter logic [15:0] A2 = 16'b1110001000010001; // ECC: 6'b110110
  parameter logic [15:0] B2 = 16'b1110001100011111; // ECC: 6'b111111

  parameter logic [15:0] A3 = 16'b1100100110010000; // ECC: 6'b011000
  parameter logic [15:0] B3 = 16'b1111110111010010; // ECC: 6'b111000

  parameter logic [15:0] A4 = 16'b0000111100100001; // ECC: 6'b010100
  parameter logic [15:0] B4 = 16'b1010111110100111; // ECC: 6'b111101

  parameter logic [15:0] A5 = 16'b1101010010110001; // ECC: 6'b110000
  parameter logic [15:0] B5 = 16'b1101011011111111; // ECC: 6'b110001

  parameter logic [15:0] A6 = 16'b0010101100110000; // ECC: 6'b100010
  parameter logic [15:0] B6 = 16'b1010101101110110; // ECC: 6'b111111

  parameter logic [15:0] A7 = 16'b0011110100110010; // ECC: 6'b010100
  parameter logic [15:0] B7 = 16'b1111111110110011; // ECC: 6'b110100

  parameter logic [15:0] A8 = 16'b1110100010110000; // ECC: 6'b101100
  parameter logic [15:0] B8 = 16'b1110111010111010; // ECC: 6'b101111

  parameter logic [15:0] A9 = 16'b1111010000011101; // ECC: 6'b000100
  parameter logic [15:0] B9 = 16'b1111010011111111; // ECC: 6'b101100

  parameter logic [15:0] A10 = 16'b1001100110100101; // ECC: 6'b011000
  parameter logic [15:0] B10 = 16'b1111111110100101; // ECC: 6'b011110

  parameter logic [15:0] A11 = 16'b1110010010000101; // ECC: 6'b110100
  parameter logic [15:0] B11 = 16'b1110010011101111; // ECC: 6'b110111

  parameter logic [15:0] A12 = 16'b0100100101110111; // ECC: 6'b100000
  parameter logic [15:0] B12 = 16'b0100111111111111; // ECC: 6'b101010

  parameter logic [15:0] A13 = 16'b0010110001110011; // ECC: 6'b000011
  parameter logic [15:0] B13 = 16'b1011111001111111; // ECC: 6'b001011

  parameter logic [15:0] A14 = 16'b1001000101101100; // ECC: 6'b101010
  parameter logic [15:0] B14 = 16'b1001110111101101; // ECC: 6'b111011

  parameter logic [15:0] A15 = 16'b0011000000001101; // ECC: 6'b100011
  parameter logic [15:0] B15 = 16'b1111001011011111; // ECC: 6'b100111

  parameter logic [15:0] A16 = 16'b1010011000010101; // ECC: 6'b001011
  parameter logic [15:0] B16 = 16'b1011011110011101; // ECC: 6'b011111

  parameter logic [15:0] A17 = 16'b0110000100101110; // ECC: 6'b000100
  parameter logic [15:0] B17 = 16'b1110010101111110; // ECC: 6'b011100

  parameter logic [15:0] A18 = 16'b1100001110110000; // ECC: 6'b001101
  parameter logic [15:0] B18 = 16'b1101001110110111; // ECC: 6'b011111

  parameter logic [15:0] A19 = 16'b1100000110000011; // ECC: 6'b000110
  parameter logic [15:0] B19 = 16'b1110010111010111; // ECC: 6'b111110


  // SEC_CM: TRANSITION.CTR.SPARSE
  // The C/D values are used for the encoded LC transition counter.
  parameter logic [15:0] C0 = 16'b1111000000100100; // ECC: 6'b001100
  parameter logic [15:0] D0 = 16'b1111110000111100; // ECC: 6'b111100

  parameter logic [15:0] C1 = 16'b0010000110000011; // ECC: 6'b110100
  parameter logic [15:0] D1 = 16'b0010001111111011; // ECC: 6'b110101

  parameter logic [15:0] C2 = 16'b1111100011000100; // ECC: 6'b110000
  parameter logic [15:0] D2 = 16'b1111100111101110; // ECC: 6'b110101

  parameter logic [15:0] C3 = 16'b1010110000011000; // ECC: 6'b110110
  parameter logic [15:0] D3 = 16'b1010110110011111; // ECC: 6'b110111

  parameter logic [15:0] C4 = 16'b0101001101001101; // ECC: 6'b001100
  parameter logic [15:0] D4 = 16'b0111111101101111; // ECC: 6'b001110

  parameter logic [15:0] C5 = 16'b0100010011010010; // ECC: 6'b110000
  parameter logic [15:0] D5 = 16'b0100010011111011; // ECC: 6'b111110

  parameter logic [15:0] C6 = 16'b1100010010100100; // ECC: 6'b101110
  parameter logic [15:0] D6 = 16'b1100111011100110; // ECC: 6'b111111

  parameter logic [15:0] C7 = 16'b0001111001100011; // ECC: 6'b000101
  parameter logic [15:0] D7 = 16'b0101111001111011; // ECC: 6'b011111

  parameter logic [15:0] C8 = 16'b0110010110010000; // ECC: 6'b000000
  parameter logic [15:0] D8 = 16'b0111011111010100; // ECC: 6'b010001

  parameter logic [15:0] C9 = 16'b0010001101100100; // ECC: 6'b010111
  parameter logic [15:0] D9 = 16'b1110011101100111; // ECC: 6'b011111

  parameter logic [15:0] C10 = 16'b0100101100000000; // ECC: 6'b000110
  parameter logic [15:0] D10 = 16'b1100101101010011; // ECC: 6'b110111

  parameter logic [15:0] C11 = 16'b1011101010000001; // ECC: 6'b000100
  parameter logic [15:0] D11 = 16'b1111111010101011; // ECC: 6'b010111

  parameter logic [15:0] C12 = 16'b0101101110101010; // ECC: 6'b010000
  parameter logic [15:0] D12 = 16'b0101111110111111; // ECC: 6'b010011

  parameter logic [15:0] C13 = 16'b0010110001101001; // ECC: 6'b001000
  parameter logic [15:0] D13 = 16'b0110111011101001; // ECC: 6'b011110

  parameter logic [15:0] C14 = 16'b1111001000010011; // ECC: 6'b100001
  parameter logic [15:0] D14 = 16'b1111001101110111; // ECC: 6'b101011

  parameter logic [15:0] C15 = 16'b0001110111110010; // ECC: 6'b100000
  parameter logic [15:0] D15 = 16'b0101110111110011; // ECC: 6'b110111

  parameter logic [15:0] C16 = 16'b1001101101100000; // ECC: 6'b110100
  parameter logic [15:0] D16 = 16'b1001111101101111; // ECC: 6'b111100

  parameter logic [15:0] C17 = 16'b0101111001101000; // ECC: 6'b110000
  parameter logic [15:0] D17 = 16'b1111111101101000; // ECC: 6'b111011

  parameter logic [15:0] C18 = 16'b0101110111000100; // ECC: 6'b010100
  parameter logic [15:0] D18 = 16'b0101110111011110; // ECC: 6'b011111

  parameter logic [15:0] C19 = 16'b0000010000000101; // ECC: 6'b101010
  parameter logic [15:0] D19 = 16'b0110010001010101; // ECC: 6'b101111

  parameter logic [15:0] C20 = 16'b0111011000101000; // ECC: 6'b011001
  parameter logic [15:0] D20 = 16'b0111011010111110; // ECC: 6'b011111

  parameter logic [15:0] C21 = 16'b0110001011101000; // ECC: 6'b100011
  parameter logic [15:0] D21 = 16'b0110101111111101; // ECC: 6'b110011

  parameter logic [15:0] C22 = 16'b1000101110001010; // ECC: 6'b101001
  parameter logic [15:0] D22 = 16'b1000111111111011; // ECC: 6'b101101

  parameter logic [15:0] C23 = 16'b1101000000001101; // ECC: 6'b010001
  parameter logic [15:0] D23 = 16'b1111101111001101; // ECC: 6'b010111


  parameter logic [15:0] ZRO = 16'h0;

  ////////////////////////
  // Derived enum types //
  ////////////////////////

  // Use lc_state_t and lc_cnt_t in interfaces as very wide enumerations ( > 64 bits )
  // are not supported for virtual interfaces by Excelium yet
  // https://github.com/lowRISC/opentitan/issues/8884 (Cadence issue: cds_46570160)
  // The enumeration types lc_state_e and lc_cnt_e are still ok in other circumstances

  typedef logic [LcStateWidth-1:0] lc_state_t;
  typedef enum lc_state_t {
    LcStRaw           = {ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO},
    LcStTestUnlocked0 = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  A3,  A2,  A1,  B0},
    LcStTestLocked0   = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  A3,  A2,  B1,  B0},
    LcStTestUnlocked1 = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  A3,  B2,  B1,  B0},
    LcStTestLocked1   = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  A6,  A5,  A4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked2 = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  A6,  A5,  B4,  B3,  B2,  B1,  B0},
    LcStTestLocked2   = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  A6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked3 = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  A7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestLocked3   = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  A8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked4 = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  A9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestLocked4   = {A19, A18, A17, A16, A15, A14, A13, A12, A11, A10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked5 = {A19, A18, A17, A16, A15, A14, A13, A12, A11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestLocked5   = {A19, A18, A17, A16, A15, A14, A13, A12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked6 = {A19, A18, A17, A16, A15, A14, A13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestLocked6   = {A19, A18, A17, A16, A15, A14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStTestUnlocked7 = {A19, A18, A17, A16, A15, B14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStDev           = {A19, A18, A17, A16, B15, B14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStProd          = {A19, A18, A17, B16, A15, B14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStProdEnd       = {A19, A18, B17, A16, A15, B14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStRma           = {B19, B18, A17, B16, B15, B14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0},
    LcStScrap         = {B19, B18, B17, B16, B15, B14, B13, B12, B11, B10,  B9,  B8,  B7,  B6,  B5,  B4,  B3,  B2,  B1,  B0}
  } lc_state_e;

  typedef logic [LcCountWidth-1:0] lc_cnt_t;
  typedef enum lc_cnt_t {
    LcCnt0  = {ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO, ZRO},
    LcCnt1  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  C3,  C2,  C1,  D0},
    LcCnt2  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  C3,  C2,  D1,  D0},
    LcCnt3  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  C3,  D2,  D1,  D0},
    LcCnt4  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  C4,  D3,  D2,  D1,  D0},
    LcCnt5  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  C5,  D4,  D3,  D2,  D1,  D0},
    LcCnt6  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  C6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt7  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  C7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt8  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  C8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt9  = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  C9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt10 = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, C10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt11 = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, C11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt12 = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, C12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt13 = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, C13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt14 = {C23, C22, C21, C20, C19, C18, C17, C16, C15, C14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt15 = {C23, C22, C21, C20, C19, C18, C17, C16, C15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt16 = {C23, C22, C21, C20, C19, C18, C17, C16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt17 = {C23, C22, C21, C20, C19, C18, C17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt18 = {C23, C22, C21, C20, C19, C18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt19 = {C23, C22, C21, C20, C19, D18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt20 = {C23, C22, C21, C20, D19, D18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt21 = {C23, C22, C21, D20, D19, D18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt22 = {C23, C22, D21, D20, D19, D18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt23 = {C23, D22, D21, D20, D19, D18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0},
    LcCnt24 = {D23, D22, D21, D20, D19, D18, D17, D16, D15, D14, D13, D12, D11, D10,  D9,  D8,  D7,  D6,  D5,  D4,  D3,  D2,  D1,  D0}
  } lc_cnt_e;

  // Decoded life cycle state, used to interface with CSRs and TAP.
  typedef enum logic [DecLcStateWidth-1:0] {
    DecLcStRaw = 0,
    DecLcStTestUnlocked0 = 1,
    DecLcStTestLocked0 = 2,
    DecLcStTestUnlocked1 = 3,
    DecLcStTestLocked1 = 4,
    DecLcStTestUnlocked2 = 5,
    DecLcStTestLocked2 = 6,
    DecLcStTestUnlocked3 = 7,
    DecLcStTestLocked3 = 8,
    DecLcStTestUnlocked4 = 9,
    DecLcStTestLocked4 = 10,
    DecLcStTestUnlocked5 = 11,
    DecLcStTestLocked5 = 12,
    DecLcStTestUnlocked6 = 13,
    DecLcStTestLocked6 = 14,
    DecLcStTestUnlocked7 = 15,
    DecLcStDev = 16,
    DecLcStProd = 17,
    DecLcStProdEnd = 18,
    DecLcStRma = 19,
    DecLcStScrap = 20,
    DecLcStPostTrans = 21,
    DecLcStEscalate = 22,
    DecLcStInvalid = 23
  } dec_lc_state_e;

  typedef dec_lc_state_e [DecLcStateNumRep-1:0] ext_dec_lc_state_t;

  typedef enum logic [DecLcIdStateWidth-1:0] {
    DecLcIdBlank,
    DecLcIdPersonalized,
    DecLcIdInvalid
  } dec_lc_id_state_e;

  typedef logic [DecLcCountWidth-1:0] dec_lc_cnt_t;


  ///////////////////////////////////////////
  // Hashed RAW unlock and all-zero tokens //
  ///////////////////////////////////////////

  parameter int LcTokenWidth = 128;
  typedef logic [LcTokenWidth-1:0] lc_token_t;

  parameter lc_token_t AllZeroToken = {
    128'h0
  };
  parameter lc_token_t RndCnstRawUnlockToken = {
    128'h51E6121C8694C6BC41F36E2175199296
  };
  parameter lc_token_t AllZeroTokenHashed = {
    128'h3852305BAECF5FF1D5C1D25F6DB9058D
  };
  parameter lc_token_t RndCnstRawUnlockTokenHashed = {
    128'hC1E437642C17A6A2C744CCF32509B8A5
  };

endpackage : lc_ctrl_state_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_clock_mux2

#(

  parameter bit NoFpgaBufG = 1'b0 // this parameter serves no function in the generic model

) (
  input        clk0_i,
  input        clk1_i,
  input        sel_i,
  output logic clk_o
);

  if (1) begin : gen_generic
    prim_generic_clock_mux2 #(
      .NoFpgaBufG(NoFpgaBufG)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_pad_wrapper
import prim_pad_wrapper_pkg::*;
#(

  // These parameters are ignored in this model.
  parameter pad_type_e PadType = BidirStd,
  parameter scan_role_e ScanRole = NoScan

) (
  // This is only used for scanmode (not used in generic models)
  input              clk_scan_i,
  input              scanmode_i,
  // Power sequencing signals (not used in generic models)
  input pad_pok_t    pok_i,
  // Main Pad signals
  inout wire         inout_io, // bidirectional pad
  output logic       in_o,     // input data
  output logic       in_raw_o, // uninverted output data
  input              ie_i,     // input enable
  input              out_i,    // output data
  input              oe_i,     // output enable
  input pad_attr_t   attr_i    // additional pad attributes
);

  if (1) begin : gen_generic
    prim_generic_pad_wrapper #(
      .PadType(PadType),
      .ScanRole(ScanRole)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_ram_1p
import prim_ram_1p_pkg::*;
#(

  parameter  int Width           = 32, // bit
  parameter  int Depth           = 128,
  parameter  int DataBitsPerMask = 1, // Number of data bits per bit of write mask
  parameter      MemInitFile     = "", // VMEM file to initialize the memory with

  localparam int Aw              = $clog2(Depth)  // derived parameter

) (
  input  logic             clk_i,

  input  logic             req_i,
  input  logic             write_i,
  input  logic [Aw-1:0]    addr_i,
  input  logic [Width-1:0] wdata_i,
  input  logic [Width-1:0] wmask_i,
  output logic [Width-1:0] rdata_o, // Read data. Data is returned one cycle after req_i is high.
  input ram_1p_cfg_t       cfg_i
);

  if (1) begin : gen_generic
    prim_generic_ram_1p #(
      .DataBitsPerMask(DataBitsPerMask),
      .Depth(Depth),
      .MemInitFile(MemInitFile),
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_rom
import prim_rom_pkg::*;
#(

  parameter  int Width       = 32,
  parameter  int Depth       = 2048, // 8kB default
  parameter      MemInitFile = "", // VMEM file to initialize the memory with

  localparam int Aw          = $clog2(Depth)

) (
  input  logic             clk_i,
  input  logic             req_i,
  input  logic [Aw-1:0]    addr_i,
  output logic [Width-1:0] rdata_o,
  input rom_cfg_t          cfg_i
);

  if (1) begin : gen_generic
    prim_generic_rom #(
      .Depth(Depth),
      .MemInitFile(MemInitFile),
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module prim_generic_flop_en #(
  parameter int               Width      = 1,
  parameter bit               EnSecBuf   = 0,
  parameter logic [Width-1:0] ResetValue = 0
) (
  input                    clk_i,
  input                    rst_ni,
  input                    en_i,
  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_o
);

  logic en;
  if (EnSecBuf) begin : gen_en_sec_buf
    prim_sec_anchor_buf #(
      .Width(1)
    ) u_en_buf (
      .in_i(en_i),
      .out_o(en)
    );
  end else begin : gen_en_no_sec_buf
    assign en = en_i;
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      q_o <= ResetValue;
    end else if (en) begin
      q_o <= d_i;
    end
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// One-hot encoder
// Outputs a one-hot encoded version of an integer input.

module prim_onehot_enc #(
  parameter int unsigned OneHotWidth = 32,
  localparam int unsigned InputWidth = $clog2(OneHotWidth)
) (
  input  logic [InputWidth-1:0]  in_i,
  input  logic                   en_i, // out_o == '0 when en_i == 0

  output logic [OneHotWidth-1:0] out_o
);

  for (genvar i = 0; i < OneHotWidth; ++i) begin : g_out
    assign out_o[i] = (in_i == i) & en_i;
  end
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// One-hot mux
// A AND/OR mux with a one-hot select input.

`include "prim_assert.sv"

module prim_onehot_mux #(
  parameter int Width  = 32,
  parameter int Inputs = 8
) (
  // Clock and reset only for assertions
  input clk_i,
  input rst_ni,

  input  logic [Width-1:0]  in_i [Inputs],
  input  logic [Inputs-1:0] sel_i, // Must be one-hot or zero
  output logic [Width-1:0]  out_o
);
  logic [Inputs-1:0] in_mux [Width];

  for (genvar b = 0; b < Width; ++b) begin : g_in_mux_outer
    logic [Inputs-1:0] out_mux_bits;

    for (genvar i = 0; i < Inputs; ++i) begin : g_in_mux_inner
      assign in_mux[b][i] = in_i[i][b];
    end

    prim_and2 #(.Width(Inputs)) u_mux_bit_and(
      .in0_i(in_mux[b]),
      .in1_i(sel_i),
      .out_o(out_mux_bits)
    );

    assign out_o[b] = |out_mux_bits;
  end

  logic unused_clk;
  logic unused_rst_n;

  // clock and reset only needed for assertion
  assign unused_clk   = clk_i;
  assign unused_rst_n = rst_ni;

  `ASSERT(SelIsOnehot_A, $onehot0(sel_i))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Onehot checker.
//
// This module checks whether the input vector oh_i is onehot0 and generates an error if not.
//
// Optionally, two additional checks can be activated:
//
// 1) EnableCheck: this check performs an OR reduction of the onehot vector, and compares
//    the result with en_i. If there is a mismatch, an error is generated.
// 2) AddrCheck: this checks whether the onehot bit is in the correct position.
//    It requires an additional address addr_i to be supplied to the module.
//
// All checks make use of an explicit binary tree implementation in order to minimize the delay.
//

`include "prim_assert.sv"

module prim_onehot_check #(
  parameter int unsigned AddrWidth   = 5,
  // The onehot width can be <= 2**AddrWidth and does not have to be a power of two.
  parameter int unsigned OneHotWidth = 2**AddrWidth,
  // If set to 0, the addr_i input will not be used for the check and can be tied off.
  parameter bit          AddrCheck   = 1,
  // If set to 0, the en_i value will not be used for the check and can be tied off.
  parameter bit          EnableCheck = 1,
  // If set to 1, the oh_i vector must always be one hot if en_i is set to 1.
  // If set to 0, the oh_i vector may be 0 if en_i is set to 1 (useful when oh_i can be masked).
  parameter bit          StrictCheck = 1,
  // This should only be disabled in special circumstances, for example
  // in non-comportable IPs where an error does not trigger an alert.
  parameter bit EnableAlertTriggerSVA = 1
) (
  // The module is combinational - the clock and reset are only used for assertions.
  input                          clk_i,
  input                          rst_ni,

  input  logic [OneHotWidth-1:0] oh_i,
  input  logic [AddrWidth-1:0]   addr_i,
  input  logic                   en_i,

  output logic                   err_o
);

  ///////////////////////
  // Binary tree logic //
  ///////////////////////

  `ASSERT_INIT(NumSources_A, OneHotWidth >= 1)
  `ASSERT_INIT(AddrWidth_A, AddrWidth >= 1)
  `ASSERT_INIT(AddrRange_A, OneHotWidth <= 2**AddrWidth)
  `ASSERT_INIT(AddrImpliesEnable_A, AddrCheck && EnableCheck || !AddrCheck)

  // Align to powers of 2 for simplicity.
  // A full binary tree with N levels has 2**N + 2**N-1 nodes.
  localparam int NumLevels = AddrWidth;
  logic [2**(NumLevels+1)-2:0] or_tree;
  logic [2**(NumLevels+1)-2:0] and_tree; // Used for the address check
  logic [2**(NumLevels+1)-2:0] err_tree; // Used for the enable check

  for (genvar level = 0; level < NumLevels+1; level++) begin : gen_tree
    //
    // level+1   C0   C1   <- "Base1" points to the first node on "level+1",
    //            \  /         these nodes are the children of the nodes one level below
    // level       Pa      <- "Base0", points to the first node on "level",
    //                         these nodes are the parents of the nodes one level above
    //
    // hence we have the following indices for the paPa, C0, C1 nodes:
    // Pa = 2**level     - 1 + offset       = Base0 + offset
    // C0 = 2**(level+1) - 1 + 2*offset     = Base1 + 2*offset
    // C1 = 2**(level+1) - 1 + 2*offset + 1 = Base1 + 2*offset + 1
    //
    localparam int Base0 = (2**level)-1;
    localparam int Base1 = (2**(level+1))-1;

    for (genvar offset = 0; offset < 2**level; offset++) begin : gen_level
      localparam int Pa = Base0 + offset;
      localparam int C0 = Base1 + 2*offset;
      localparam int C1 = Base1 + 2*offset + 1;

      // This assigns the input values, their corresponding IDs and valid signals to the tree leafs.
      if (level == NumLevels) begin : gen_leafs
        if (offset < OneHotWidth) begin : gen_assign
          assign or_tree[Pa]  = oh_i[offset];
          assign and_tree[Pa] = oh_i[offset];
        end else begin : gen_tie_off
          assign or_tree[Pa]  = 1'b0;
          assign and_tree[Pa] = 1'b0;
        end
        assign err_tree[Pa] = 1'b0;
      // This creates the node assignments.
      end else begin : gen_nodes
        assign or_tree[Pa]  = or_tree[C0] || or_tree[C1];
        assign and_tree[Pa] = (!addr_i[AddrWidth-1-level] && and_tree[C0]) ||
                              (addr_i[AddrWidth-1-level] && and_tree[C1]);
        assign err_tree[Pa] = (or_tree[C0] && or_tree[C1]) || err_tree[C0] || err_tree[C1];
      end
    end : gen_level
  end : gen_tree

  ///////////////////
  // Onehot Checks //
  ///////////////////

  logic enable_err, addr_err, oh0_err;
  assign err_o = oh0_err || enable_err || addr_err;

  // Check that no more than 1 bit is set in the vector.
  assign oh0_err = err_tree[0];
  `ASSERT(Onehot0Check_A, !$onehot0(oh_i) |-> err_o)

  // Check that en_i agrees with (|oh_i).
  // Note: if StrictCheck 0, the oh_i vector may be all-zero if en_i == 1 (but not vice versa).
  if (EnableCheck) begin : gen_enable_check
    if (StrictCheck) begin : gen_strict
      assign enable_err = or_tree[0] ^ en_i;
      `ASSERT(EnableCheck_A, (|oh_i) != en_i |-> err_o)
    end else begin : gen_not_strict
      assign enable_err = !en_i && or_tree[0];
      `ASSERT(EnableCheck_A, !en_i && (|oh_i) |-> err_o)
    end
  end else begin : gen_no_enable_check
    logic unused_or_tree;
    assign unused_or_tree = ^or_tree;
    assign enable_err = 1'b0;
  end

  // Check that the set bit is actually in the correct position.
  if (AddrCheck) begin : gen_addr_check_strict
    assign addr_err = or_tree[0] ^ and_tree[0];
    `ASSERT(AddrCheck_A, oh_i[addr_i] != (|oh_i) |-> err_o)
  end else begin : gen_no_addr_check_strict
    logic unused_and_tree;
    assign unused_and_tree = ^and_tree;
    assign addr_err = 1'b0;
  end

  // This logic that will be assign to one, when user adds macro
  // ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ALERT to check the error with alert, in case that
  // prim_onehot_check is used in design without adding this assertion check.
  `ifdef INC_ASSERT
  `ifndef PRIM_DEFAULT_IMPL
    `define PRIM_DEFAULT_IMPL prim_pkg::ImplGeneric
  `endif
  parameter prim_pkg::impl_e Impl = `PRIM_DEFAULT_IMPL;

  logic unused_assert_connected;
  // TODO(#13337): only check generic for now. The path of this prim in other Impl may differ
  if (Impl == prim_pkg::ImplGeneric) begin : gen_generic
    `ASSERT_INIT_NET(AssertConnected_A, unused_assert_connected === 1'b1 || !EnableAlertTriggerSVA)
  end
  `endif
endmodule : prim_onehot_check


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// This file is auto-generated.
// Used parser: Fallback (regex)


// This is to prevent AscentLint warnings in the generated
// abstract prim wrapper. These warnings occur due to the .*
// use. TODO: we may want to move these inline waivers
// into a separate, generated waiver file for consistency.
//ri lint_check_off OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ
module prim_flop_en

#(

  parameter int               Width      = 1,
  parameter bit               EnSecBuf   = 0,
  parameter logic [Width-1:0] ResetValue = 0

) (
  input                    clk_i,
  input                    rst_ni,
  input                    en_i,
  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_o
);

  if (1) begin : gen_generic
    prim_generic_flop_en #(
      .EnSecBuf(EnSecBuf),
      .ResetValue(ResetValue),
      .Width(Width)
    ) u_impl_generic (
      .*
    );

  end

endmodule
//ri lint_check_on OUTPUT_NOT_DRIVEN INPUT_NOT_READ HIER_BRANCH_NOT_READ


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Convenience module for wrapping prim_and2 for use in blanking.
// When en_i == 1 the input is fed through to the output.
// When en_i == 0 the output is 0.
module prim_blanker #(
  parameter int Width = 1
) (
  input  logic [Width-1:0] in_i,
  input  logic             en_i,
  output logic [Width-1:0] out_o
);
  prim_and2 #(.Width(Width)) u_blank_and (
    .in0_i(in_i),
    .in1_i({Width{en_i}}),
    .out_o
  );
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Hardened LFSR module that instantiates two LFSRs of the same type.
// The state vector of both LFSRs is constantly checked and an error is asserted if the
// two states are inconsistent.

module prim_double_lfsr #(
  // prim_lfsr parameters - refer to prim_lfsr for their meaning/
  parameter                    LfsrType     = "GAL_XOR",
  parameter int unsigned       LfsrDw       = 32,
  localparam int unsigned      LfsrIdxDw    = $clog2(LfsrDw),
  parameter int unsigned       EntropyDw    =  8,
  parameter int unsigned       StateOutDw   =  8,
  parameter logic [LfsrDw-1:0] DefaultSeed  = LfsrDw'(1),
  parameter logic [LfsrDw-1:0] CustomCoeffs = '0,
  parameter bit                StatePermEn  = 1'b0,
  parameter logic [LfsrDw-1:0][LfsrIdxDw-1:0] StatePerm = '0,
  parameter bit                MaxLenSVA    = 1'b1,
  parameter bit                LockupSVA    = 1'b1,
  parameter bit                ExtSeedSVA   = 1'b1,
  parameter bit                NonLinearOut = 1'b0,
  // This should only be disabled in special circumstances, for example
  // in non-comportable IPs where an error does not trigger an alert.
  parameter bit                EnableAlertTriggerSVA = 1
) (
  input                         clk_i,
  input                         rst_ni,
  input                         seed_en_i,
  input        [LfsrDw-1:0]     seed_i,
  input                         lfsr_en_i,
  input        [EntropyDw-1:0]  entropy_i,
  output logic [StateOutDw-1:0] state_o,
  // Asserted if the parallel LFSR states are inconsistent.
  output logic                  err_o
);


  logic [1:0][LfsrDw-1:0] lfsr_state;
  // We employ redundant LFSRs to guard against FI attacks.
  for (genvar k = 0; k < 2; k++) begin : gen_double_lfsr
    // Instantiate size_only buffers to prevent
    // optimization / merging of redundant logic.
    logic lfsr_en_buf, seed_en_buf;
    logic [EntropyDw-1:0] entropy_buf;
    logic [LfsrDw-1:0] seed_buf, lfsr_state_unbuf;
    prim_buf #(
      .Width(EntropyDw + LfsrDw + 2)
    ) u_prim_buf_input (
      .in_i({seed_en_i, seed_i, lfsr_en_i, entropy_i}),
      .out_o({seed_en_buf, seed_buf, lfsr_en_buf, entropy_buf})
    );

    prim_lfsr #(
      .LfsrType(LfsrType),
      .LfsrDw(LfsrDw),
      .EntropyDw(EntropyDw),
      // output the full width so that the states can be cross checked.
      .StateOutDw(LfsrDw),
      .DefaultSeed(DefaultSeed),
      .CustomCoeffs(CustomCoeffs),
      .StatePermEn(StatePermEn),
      .StatePerm(StatePerm),
      .MaxLenSVA(MaxLenSVA),
      .LockupSVA(LockupSVA),
      .ExtSeedSVA(ExtSeedSVA),
      .NonLinearOut(NonLinearOut)
    ) u_prim_lfsr (
      .clk_i,
      .rst_ni,
      .seed_en_i  ( seed_en_buf      ),
      .seed_i     ( seed_buf         ),
      .lfsr_en_i  ( lfsr_en_buf      ),
      .entropy_i  ( entropy_buf      ),
      .state_o    ( lfsr_state_unbuf )
    );

    prim_buf #(
      .Width(LfsrDw)
    ) u_prim_buf_output (
      .in_i(lfsr_state_unbuf),
      .out_o(lfsr_state[k])
    );
  end

`ifdef SIMULATION
`ifndef VERILATOR
  // Ensure both LFSRs start off with the same default seed. if randomized in simulations.
  initial begin : p_sync_lfsr_default_seed
    wait (!$isunknown(gen_double_lfsr[0].u_prim_lfsr.DefaultSeedLocal));
    wait (!$isunknown(gen_double_lfsr[1].u_prim_lfsr.DefaultSeedLocal));
    gen_double_lfsr[1].u_prim_lfsr.DefaultSeedLocal =
        gen_double_lfsr[0].u_prim_lfsr.DefaultSeedLocal;
    $display("%m: Updated gen_double_lfsr[1].u_prim_lfsr.DefaultSeedLocal = 0x%0h",
        gen_double_lfsr[1].u_prim_lfsr.DefaultSeedLocal);
  end
`endif
`endif

  // Output the state from the first LFSR
  assign state_o = lfsr_state[0][StateOutDw-1:0];
  assign err_o = lfsr_state[0] != lfsr_state[1];

  // This logic that will be assign to one, when user adds macro
  // ASSERT_PRIM_DOUBLE_LFSR_ERROR_TRIGGER_ALERT to check the error with alert, in case that
  // prim_double_lfsr is used in design without adding this assertion check.
  `ifdef INC_ASSERT
  logic unused_assert_connected;

  `ASSERT_INIT_NET(AssertConnected_A, unused_assert_connected === 1'b1 || !EnableAlertTriggerSVA)
  `endif
endmodule : prim_double_lfsr


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Generic double-synchronizer flop
// This may need to be moved to prim_generic if libraries have a specific cell
// for synchronization

module prim_flop_2sync #(
  parameter int               Width      = 16,
  parameter logic [Width-1:0] ResetValue = '0,
  parameter bit               EnablePrimCdcRand = 1
) (
  input                    clk_i,
  input                    rst_ni,
  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_o
);

  logic [Width-1:0] d_o;
  logic [Width-1:0] intq;

`ifdef SIMULATION

  prim_cdc_rand_delay #(
    .DataWidth(Width),
    .Enable(EnablePrimCdcRand)
  ) u_prim_cdc_rand_delay (
    .clk_i,
    .rst_ni,
    .src_data_i(d_i),
    .prev_data_i(intq),
    .dst_data_o(d_o)
  );
`else // !`ifdef SIMULATION
  logic unused_sig;
  assign unused_sig = EnablePrimCdcRand;
  always_comb d_o = d_i;
`endif // !`ifdef SIMULATION

  prim_flop #(
    .Width(Width),
    .ResetValue(ResetValue)
  ) u_sync_1 (
    .clk_i,
    .rst_ni,
    .d_i(d_o),
    .q_o(intq)
  );

  prim_flop #(
    .Width(Width),
    .ResetValue(ResetValue)
  ) u_sync_2 (
    .clk_i,
    .rst_ni,
    .d_i(intq),
    .q_o
  );

endmodule : prim_flop_2sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// This package defines common multibit signal types, active high and active low values and
// the corresponding functions to test whether the values are set or not.

`include "prim_assert.sv"

package prim_mubi_pkg;

  //////////////////////////////////////////////
  // 4 Bit Multibit Type and Functions //
  //////////////////////////////////////////////

  parameter int MuBi4Width = 4;
  typedef enum logic [MuBi4Width-1:0] {
    MuBi4True = 4'h6, // enabled
    MuBi4False = 4'h9  // disabled
  } mubi4_t;

  // This is a prerequisite for the multibit functions below to work.
  `ASSERT_STATIC_IN_PACKAGE(CheckMuBi4ValsComplementary_A, MuBi4True == ~MuBi4False)

  // Test whether the value is supplied is one of the valid enumerations
  function automatic logic mubi4_test_invalid(mubi4_t val);
    return ~(val inside {MuBi4True, MuBi4False});
  endfunction : mubi4_test_invalid

  // Convert a 1 input value to a mubi output
  function automatic mubi4_t mubi4_bool_to_mubi(logic val);
    return (val ? MuBi4True : MuBi4False);
  endfunction : mubi4_bool_to_mubi

  // Test whether the multibit value signals an "enabled" condition.
  // The strict version of this function requires
  // the multibit value to equal True.
  function automatic logic mubi4_test_true_strict(mubi4_t val);
    return MuBi4True == val;
  endfunction : mubi4_test_true_strict

  // Test whether the multibit value signals a "disabled" condition.
  // The strict version of this function requires
  // the multibit value to equal False.
  function automatic logic mubi4_test_false_strict(mubi4_t val);
    return MuBi4False == val;
  endfunction : mubi4_test_false_strict

  // Test whether the multibit value signals an "enabled" condition.
  // The loose version of this function interprets all
  // values other than False as "enabled".
  function automatic logic mubi4_test_true_loose(mubi4_t val);
    return MuBi4False != val;
  endfunction : mubi4_test_true_loose

  // Test whether the multibit value signals a "disabled" condition.
  // The loose version of this function interprets all
  // values other than True as "disabled".
  function automatic logic mubi4_test_false_loose(mubi4_t val);
    return MuBi4True != val;
  endfunction : mubi4_test_false_loose


  // Performs a logical OR operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | act
  // !act | act  | act
  // act  | act  | act
  //
  function automatic mubi4_t mubi4_or(mubi4_t a, mubi4_t b, mubi4_t act);
    logic [MuBi4Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi4Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] || b_in[k];
      end else begin
        out[k] = a_in[k] && b_in[k];
      end
    end
    return mubi4_t'(out);
  endfunction : mubi4_or

  // Performs a logical AND operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | !act
  // !act | act  | !act
  // act  | act  | act
  //
  function automatic mubi4_t mubi4_and(mubi4_t a, mubi4_t b, mubi4_t act);
    logic [MuBi4Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi4Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] && b_in[k];
      end else begin
        out[k] = a_in[k] || b_in[k];
      end
    end
    return mubi4_t'(out);
  endfunction : mubi4_and

  // Performs a logical OR operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi4_t mubi4_or_hi(mubi4_t a, mubi4_t b);
    return mubi4_or(a, b, MuBi4True);
  endfunction : mubi4_or_hi

  // Performs a logical AND operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi4_t mubi4_and_hi(mubi4_t a, mubi4_t b);
    return mubi4_and(a, b, MuBi4True);
  endfunction : mubi4_and_hi

  // Performs a logical OR operation between two multibit values.
  // This treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi4_t mubi4_or_lo(mubi4_t a, mubi4_t b);
    return mubi4_or(a, b, MuBi4False);
  endfunction : mubi4_or_lo

  // Performs a logical AND operation between two multibit values.
  // Tlos treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi4_t mubi4_and_lo(mubi4_t a, mubi4_t b);
    return mubi4_and(a, b, MuBi4False);
  endfunction : mubi4_and_lo

  //////////////////////////////////////////////
  // 8 Bit Multibit Type and Functions //
  //////////////////////////////////////////////

  parameter int MuBi8Width = 8;
  typedef enum logic [MuBi8Width-1:0] {
    MuBi8True = 8'h96, // enabled
    MuBi8False = 8'h69  // disabled
  } mubi8_t;

  // This is a prerequisite for the multibit functions below to work.
  `ASSERT_STATIC_IN_PACKAGE(CheckMuBi8ValsComplementary_A, MuBi8True == ~MuBi8False)

  // Test whether the value is supplied is one of the valid enumerations
  function automatic logic mubi8_test_invalid(mubi8_t val);
    return ~(val inside {MuBi8True, MuBi8False});
  endfunction : mubi8_test_invalid

  // Convert a 1 input value to a mubi output
  function automatic mubi8_t mubi8_bool_to_mubi(logic val);
    return (val ? MuBi8True : MuBi8False);
  endfunction : mubi8_bool_to_mubi

  // Test whether the multibit value signals an "enabled" condition.
  // The strict version of this function requires
  // the multibit value to equal True.
  function automatic logic mubi8_test_true_strict(mubi8_t val);
    return MuBi8True == val;
  endfunction : mubi8_test_true_strict

  // Test whether the multibit value signals a "disabled" condition.
  // The strict version of this function requires
  // the multibit value to equal False.
  function automatic logic mubi8_test_false_strict(mubi8_t val);
    return MuBi8False == val;
  endfunction : mubi8_test_false_strict

  // Test whether the multibit value signals an "enabled" condition.
  // The loose version of this function interprets all
  // values other than False as "enabled".
  function automatic logic mubi8_test_true_loose(mubi8_t val);
    return MuBi8False != val;
  endfunction : mubi8_test_true_loose

  // Test whether the multibit value signals a "disabled" condition.
  // The loose version of this function interprets all
  // values other than True as "disabled".
  function automatic logic mubi8_test_false_loose(mubi8_t val);
    return MuBi8True != val;
  endfunction : mubi8_test_false_loose


  // Performs a logical OR operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | act
  // !act | act  | act
  // act  | act  | act
  //
  function automatic mubi8_t mubi8_or(mubi8_t a, mubi8_t b, mubi8_t act);
    logic [MuBi8Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi8Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] || b_in[k];
      end else begin
        out[k] = a_in[k] && b_in[k];
      end
    end
    return mubi8_t'(out);
  endfunction : mubi8_or

  // Performs a logical AND operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | !act
  // !act | act  | !act
  // act  | act  | act
  //
  function automatic mubi8_t mubi8_and(mubi8_t a, mubi8_t b, mubi8_t act);
    logic [MuBi8Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi8Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] && b_in[k];
      end else begin
        out[k] = a_in[k] || b_in[k];
      end
    end
    return mubi8_t'(out);
  endfunction : mubi8_and

  // Performs a logical OR operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi8_t mubi8_or_hi(mubi8_t a, mubi8_t b);
    return mubi8_or(a, b, MuBi8True);
  endfunction : mubi8_or_hi

  // Performs a logical AND operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi8_t mubi8_and_hi(mubi8_t a, mubi8_t b);
    return mubi8_and(a, b, MuBi8True);
  endfunction : mubi8_and_hi

  // Performs a logical OR operation between two multibit values.
  // This treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi8_t mubi8_or_lo(mubi8_t a, mubi8_t b);
    return mubi8_or(a, b, MuBi8False);
  endfunction : mubi8_or_lo

  // Performs a logical AND operation between two multibit values.
  // Tlos treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi8_t mubi8_and_lo(mubi8_t a, mubi8_t b);
    return mubi8_and(a, b, MuBi8False);
  endfunction : mubi8_and_lo

  //////////////////////////////////////////////
  // 12 Bit Multibit Type and Functions //
  //////////////////////////////////////////////

  parameter int MuBi12Width = 12;
  typedef enum logic [MuBi12Width-1:0] {
    MuBi12True = 12'h696, // enabled
    MuBi12False = 12'h969  // disabled
  } mubi12_t;

  // This is a prerequisite for the multibit functions below to work.
  `ASSERT_STATIC_IN_PACKAGE(CheckMuBi12ValsComplementary_A, MuBi12True == ~MuBi12False)

  // Test whether the value is supplied is one of the valid enumerations
  function automatic logic mubi12_test_invalid(mubi12_t val);
    return ~(val inside {MuBi12True, MuBi12False});
  endfunction : mubi12_test_invalid

  // Convert a 1 input value to a mubi output
  function automatic mubi12_t mubi12_bool_to_mubi(logic val);
    return (val ? MuBi12True : MuBi12False);
  endfunction : mubi12_bool_to_mubi

  // Test whether the multibit value signals an "enabled" condition.
  // The strict version of this function requires
  // the multibit value to equal True.
  function automatic logic mubi12_test_true_strict(mubi12_t val);
    return MuBi12True == val;
  endfunction : mubi12_test_true_strict

  // Test whether the multibit value signals a "disabled" condition.
  // The strict version of this function requires
  // the multibit value to equal False.
  function automatic logic mubi12_test_false_strict(mubi12_t val);
    return MuBi12False == val;
  endfunction : mubi12_test_false_strict

  // Test whether the multibit value signals an "enabled" condition.
  // The loose version of this function interprets all
  // values other than False as "enabled".
  function automatic logic mubi12_test_true_loose(mubi12_t val);
    return MuBi12False != val;
  endfunction : mubi12_test_true_loose

  // Test whether the multibit value signals a "disabled" condition.
  // The loose version of this function interprets all
  // values other than True as "disabled".
  function automatic logic mubi12_test_false_loose(mubi12_t val);
    return MuBi12True != val;
  endfunction : mubi12_test_false_loose


  // Performs a logical OR operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | act
  // !act | act  | act
  // act  | act  | act
  //
  function automatic mubi12_t mubi12_or(mubi12_t a, mubi12_t b, mubi12_t act);
    logic [MuBi12Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi12Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] || b_in[k];
      end else begin
        out[k] = a_in[k] && b_in[k];
      end
    end
    return mubi12_t'(out);
  endfunction : mubi12_or

  // Performs a logical AND operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | !act
  // !act | act  | !act
  // act  | act  | act
  //
  function automatic mubi12_t mubi12_and(mubi12_t a, mubi12_t b, mubi12_t act);
    logic [MuBi12Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi12Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] && b_in[k];
      end else begin
        out[k] = a_in[k] || b_in[k];
      end
    end
    return mubi12_t'(out);
  endfunction : mubi12_and

  // Performs a logical OR operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi12_t mubi12_or_hi(mubi12_t a, mubi12_t b);
    return mubi12_or(a, b, MuBi12True);
  endfunction : mubi12_or_hi

  // Performs a logical AND operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi12_t mubi12_and_hi(mubi12_t a, mubi12_t b);
    return mubi12_and(a, b, MuBi12True);
  endfunction : mubi12_and_hi

  // Performs a logical OR operation between two multibit values.
  // This treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi12_t mubi12_or_lo(mubi12_t a, mubi12_t b);
    return mubi12_or(a, b, MuBi12False);
  endfunction : mubi12_or_lo

  // Performs a logical AND operation between two multibit values.
  // Tlos treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi12_t mubi12_and_lo(mubi12_t a, mubi12_t b);
    return mubi12_and(a, b, MuBi12False);
  endfunction : mubi12_and_lo

  //////////////////////////////////////////////
  // 16 Bit Multibit Type and Functions //
  //////////////////////////////////////////////

  parameter int MuBi16Width = 16;
  typedef enum logic [MuBi16Width-1:0] {
    MuBi16True = 16'h9696, // enabled
    MuBi16False = 16'h6969  // disabled
  } mubi16_t;

  // This is a prerequisite for the multibit functions below to work.
  `ASSERT_STATIC_IN_PACKAGE(CheckMuBi16ValsComplementary_A, MuBi16True == ~MuBi16False)

  // Test whether the value is supplied is one of the valid enumerations
  function automatic logic mubi16_test_invalid(mubi16_t val);
    return ~(val inside {MuBi16True, MuBi16False});
  endfunction : mubi16_test_invalid

  // Convert a 1 input value to a mubi output
  function automatic mubi16_t mubi16_bool_to_mubi(logic val);
    return (val ? MuBi16True : MuBi16False);
  endfunction : mubi16_bool_to_mubi

  // Test whether the multibit value signals an "enabled" condition.
  // The strict version of this function requires
  // the multibit value to equal True.
  function automatic logic mubi16_test_true_strict(mubi16_t val);
    return MuBi16True == val;
  endfunction : mubi16_test_true_strict

  // Test whether the multibit value signals a "disabled" condition.
  // The strict version of this function requires
  // the multibit value to equal False.
  function automatic logic mubi16_test_false_strict(mubi16_t val);
    return MuBi16False == val;
  endfunction : mubi16_test_false_strict

  // Test whether the multibit value signals an "enabled" condition.
  // The loose version of this function interprets all
  // values other than False as "enabled".
  function automatic logic mubi16_test_true_loose(mubi16_t val);
    return MuBi16False != val;
  endfunction : mubi16_test_true_loose

  // Test whether the multibit value signals a "disabled" condition.
  // The loose version of this function interprets all
  // values other than True as "disabled".
  function automatic logic mubi16_test_false_loose(mubi16_t val);
    return MuBi16True != val;
  endfunction : mubi16_test_false_loose


  // Performs a logical OR operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | act
  // !act | act  | act
  // act  | act  | act
  //
  function automatic mubi16_t mubi16_or(mubi16_t a, mubi16_t b, mubi16_t act);
    logic [MuBi16Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi16Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] || b_in[k];
      end else begin
        out[k] = a_in[k] && b_in[k];
      end
    end
    return mubi16_t'(out);
  endfunction : mubi16_or

  // Performs a logical AND operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | !act
  // !act | act  | !act
  // act  | act  | act
  //
  function automatic mubi16_t mubi16_and(mubi16_t a, mubi16_t b, mubi16_t act);
    logic [MuBi16Width-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < MuBi16Width; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] && b_in[k];
      end else begin
        out[k] = a_in[k] || b_in[k];
      end
    end
    return mubi16_t'(out);
  endfunction : mubi16_and

  // Performs a logical OR operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi16_t mubi16_or_hi(mubi16_t a, mubi16_t b);
    return mubi16_or(a, b, MuBi16True);
  endfunction : mubi16_or_hi

  // Performs a logical AND operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi16_t mubi16_and_hi(mubi16_t a, mubi16_t b);
    return mubi16_and(a, b, MuBi16True);
  endfunction : mubi16_and_hi

  // Performs a logical OR operation between two multibit values.
  // This treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi16_t mubi16_or_lo(mubi16_t a, mubi16_t b);
    return mubi16_or(a, b, MuBi16False);
  endfunction : mubi16_or_lo

  // Performs a logical AND operation between two multibit values.
  // Tlos treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic mubi16_t mubi16_and_lo(mubi16_t a, mubi16_t b);
    return mubi16_and(a, b, MuBi16False);
  endfunction : mubi16_and_lo

endpackage : prim_mubi_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Multibit sender module. This module is instantiates a hand-picked flop cell for each bit in the
// multibit signal such that tools do not optimize the multibit encoding.

`include "prim_assert.sv"

module prim_mubi4_sender
  import prim_mubi_pkg::*;
#(
  // This flops the output if set to 1.
  // In special cases where the sender is in the same clock domain as the receiver,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // Enable anchor buffer
  parameter bit EnSecBuf = 0,
  // Reset value for the sender flops
  parameter mubi4_t ResetValue = MuBi4False
) (
  input          clk_i,
  input          rst_ni,
  input  mubi4_t mubi_i,
  output mubi4_t mubi_o
);

  logic [MuBi4Width-1:0] mubi, mubi_int, mubi_out;
  assign mubi = MuBi4Width'(mubi_i);

  // first generation block decides whether a flop should be present
  if (AsyncOn) begin : gen_flops
    prim_flop #(
      .Width(MuBi4Width),
      .ResetValue(MuBi4Width'(ResetValue))
    ) u_prim_flop (
      .clk_i,
      .rst_ni,
      .d_i   ( mubi     ),
      .q_o   ( mubi_int )
    );
  end else begin : gen_no_flops
    assign mubi_int = mubi;

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for sythesis since it is unloaded.
    mubi4_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi4False;
      end else begin
         unused_logic <= mubi_i;
      end
    end
  end

  // second generation block determines output buffer type
  // 1. If EnSecBuf -> always leads to a sec buffer regardless of first block
  // 2. If not EnSecBuf and not AsyncOn -> use normal buffer
  // 3. If not EnSecBuf and AsyncOn -> feed through
  if (EnSecBuf) begin : gen_sec_buf
    prim_sec_anchor_buf #(
      .Width(4)
    ) u_prim_sec_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else if (!AsyncOn) begin : gen_prim_buf
    prim_buf #(
      .Width(4)
    ) u_prim_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else begin : gen_feedthru
    assign mubi_out = mubi_int;
  end

  assign mubi_o = mubi4_t'(mubi_out);

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi4_sender


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Double-synchronizer flop for multibit signals with additional output buffers.

`include "prim_assert.sv"

module prim_mubi4_sync
  import prim_mubi_pkg::*;
#(
  // Number of separately buffered output signals.
  // The buffer cells have a don't touch constraint
  // on them such that synthesis tools won't collapse
  // all copies into one signal.
  parameter int NumCopies = 1,
  // This instantiates the synchronizer flops if set to 1.
  // In special cases where the receiver is in the same clock domain as the sender,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // This controls whether the mubi module institutes stability checks when
  // AsyncOn is set.  If stability checks are on, a 3rd stage of storage is
  // added after the synchronizers and the outputs only updated if the 3rd
  // stage and sychronizer agree.  If they do not agree, the ResetValue is
  // output instead.
  parameter bit StabilityCheck = 0,
  // Reset value for the sync flops
  parameter mubi4_t ResetValue = MuBi4False
) (
  input                          clk_i,
  input                          rst_ni,
  input  mubi4_t                 mubi_i,
  output mubi4_t [NumCopies-1:0] mubi_o
);

  `ASSERT_INIT(NumCopiesMustBeGreaterZero_A, NumCopies > 0)

  logic [MuBi4Width-1:0] mubi;
  if (AsyncOn) begin : gen_flops
    logic [MuBi4Width-1:0] mubi_sync;
    prim_flop_2sync #(
      .Width(MuBi4Width),
      .ResetValue(MuBi4Width'(ResetValue))
    ) u_prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(MuBi4Width'(mubi_i)),
      .q_o(mubi_sync)
    );

    if (StabilityCheck) begin : gen_stable_chks
      logic [MuBi4Width-1:0] mubi_q;
      prim_flop #(
        .Width(MuBi4Width),
        .ResetValue(MuBi4Width'(ResetValue))
      ) u_prim_flop_3rd_stage (
        .clk_i,
        .rst_ni,
        .d_i(mubi_sync),
        .q_o(mubi_q)
      );

      logic [MuBi4Width-1:0] sig_unstable;
      prim_xor2 #(
        .Width(MuBi4Width)
      ) u_mubi_xor (
        .in0_i(mubi_sync),
        .in1_i(mubi_q),
        .out_o(sig_unstable)
      );

      logic [MuBi4Width-1:0] reset_value;
      assign reset_value = ResetValue;

      for (genvar k = 0; k < MuBi4Width; k++) begin : gen_bufs_muxes
        logic [MuBi4Width-1:0] sig_unstable_buf;

        // each mux gets its own buffered output, this ensures the OR-ing
        // cannot be defeated in one place.
        prim_sec_anchor_buf #(
          .Width(MuBi4Width)
        ) u_sig_unstable_buf (
          .in_i(sig_unstable),
          .out_o(sig_unstable_buf)
        );

        // if any xor indicates signal is unstable, output the reset
        // value. note that the input and output signals of this mux
        // are driven/read by constrained primitive cells (regs, buffers),
        // hence this mux can be implemented behaviorally.
        assign mubi[k] = (|sig_unstable_buf) ? reset_value[k] : mubi_q[k];
      end

// Note regarding SVAs below:
//
// 1) Without the sampled rst_ni pre-condition, this may cause false assertion failures right after
// a reset release, since the "disable iff" condition with the rst_ni is sampled in the "observed"
// SV scheduler region after all assignments have been evaluated (see also LRM section 16.12, page
// 423). This is a simulation artifact due to reset synchronization in RTL, which releases rst_ni
// on the active clock edge. This causes the assertion to evaluate although the reset was actually
// 0 when entering this simulation cycle.
//
// 2) Similarly to 1) there can be sampling mismatches of the lc_en_i signal since that signal may
// originate from a different clock domain. I.e., in cases where the lc_en_i signal changes exactly
// at the same time that the clk_i signal rises, the SVA will not pick up that change in that clock
// cycle, whereas RTL will because SVAs sample values in the "preponed" region. To that end we make
// use of an RTL helper variable to sample the lc_en_i signal, hence ensuring that there are no
// sampling mismatches.
`ifdef INC_ASSERT
      mubi4_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputIfUnstable_A, sig_unstable |-> mubi_o == {NumCopies{reset_value}})
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##[3:4] sig_unstable || mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}})
`endif
    end else begin : gen_no_stable_chks
      assign mubi = mubi_sync;
`ifdef INC_ASSERT
      mubi4_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##3 (mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}} ||
                              $past(mubi_in_sva_q, 2) != $past(mubi_in_sva_q, 1)))
`endif
    end
  end else begin : gen_no_flops

    //VCS coverage off
    // pragma coverage off

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for synthesis since it is unloaded.
    mubi4_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi4False;
      end else begin
         unused_logic <= mubi_i;
      end
    end

    //VCS coverage on
    // pragma coverage on

    assign mubi = MuBi4Width'(mubi_i);

    `ASSERT(OutputDelay_A, mubi_o == {NumCopies{mubi_i}})
  end

  for (genvar j = 0; j < NumCopies; j++) begin : gen_buffs
    logic [MuBi4Width-1:0] mubi_out;
    for (genvar k = 0; k < MuBi4Width; k++) begin : gen_bits
      prim_buf u_prim_buf (
        .in_i(mubi[k]),
        .out_o(mubi_out[k])
      );
    end
    assign mubi_o[j] = mubi4_t'(mubi_out);
  end

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi4_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Decoder for multibit control signals with additional input buffers.

`include "prim_assert.sv"

module prim_mubi4_dec
  import prim_mubi_pkg::*;
#(
  parameter bit TestTrue = 1,
  parameter bit TestStrict = 1
) (
  input  mubi4_t mubi_i,
  output logic           mubi_dec_o
);

logic [MuBi4Width-1:0] mubi, mubi_out;
assign mubi = MuBi4Width'(mubi_i);

// The buffer cells have a don't touch constraint on them
// such that synthesis tools won't collapse them
for (genvar k = 0; k < MuBi4Width; k++) begin : gen_bits
  prim_buf u_prim_buf (
    .in_i  ( mubi[k]     ),
    .out_o ( mubi_out[k] )
  );
end

if (TestTrue && TestStrict) begin : gen_test_true_strict
  assign mubi_dec_o = mubi4_test_true_strict(mubi4_t'(mubi_out));
end else if (TestTrue && !TestStrict) begin : gen_test_true_loose
  assign mubi_dec_o = mubi4_test_true_loose(mubi4_t'(mubi_out));
end else if (!TestTrue && TestStrict) begin : gen_test_false_strict
  assign mubi_dec_o = mubi4_test_false_strict(mubi4_t'(mubi_out));
end else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
  assign mubi_dec_o = mubi4_test_false_loose(mubi4_t'(mubi_out));
end else begin : gen_unknown_config
  `ASSERT_INIT(UnknownConfig_A, 0)
end

endmodule : prim_mubi4_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Multibit sender module. This module is instantiates a hand-picked flop cell for each bit in the
// multibit signal such that tools do not optimize the multibit encoding.

`include "prim_assert.sv"

module prim_mubi8_sender
  import prim_mubi_pkg::*;
#(
  // This flops the output if set to 1.
  // In special cases where the sender is in the same clock domain as the receiver,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // Enable anchor buffer
  parameter bit EnSecBuf = 0,
  // Reset value for the sender flops
  parameter mubi8_t ResetValue = MuBi8False
) (
  input          clk_i,
  input          rst_ni,
  input  mubi8_t mubi_i,
  output mubi8_t mubi_o
);

  logic [MuBi8Width-1:0] mubi, mubi_int, mubi_out;
  assign mubi = MuBi8Width'(mubi_i);

  // first generation block decides whether a flop should be present
  if (AsyncOn) begin : gen_flops
    prim_flop #(
      .Width(MuBi8Width),
      .ResetValue(MuBi8Width'(ResetValue))
    ) u_prim_flop (
      .clk_i,
      .rst_ni,
      .d_i   ( mubi     ),
      .q_o   ( mubi_int )
    );
  end else begin : gen_no_flops
    assign mubi_int = mubi;

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for sythesis since it is unloaded.
    mubi8_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi8False;
      end else begin
         unused_logic <= mubi_i;
      end
    end
  end

  // second generation block determines output buffer type
  // 1. If EnSecBuf -> always leads to a sec buffer regardless of first block
  // 2. If not EnSecBuf and not AsyncOn -> use normal buffer
  // 3. If not EnSecBuf and AsyncOn -> feed through
  if (EnSecBuf) begin : gen_sec_buf
    prim_sec_anchor_buf #(
      .Width(8)
    ) u_prim_sec_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else if (!AsyncOn) begin : gen_prim_buf
    prim_buf #(
      .Width(8)
    ) u_prim_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else begin : gen_feedthru
    assign mubi_out = mubi_int;
  end

  assign mubi_o = mubi8_t'(mubi_out);

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi8_sender


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Double-synchronizer flop for multibit signals with additional output buffers.

`include "prim_assert.sv"

module prim_mubi8_sync
  import prim_mubi_pkg::*;
#(
  // Number of separately buffered output signals.
  // The buffer cells have a don't touch constraint
  // on them such that synthesis tools won't collapse
  // all copies into one signal.
  parameter int NumCopies = 1,
  // This instantiates the synchronizer flops if set to 1.
  // In special cases where the receiver is in the same clock domain as the sender,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // This controls whether the mubi module institutes stability checks when
  // AsyncOn is set.  If stability checks are on, a 3rd stage of storage is
  // added after the synchronizers and the outputs only updated if the 3rd
  // stage and sychronizer agree.  If they do not agree, the ResetValue is
  // output instead.
  parameter bit StabilityCheck = 0,
  // Reset value for the sync flops
  parameter mubi8_t ResetValue = MuBi8False
) (
  input                          clk_i,
  input                          rst_ni,
  input  mubi8_t                 mubi_i,
  output mubi8_t [NumCopies-1:0] mubi_o
);

  `ASSERT_INIT(NumCopiesMustBeGreaterZero_A, NumCopies > 0)

  logic [MuBi8Width-1:0] mubi;
  if (AsyncOn) begin : gen_flops
    logic [MuBi8Width-1:0] mubi_sync;
    prim_flop_2sync #(
      .Width(MuBi8Width),
      .ResetValue(MuBi8Width'(ResetValue))
    ) u_prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(MuBi8Width'(mubi_i)),
      .q_o(mubi_sync)
    );

    if (StabilityCheck) begin : gen_stable_chks
      logic [MuBi8Width-1:0] mubi_q;
      prim_flop #(
        .Width(MuBi8Width),
        .ResetValue(MuBi8Width'(ResetValue))
      ) u_prim_flop_3rd_stage (
        .clk_i,
        .rst_ni,
        .d_i(mubi_sync),
        .q_o(mubi_q)
      );

      logic [MuBi8Width-1:0] sig_unstable;
      prim_xor2 #(
        .Width(MuBi8Width)
      ) u_mubi_xor (
        .in0_i(mubi_sync),
        .in1_i(mubi_q),
        .out_o(sig_unstable)
      );

      logic [MuBi8Width-1:0] reset_value;
      assign reset_value = ResetValue;

      for (genvar k = 0; k < MuBi8Width; k++) begin : gen_bufs_muxes
        logic [MuBi8Width-1:0] sig_unstable_buf;

        // each mux gets its own buffered output, this ensures the OR-ing
        // cannot be defeated in one place.
        prim_sec_anchor_buf #(
          .Width(MuBi8Width)
        ) u_sig_unstable_buf (
          .in_i(sig_unstable),
          .out_o(sig_unstable_buf)
        );

        // if any xor indicates signal is unstable, output the reset
        // value. note that the input and output signals of this mux
        // are driven/read by constrained primitive cells (regs, buffers),
        // hence this mux can be implemented behaviorally.
        assign mubi[k] = (|sig_unstable_buf) ? reset_value[k] : mubi_q[k];
      end

// Note regarding SVAs below:
//
// 1) Without the sampled rst_ni pre-condition, this may cause false assertion failures right after
// a reset release, since the "disable iff" condition with the rst_ni is sampled in the "observed"
// SV scheduler region after all assignments have been evaluated (see also LRM section 16.12, page
// 423). This is a simulation artifact due to reset synchronization in RTL, which releases rst_ni
// on the active clock edge. This causes the assertion to evaluate although the reset was actually
// 0 when entering this simulation cycle.
//
// 2) Similarly to 1) there can be sampling mismatches of the lc_en_i signal since that signal may
// originate from a different clock domain. I.e., in cases where the lc_en_i signal changes exactly
// at the same time that the clk_i signal rises, the SVA will not pick up that change in that clock
// cycle, whereas RTL will because SVAs sample values in the "preponed" region. To that end we make
// use of an RTL helper variable to sample the lc_en_i signal, hence ensuring that there are no
// sampling mismatches.
`ifdef INC_ASSERT
      mubi8_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputIfUnstable_A, sig_unstable |-> mubi_o == {NumCopies{reset_value}})
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##[3:4] sig_unstable || mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}})
`endif
    end else begin : gen_no_stable_chks
      assign mubi = mubi_sync;
`ifdef INC_ASSERT
      mubi8_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##3 (mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}} ||
                              $past(mubi_in_sva_q, 2) != $past(mubi_in_sva_q, 1)))
`endif
    end
  end else begin : gen_no_flops

    //VCS coverage off
    // pragma coverage off

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for synthesis since it is unloaded.
    mubi8_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi8False;
      end else begin
         unused_logic <= mubi_i;
      end
    end

    //VCS coverage on
    // pragma coverage on

    assign mubi = MuBi8Width'(mubi_i);

    `ASSERT(OutputDelay_A, mubi_o == {NumCopies{mubi_i}})
  end

  for (genvar j = 0; j < NumCopies; j++) begin : gen_buffs
    logic [MuBi8Width-1:0] mubi_out;
    for (genvar k = 0; k < MuBi8Width; k++) begin : gen_bits
      prim_buf u_prim_buf (
        .in_i(mubi[k]),
        .out_o(mubi_out[k])
      );
    end
    assign mubi_o[j] = mubi8_t'(mubi_out);
  end

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi8_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Decoder for multibit control signals with additional input buffers.

`include "prim_assert.sv"

module prim_mubi8_dec
  import prim_mubi_pkg::*;
#(
  parameter bit TestTrue = 1,
  parameter bit TestStrict = 1
) (
  input  mubi8_t mubi_i,
  output logic           mubi_dec_o
);

logic [MuBi8Width-1:0] mubi, mubi_out;
assign mubi = MuBi8Width'(mubi_i);

// The buffer cells have a don't touch constraint on them
// such that synthesis tools won't collapse them
for (genvar k = 0; k < MuBi8Width; k++) begin : gen_bits
  prim_buf u_prim_buf (
    .in_i  ( mubi[k]     ),
    .out_o ( mubi_out[k] )
  );
end

if (TestTrue && TestStrict) begin : gen_test_true_strict
  assign mubi_dec_o = mubi8_test_true_strict(mubi8_t'(mubi_out));
end else if (TestTrue && !TestStrict) begin : gen_test_true_loose
  assign mubi_dec_o = mubi8_test_true_loose(mubi8_t'(mubi_out));
end else if (!TestTrue && TestStrict) begin : gen_test_false_strict
  assign mubi_dec_o = mubi8_test_false_strict(mubi8_t'(mubi_out));
end else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
  assign mubi_dec_o = mubi8_test_false_loose(mubi8_t'(mubi_out));
end else begin : gen_unknown_config
  `ASSERT_INIT(UnknownConfig_A, 0)
end

endmodule : prim_mubi8_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Multibit sender module. This module is instantiates a hand-picked flop cell for each bit in the
// multibit signal such that tools do not optimize the multibit encoding.

`include "prim_assert.sv"

module prim_mubi12_sender
  import prim_mubi_pkg::*;
#(
  // This flops the output if set to 1.
  // In special cases where the sender is in the same clock domain as the receiver,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // Enable anchor buffer
  parameter bit EnSecBuf = 0,
  // Reset value for the sender flops
  parameter mubi12_t ResetValue = MuBi12False
) (
  input          clk_i,
  input          rst_ni,
  input  mubi12_t mubi_i,
  output mubi12_t mubi_o
);

  logic [MuBi12Width-1:0] mubi, mubi_int, mubi_out;
  assign mubi = MuBi12Width'(mubi_i);

  // first generation block decides whether a flop should be present
  if (AsyncOn) begin : gen_flops
    prim_flop #(
      .Width(MuBi12Width),
      .ResetValue(MuBi12Width'(ResetValue))
    ) u_prim_flop (
      .clk_i,
      .rst_ni,
      .d_i   ( mubi     ),
      .q_o   ( mubi_int )
    );
  end else begin : gen_no_flops
    assign mubi_int = mubi;

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for sythesis since it is unloaded.
    mubi12_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi12False;
      end else begin
         unused_logic <= mubi_i;
      end
    end
  end

  // second generation block determines output buffer type
  // 1. If EnSecBuf -> always leads to a sec buffer regardless of first block
  // 2. If not EnSecBuf and not AsyncOn -> use normal buffer
  // 3. If not EnSecBuf and AsyncOn -> feed through
  if (EnSecBuf) begin : gen_sec_buf
    prim_sec_anchor_buf #(
      .Width(12)
    ) u_prim_sec_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else if (!AsyncOn) begin : gen_prim_buf
    prim_buf #(
      .Width(12)
    ) u_prim_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else begin : gen_feedthru
    assign mubi_out = mubi_int;
  end

  assign mubi_o = mubi12_t'(mubi_out);

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi12_sender


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Double-synchronizer flop for multibit signals with additional output buffers.

`include "prim_assert.sv"

module prim_mubi12_sync
  import prim_mubi_pkg::*;
#(
  // Number of separately buffered output signals.
  // The buffer cells have a don't touch constraint
  // on them such that synthesis tools won't collapse
  // all copies into one signal.
  parameter int NumCopies = 1,
  // This instantiates the synchronizer flops if set to 1.
  // In special cases where the receiver is in the same clock domain as the sender,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // This controls whether the mubi module institutes stability checks when
  // AsyncOn is set.  If stability checks are on, a 3rd stage of storage is
  // added after the synchronizers and the outputs only updated if the 3rd
  // stage and sychronizer agree.  If they do not agree, the ResetValue is
  // output instead.
  parameter bit StabilityCheck = 0,
  // Reset value for the sync flops
  parameter mubi12_t ResetValue = MuBi12False
) (
  input                          clk_i,
  input                          rst_ni,
  input  mubi12_t                 mubi_i,
  output mubi12_t [NumCopies-1:0] mubi_o
);

  `ASSERT_INIT(NumCopiesMustBeGreaterZero_A, NumCopies > 0)

  logic [MuBi12Width-1:0] mubi;
  if (AsyncOn) begin : gen_flops
    logic [MuBi12Width-1:0] mubi_sync;
    prim_flop_2sync #(
      .Width(MuBi12Width),
      .ResetValue(MuBi12Width'(ResetValue))
    ) u_prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(MuBi12Width'(mubi_i)),
      .q_o(mubi_sync)
    );

    if (StabilityCheck) begin : gen_stable_chks
      logic [MuBi12Width-1:0] mubi_q;
      prim_flop #(
        .Width(MuBi12Width),
        .ResetValue(MuBi12Width'(ResetValue))
      ) u_prim_flop_3rd_stage (
        .clk_i,
        .rst_ni,
        .d_i(mubi_sync),
        .q_o(mubi_q)
      );

      logic [MuBi12Width-1:0] sig_unstable;
      prim_xor2 #(
        .Width(MuBi12Width)
      ) u_mubi_xor (
        .in0_i(mubi_sync),
        .in1_i(mubi_q),
        .out_o(sig_unstable)
      );

      logic [MuBi12Width-1:0] reset_value;
      assign reset_value = ResetValue;

      for (genvar k = 0; k < MuBi12Width; k++) begin : gen_bufs_muxes
        logic [MuBi12Width-1:0] sig_unstable_buf;

        // each mux gets its own buffered output, this ensures the OR-ing
        // cannot be defeated in one place.
        prim_sec_anchor_buf #(
          .Width(MuBi12Width)
        ) u_sig_unstable_buf (
          .in_i(sig_unstable),
          .out_o(sig_unstable_buf)
        );

        // if any xor indicates signal is unstable, output the reset
        // value. note that the input and output signals of this mux
        // are driven/read by constrained primitive cells (regs, buffers),
        // hence this mux can be implemented behaviorally.
        assign mubi[k] = (|sig_unstable_buf) ? reset_value[k] : mubi_q[k];
      end

// Note regarding SVAs below:
//
// 1) Without the sampled rst_ni pre-condition, this may cause false assertion failures right after
// a reset release, since the "disable iff" condition with the rst_ni is sampled in the "observed"
// SV scheduler region after all assignments have been evaluated (see also LRM section 16.12, page
// 423). This is a simulation artifact due to reset synchronization in RTL, which releases rst_ni
// on the active clock edge. This causes the assertion to evaluate although the reset was actually
// 0 when entering this simulation cycle.
//
// 2) Similarly to 1) there can be sampling mismatches of the lc_en_i signal since that signal may
// originate from a different clock domain. I.e., in cases where the lc_en_i signal changes exactly
// at the same time that the clk_i signal rises, the SVA will not pick up that change in that clock
// cycle, whereas RTL will because SVAs sample values in the "preponed" region. To that end we make
// use of an RTL helper variable to sample the lc_en_i signal, hence ensuring that there are no
// sampling mismatches.
`ifdef INC_ASSERT
      mubi12_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputIfUnstable_A, sig_unstable |-> mubi_o == {NumCopies{reset_value}})
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##[3:4] sig_unstable || mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}})
`endif
    end else begin : gen_no_stable_chks
      assign mubi = mubi_sync;
`ifdef INC_ASSERT
      mubi12_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##3 (mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}} ||
                              $past(mubi_in_sva_q, 2) != $past(mubi_in_sva_q, 1)))
`endif
    end
  end else begin : gen_no_flops

    //VCS coverage off
    // pragma coverage off

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for synthesis since it is unloaded.
    mubi12_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi12False;
      end else begin
         unused_logic <= mubi_i;
      end
    end

    //VCS coverage on
    // pragma coverage on

    assign mubi = MuBi12Width'(mubi_i);

    `ASSERT(OutputDelay_A, mubi_o == {NumCopies{mubi_i}})
  end

  for (genvar j = 0; j < NumCopies; j++) begin : gen_buffs
    logic [MuBi12Width-1:0] mubi_out;
    for (genvar k = 0; k < MuBi12Width; k++) begin : gen_bits
      prim_buf u_prim_buf (
        .in_i(mubi[k]),
        .out_o(mubi_out[k])
      );
    end
    assign mubi_o[j] = mubi12_t'(mubi_out);
  end

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi12_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Decoder for multibit control signals with additional input buffers.

`include "prim_assert.sv"

module prim_mubi12_dec
  import prim_mubi_pkg::*;
#(
  parameter bit TestTrue = 1,
  parameter bit TestStrict = 1
) (
  input  mubi12_t mubi_i,
  output logic           mubi_dec_o
);

logic [MuBi12Width-1:0] mubi, mubi_out;
assign mubi = MuBi12Width'(mubi_i);

// The buffer cells have a don't touch constraint on them
// such that synthesis tools won't collapse them
for (genvar k = 0; k < MuBi12Width; k++) begin : gen_bits
  prim_buf u_prim_buf (
    .in_i  ( mubi[k]     ),
    .out_o ( mubi_out[k] )
  );
end

if (TestTrue && TestStrict) begin : gen_test_true_strict
  assign mubi_dec_o = mubi12_test_true_strict(mubi12_t'(mubi_out));
end else if (TestTrue && !TestStrict) begin : gen_test_true_loose
  assign mubi_dec_o = mubi12_test_true_loose(mubi12_t'(mubi_out));
end else if (!TestTrue && TestStrict) begin : gen_test_false_strict
  assign mubi_dec_o = mubi12_test_false_strict(mubi12_t'(mubi_out));
end else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
  assign mubi_dec_o = mubi12_test_false_loose(mubi12_t'(mubi_out));
end else begin : gen_unknown_config
  `ASSERT_INIT(UnknownConfig_A, 0)
end

endmodule : prim_mubi12_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Multibit sender module. This module is instantiates a hand-picked flop cell for each bit in the
// multibit signal such that tools do not optimize the multibit encoding.

`include "prim_assert.sv"

module prim_mubi16_sender
  import prim_mubi_pkg::*;
#(
  // This flops the output if set to 1.
  // In special cases where the sender is in the same clock domain as the receiver,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // Enable anchor buffer
  parameter bit EnSecBuf = 0,
  // Reset value for the sender flops
  parameter mubi16_t ResetValue = MuBi16False
) (
  input          clk_i,
  input          rst_ni,
  input  mubi16_t mubi_i,
  output mubi16_t mubi_o
);

  logic [MuBi16Width-1:0] mubi, mubi_int, mubi_out;
  assign mubi = MuBi16Width'(mubi_i);

  // first generation block decides whether a flop should be present
  if (AsyncOn) begin : gen_flops
    prim_flop #(
      .Width(MuBi16Width),
      .ResetValue(MuBi16Width'(ResetValue))
    ) u_prim_flop (
      .clk_i,
      .rst_ni,
      .d_i   ( mubi     ),
      .q_o   ( mubi_int )
    );
  end else begin : gen_no_flops
    assign mubi_int = mubi;

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for sythesis since it is unloaded.
    mubi16_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi16False;
      end else begin
         unused_logic <= mubi_i;
      end
    end
  end

  // second generation block determines output buffer type
  // 1. If EnSecBuf -> always leads to a sec buffer regardless of first block
  // 2. If not EnSecBuf and not AsyncOn -> use normal buffer
  // 3. If not EnSecBuf and AsyncOn -> feed through
  if (EnSecBuf) begin : gen_sec_buf
    prim_sec_anchor_buf #(
      .Width(16)
    ) u_prim_sec_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else if (!AsyncOn) begin : gen_prim_buf
    prim_buf #(
      .Width(16)
    ) u_prim_buf (
      .in_i(mubi_int),
      .out_o(mubi_out)
    );
  end else begin : gen_feedthru
    assign mubi_out = mubi_int;
  end

  assign mubi_o = mubi16_t'(mubi_out);

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi16_sender


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Double-synchronizer flop for multibit signals with additional output buffers.

`include "prim_assert.sv"

module prim_mubi16_sync
  import prim_mubi_pkg::*;
#(
  // Number of separately buffered output signals.
  // The buffer cells have a don't touch constraint
  // on them such that synthesis tools won't collapse
  // all copies into one signal.
  parameter int NumCopies = 1,
  // This instantiates the synchronizer flops if set to 1.
  // In special cases where the receiver is in the same clock domain as the sender,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // This controls whether the mubi module institutes stability checks when
  // AsyncOn is set.  If stability checks are on, a 3rd stage of storage is
  // added after the synchronizers and the outputs only updated if the 3rd
  // stage and sychronizer agree.  If they do not agree, the ResetValue is
  // output instead.
  parameter bit StabilityCheck = 0,
  // Reset value for the sync flops
  parameter mubi16_t ResetValue = MuBi16False
) (
  input                          clk_i,
  input                          rst_ni,
  input  mubi16_t                 mubi_i,
  output mubi16_t [NumCopies-1:0] mubi_o
);

  `ASSERT_INIT(NumCopiesMustBeGreaterZero_A, NumCopies > 0)

  logic [MuBi16Width-1:0] mubi;
  if (AsyncOn) begin : gen_flops
    logic [MuBi16Width-1:0] mubi_sync;
    prim_flop_2sync #(
      .Width(MuBi16Width),
      .ResetValue(MuBi16Width'(ResetValue))
    ) u_prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(MuBi16Width'(mubi_i)),
      .q_o(mubi_sync)
    );

    if (StabilityCheck) begin : gen_stable_chks
      logic [MuBi16Width-1:0] mubi_q;
      prim_flop #(
        .Width(MuBi16Width),
        .ResetValue(MuBi16Width'(ResetValue))
      ) u_prim_flop_3rd_stage (
        .clk_i,
        .rst_ni,
        .d_i(mubi_sync),
        .q_o(mubi_q)
      );

      logic [MuBi16Width-1:0] sig_unstable;
      prim_xor2 #(
        .Width(MuBi16Width)
      ) u_mubi_xor (
        .in0_i(mubi_sync),
        .in1_i(mubi_q),
        .out_o(sig_unstable)
      );

      logic [MuBi16Width-1:0] reset_value;
      assign reset_value = ResetValue;

      for (genvar k = 0; k < MuBi16Width; k++) begin : gen_bufs_muxes
        logic [MuBi16Width-1:0] sig_unstable_buf;

        // each mux gets its own buffered output, this ensures the OR-ing
        // cannot be defeated in one place.
        prim_sec_anchor_buf #(
          .Width(MuBi16Width)
        ) u_sig_unstable_buf (
          .in_i(sig_unstable),
          .out_o(sig_unstable_buf)
        );

        // if any xor indicates signal is unstable, output the reset
        // value. note that the input and output signals of this mux
        // are driven/read by constrained primitive cells (regs, buffers),
        // hence this mux can be implemented behaviorally.
        assign mubi[k] = (|sig_unstable_buf) ? reset_value[k] : mubi_q[k];
      end

// Note regarding SVAs below:
//
// 1) Without the sampled rst_ni pre-condition, this may cause false assertion failures right after
// a reset release, since the "disable iff" condition with the rst_ni is sampled in the "observed"
// SV scheduler region after all assignments have been evaluated (see also LRM section 16.12, page
// 423). This is a simulation artifact due to reset synchronization in RTL, which releases rst_ni
// on the active clock edge. This causes the assertion to evaluate although the reset was actually
// 0 when entering this simulation cycle.
//
// 2) Similarly to 1) there can be sampling mismatches of the lc_en_i signal since that signal may
// originate from a different clock domain. I.e., in cases where the lc_en_i signal changes exactly
// at the same time that the clk_i signal rises, the SVA will not pick up that change in that clock
// cycle, whereas RTL will because SVAs sample values in the "preponed" region. To that end we make
// use of an RTL helper variable to sample the lc_en_i signal, hence ensuring that there are no
// sampling mismatches.
`ifdef INC_ASSERT
      mubi16_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputIfUnstable_A, sig_unstable |-> mubi_o == {NumCopies{reset_value}})
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##[3:4] sig_unstable || mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}})
`endif
    end else begin : gen_no_stable_chks
      assign mubi = mubi_sync;
`ifdef INC_ASSERT
      mubi16_t mubi_in_sva_q;
      always_ff @(posedge clk_i) begin
        mubi_in_sva_q <= mubi_i;
      end
      `ASSERT(OutputDelay_A,
              rst_ni |-> ##3 (mubi_o == {NumCopies{$past(mubi_in_sva_q, 2)}} ||
                              $past(mubi_in_sva_q, 2) != $past(mubi_in_sva_q, 1)))
`endif
    end
  end else begin : gen_no_flops

    //VCS coverage off
    // pragma coverage off

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // This logic will be removed for synthesis since it is unloaded.
    mubi16_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= MuBi16False;
      end else begin
         unused_logic <= mubi_i;
      end
    end

    //VCS coverage on
    // pragma coverage on

    assign mubi = MuBi16Width'(mubi_i);

    `ASSERT(OutputDelay_A, mubi_o == {NumCopies{mubi_i}})
  end

  for (genvar j = 0; j < NumCopies; j++) begin : gen_buffs
    logic [MuBi16Width-1:0] mubi_out;
    for (genvar k = 0; k < MuBi16Width; k++) begin : gen_bits
      prim_buf u_prim_buf (
        .in_i(mubi[k]),
        .out_o(mubi_out[k])
      );
    end
    assign mubi_o[j] = mubi16_t'(mubi_out);
  end

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, mubi_o)

endmodule : prim_mubi16_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
//    util/design/gen-mubi.py
//
// Decoder for multibit control signals with additional input buffers.

`include "prim_assert.sv"

module prim_mubi16_dec
  import prim_mubi_pkg::*;
#(
  parameter bit TestTrue = 1,
  parameter bit TestStrict = 1
) (
  input  mubi16_t mubi_i,
  output logic           mubi_dec_o
);

logic [MuBi16Width-1:0] mubi, mubi_out;
assign mubi = MuBi16Width'(mubi_i);

// The buffer cells have a don't touch constraint on them
// such that synthesis tools won't collapse them
for (genvar k = 0; k < MuBi16Width; k++) begin : gen_bits
  prim_buf u_prim_buf (
    .in_i  ( mubi[k]     ),
    .out_o ( mubi_out[k] )
  );
end

if (TestTrue && TestStrict) begin : gen_test_true_strict
  assign mubi_dec_o = mubi16_test_true_strict(mubi16_t'(mubi_out));
end else if (TestTrue && !TestStrict) begin : gen_test_true_loose
  assign mubi_dec_o = mubi16_test_true_loose(mubi16_t'(mubi_out));
end else if (!TestTrue && TestStrict) begin : gen_test_false_strict
  assign mubi_dec_o = mubi16_test_false_strict(mubi16_t'(mubi_out));
end else if (!TestTrue && !TestStrict) begin : gen_test_false_loose
  assign mubi_dec_o = mubi16_test_false_loose(mubi16_t'(mubi_out));
end else begin : gen_unknown_config
  `ASSERT_INIT(UnknownConfig_A, 0)
end

endmodule : prim_mubi16_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Spurious write-enable checker for autogenerated CSR node.
// This module has additional simulation features for error injection testing.

`include "prim_assert.sv"

module prim_reg_we_check #(
  parameter int unsigned OneHotWidth  = 32
) (
  // The module is combinational - the clock and reset are only used for assertions.
  input                          clk_i,
  input                          rst_ni,

  input  logic [OneHotWidth-1:0] oh_i,
  input  logic                   en_i,

  output logic                   err_o
);

  // Prevent optimization of the onehot input buffer.
  logic [OneHotWidth-1:0] oh_buf;
  prim_buf #(
    .Width(OneHotWidth)
  ) u_prim_buf (
    .in_i(oh_i),
    .out_o(oh_buf)
  );

  prim_onehot_check #(
    .OneHotWidth(OneHotWidth),
    .AddrWidth  (prim_util_pkg::vbits(OneHotWidth)),
    .EnableCheck(1),
    // Since certain peripherals may have a very large address space
    // (e.g. > 20bit), the inverse address decoding check (which is
    // essentially an indexing operation) does not scale well and is
    // hence omitted.
    .AddrCheck(0),
    // Due to REGWEN masking of write enable strobes,
    // we do not perform strict checks. I.e., we allow cases
    // where en_i is set to 1, but the oh_i vector is all-zeroes.
    .StrictCheck(0)
  ) u_prim_onehot_check (
    .clk_i,
    .rst_ni,
    .oh_i(oh_buf),
    .addr_i('0),
    .en_i,
    .err_o
  );

endmodule : prim_reg_we_check


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

`include "prim_assert.sv"

package lc_ctrl_pkg;

  import prim_util_pkg::vbits;
  import lc_ctrl_state_pkg::*;

  ///////////////////////////////////////
  // Netlist Constants (Hashed Tokens) //
  ///////////////////////////////////////

  parameter int NumTokens = 6;
  parameter int TokenIdxWidth = vbits(NumTokens);
  typedef enum logic [TokenIdxWidth-1:0] {
    // This is the index for the hashed all-zero constant.
    // All unconditional transitions use this token.
    ZeroTokenIdx       = 3'h0,
    RawUnlockTokenIdx  = 3'h1,
    TestUnlockTokenIdx = 3'h2,
    TestExitTokenIdx   = 3'h3,
    RmaTokenIdx        = 3'h4,
    // This is the index for an all-zero value (i.e., hashed value = '0).
    // This is used as an additional blocker for some invalid state transition edges.
    InvalidTokenIdx    = 3'h5
  } token_idx_e;

  parameter int TokenMuxBits = 2**TokenIdxWidth*LcTokenWidth;
  typedef logic [TokenMuxBits-1:0] lc_token_mux_t;

  ////////////////////////////////
  // Typedefs for LC Interfaces //
  ////////////////////////////////

  parameter int TxWidth = 4;

  // Note that changing this encoding has implications on isolation cell
  // values in RTL. Do not change this unless absolutely needed.
  typedef enum logic [TxWidth-1:0] {
    On  = 4'b0101,
    Off = 4'b1010
  } lc_tx_t;
  parameter lc_tx_t LC_TX_DEFAULT = lc_tx_t'(Off);

  parameter int RmaSeedWidth = 32;
  typedef logic [RmaSeedWidth-1:0] lc_flash_rma_seed_t;
  parameter lc_flash_rma_seed_t LC_FLASH_RMA_SEED_DEFAULT = '0;

  parameter int LcKeymgrDivWidth = 128;
  typedef logic [LcKeymgrDivWidth-1:0] lc_keymgr_div_t;

  typedef struct packed {
    logic [lc_ctrl_reg_pkg::SiliconCreatorIdWidth-1:0] silicon_creator_id;
    logic [lc_ctrl_reg_pkg::ProductIdWidth-1:0]        product_id;
    logic [lc_ctrl_reg_pkg::RevisionIdWidth-1:0]       revision_id;
    logic [32-lc_ctrl_reg_pkg::RevisionIdWidth-1:0]    reserved;
  } lc_hw_rev_t;

  /////////////////////////////////////////////
  // Helper Functions for Life Cycle Signals //
  /////////////////////////////////////////////

  // This is a prerequisite for the multibit functions below to work.
  `ASSERT_STATIC_IN_PACKAGE(CheckLcTxValsComplementary_A, On == ~Off)
  // Check for bit-width matching between lc_tx_t and mubi4_t
  `ASSERT_STATIC_IN_PACKAGE(LcMuBiWidthCheck_A, $bits(TxWidth) == $bits(prim_mubi_pkg::MuBi4Width))

  // Convert a life cycle signal to mubi4
  // If in the future other versions are desired, this should really be
  // moved to prim_mubi_pkg
  //
  // The On ^ MuBi4True determines the bit differences between
  // an lc_ctrl_pkg::On and prim_mubi_pkg::MuBi4True.
  // Once the required inversions are determined, it is then applied
  // to the incoming value.  If the incoming value is true, it will
  // appropriately flip to the correct MuBiValue.
  // Since the false value is always complement of the true value,
  // this mechanism will also work for the other polarity.
  function automatic prim_mubi_pkg::mubi4_t lc_to_mubi4(lc_tx_t val);
    return prim_mubi_pkg::mubi4_t'(val ^ (On ^ prim_mubi_pkg::MuBi4True));
  endfunction : lc_to_mubi4

  function automatic lc_tx_t mubi4_to_lc(prim_mubi_pkg::mubi4_t val);
    return lc_tx_t'(val ^ (prim_mubi_pkg::MuBi4True ^ On));
  endfunction : mubi4_to_lc

  // same function as above, but for an input that is MuBi4True, return Off
  // for an input that is MuBi4False, return On
  function automatic lc_tx_t mubi4_to_lc_inv(prim_mubi_pkg::mubi4_t val);
    return lc_tx_t'(val ^ (prim_mubi_pkg::MuBi4True ^ Off));
  endfunction : mubi4_to_lc_inv

  // Test whether the value is supplied is one of the valid enumerations
  function automatic logic lc_tx_test_invalid(lc_tx_t val);
    return ~(val inside {On, Off});
  endfunction : lc_tx_test_invalid

  // Convert a 1 input value to a lc_tx output
  function automatic lc_tx_t lc_tx_bool_to_lc_tx(logic val);
    return (val ? On : Off);
  endfunction : lc_tx_bool_to_lc_tx

  // Test whether the multibit value signals an "enabled" condition.
  // The strict version of this function requires
  // the multibit value to equal True.
  function automatic logic lc_tx_test_true_strict(lc_tx_t val);
    return On == val;
  endfunction : lc_tx_test_true_strict

  // Test whether the multibit value signals a "disabled" condition.
  // The strict version of this function requires
  // the multibit value to equal False.
  function automatic logic lc_tx_test_false_strict(lc_tx_t val);
    return Off == val;
  endfunction : lc_tx_test_false_strict

  // Test whether the multibit value signals an "enabled" condition.
  // The loose version of this function interprets all
  // values other than False as "enabled".
  function automatic logic lc_tx_test_true_loose(lc_tx_t val);
    return Off != val;
  endfunction : lc_tx_test_true_loose

  // Test whether the multibit value signals a "disabled" condition.
  // The loose version of this function interprets all
  // values other than True as "disabled".
  function automatic logic lc_tx_test_false_loose(lc_tx_t val);
    return On != val;
  endfunction : lc_tx_test_false_loose


  // Performs a logical OR operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | act
  // !act | act  | act
  // act  | act  | act
  //
  // Note: due to the nature of the lc_tx_or() function, it is possible that two
  // non-strictly "act" values may produce a strictly "act" value. If this is
  // of concern, e.g. if the output is consumed with a strict check on "act",
  // consider using the prim_lc_or_hardened primitive instead.
  function automatic lc_tx_t lc_tx_or(lc_tx_t a, lc_tx_t b, lc_tx_t act);
    logic [TxWidth-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < TxWidth; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] || b_in[k];
      end else begin
        out[k] = a_in[k] && b_in[k];
      end
    end
    return lc_tx_t'(out);
  endfunction : lc_tx_or

  // Performs a logical AND operation between two multibit values.
  // This treats "act" as logical 1, and all other values are
  // treated as 0. Truth table:
  //
  // A    | B    | OUT
  //------+------+-----
  // !act | !act | !act
  // act  | !act | !act
  // !act | act  | !act
  // act  | act  | act
  //
  // Noite: The lc_tx_and() function does not suffer from the strictness problem
  // that the lc_tx_or function above does, since only one output value in the
  // truth table is strictly "act". It can hence be used in most scenarios without issues.
  // If however the lc_tx_and() function should be strictly rectifying (i.e., only
  // output "act" or ~"act"), the prim_lc_and_hardened can be used.
  function automatic lc_tx_t lc_tx_and(lc_tx_t a, lc_tx_t b, lc_tx_t act);
    logic [TxWidth-1:0] a_in, b_in, act_in, out;
    a_in = a;
    b_in = b;
    act_in = act;
    for (int k = 0; k < TxWidth; k++) begin
      if (act_in[k]) begin
        out[k] = a_in[k] && b_in[k];
      end else begin
        out[k] = a_in[k] || b_in[k];
      end
    end
    return lc_tx_t'(out);
  endfunction : lc_tx_and

  // Performs a logical OR operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic lc_tx_t lc_tx_or_hi(lc_tx_t a, lc_tx_t b);
    return lc_tx_or(a, b, On);
  endfunction : lc_tx_or_hi

  // Performs a logical AND operation between two multibit values.
  // This treats "True" as logical 1, and all other values are
  // treated as 0.
  function automatic lc_tx_t lc_tx_and_hi(lc_tx_t a, lc_tx_t b);
    return lc_tx_and(a, b, On);
  endfunction : lc_tx_and_hi

  // Performs a logical OR operation between two multibit values.
  // This treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic lc_tx_t lc_tx_or_lo(lc_tx_t a, lc_tx_t b);
    return lc_tx_or(a, b, Off);
  endfunction : lc_tx_or_lo

  // Performs a logical AND operation between two multibit values.
  // Tlos treats "False" as logical 1, and all other values are
  // treated as 0.
  function automatic lc_tx_t lc_tx_and_lo(lc_tx_t a, lc_tx_t b);
    return lc_tx_and(a, b, Off);
  endfunction : lc_tx_and_lo

  // Inverts the logical meaning of the multibit value.
  function automatic lc_tx_t lc_tx_inv(lc_tx_t a);
    return lc_tx_t'(~TxWidth'(a));
  endfunction : lc_tx_inv

  ////////////////////
  // Main FSM State //
  ////////////////////

  // SEC_CM: MAIN.FSM.SPARSE
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 15 -n 16 \
  //      -s 2934212379 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: ||||||| (7.62%)
  //  6: ||||||||| (9.52%)
  //  7: |||||||||||||||| (17.14%)
  //  8: |||||||||||||||||||| (20.95%)
  //  9: ||||||||||||||||| (18.10%)
  // 10: ||||||||||||| (14.29%)
  // 11: |||||| (6.67%)
  // 12: ||| (3.81%)
  // 13: | (1.90%)
  // 14: --
  // 15: --
  // 16: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 13
  // Minimum Hamming weight: 3
  // Maximum Hamming weight: 11
  //
  localparam int FsmStateWidth = 16;
  typedef enum logic [FsmStateWidth-1:0] {
    ResetSt       = 16'b1111011010111100,
    IdleSt        = 16'b0000011110101101,
    ClkMuxSt      = 16'b1100111011001001,
    CntIncrSt     = 16'b0011001111000111,
    CntProgSt     = 16'b0000110001010100,
    TransCheckSt  = 16'b0110111010110000,
    TokenHashSt   = 16'b1101001000111111,
    FlashRmaSt    = 16'b1110100010001111,
    TokenCheck0St = 16'b0010000011000000,
    TokenCheck1St = 16'b1101010101101111,
    TransProgSt   = 16'b1000000110101011,
    PostTransSt   = 16'b0110110100101100,
    ScrapSt       = 16'b1010100001010001,
    EscalateSt    = 16'b1011110110011011,
    InvalidSt     = 16'b0011000101001100
  } fsm_state_e;

  ///////////////////////////////////////////
  // Manufacturing State Transition Matrix //
  ///////////////////////////////////////////

  // Helper macro to assemble the token index matrix below.
  // From TEST_UNLOCKED(N)
  // -> SCRAP, RMA
  // -> PROD, PROD_END, DEV
  // -> TEST_UNLOCKED(N+1)-7
  // -> TEST_LOCKED(N)-6
  // -> TEST_UNLOCKED0-(N), RAW
  `define TEST_UNLOCKED(idx)         \
        {2{ZeroTokenIdx}},           \
        {3{TestExitTokenIdx}},       \
        {(7-idx){InvalidTokenIdx,    \
                 ZeroTokenIdx}},     \
        {(2*idx+2){InvalidTokenIdx}}

  // Helper macro to assemble the token index matrix below.
  // From TEST_LOCKED(N)
  // -> SCRAP
  // -> RMA
  // -> PROD, PROD_END, DEV
  // -> TEST_UNLOCKED(N+1)-7
  // -> TEST_LOCKED(N)-6
  // -> TEST_UNLOCKED0-(N), RAW
  `define TEST_LOCKED(idx)         \
      ZeroTokenIdx,                \
      InvalidTokenIdx,             \
      {3{TestExitTokenIdx}},       \
      {(7-idx){TestUnlockTokenIdx, \
               InvalidTokenIdx}},  \
      {(2*idx+2){InvalidTokenIdx}}

  // The token index matrix below encodes 1) which transition edges are valid and 2) which token
  // to use for a given transition edge. Note that unconditional but otherwise valid transitions
  // are assigned the ZeroTokenIdx, whereas invalid transitions are assigned an InvalidTokenIdx.
  parameter token_idx_e [NumLcStates-1:0][NumLcStates-1:0] TransTokenIdxMatrix = {
    // SCRAP
    {21{InvalidTokenIdx}}, // -> TEST_LOCKED0-6, TEST_UNLOCKED0-7, DEV, PROD, PROD_END, RMA, SCRAP
    // RMA
    ZeroTokenIdx,          // -> SCRAP
    {20{InvalidTokenIdx}}, // -> TEST_LOCKED0-6, TEST_UNLOCKED0-7, DEV, PROD, PROD_END, RMA
    // PROD_END
    ZeroTokenIdx,          // -> SCRAP
    {20{InvalidTokenIdx}}, // -> TEST_LOCKED0-6, TEST_UNLOCKED0-7, DEV, PROD, PROD_END, RMA
    // PROD
    ZeroTokenIdx,          // -> SCRAP
    RmaTokenIdx,           // -> RMA
    {19{InvalidTokenIdx}}, // -> TEST_LOCKED0-6, TEST_UNLOCKED0-7, DEV, PROD, PROD_END
    // DEV
    ZeroTokenIdx,          // -> SCRAP
    RmaTokenIdx,           // -> RMA
    {19{InvalidTokenIdx}}, // -> TEST_LOCKED0-6, TEST_UNLOCKED0-7, DEV, PROD, PROD_END
    // TEST_UNLOCKED0-7, TEST_LOCKED0-6
    `TEST_UNLOCKED(7),
    `TEST_LOCKED(6),
    `TEST_UNLOCKED(6),
    `TEST_LOCKED(5),
    `TEST_UNLOCKED(5),
    `TEST_LOCKED(4),
    `TEST_UNLOCKED(4),
    `TEST_LOCKED(3),
    `TEST_UNLOCKED(3),
    `TEST_LOCKED(2),
    `TEST_UNLOCKED(2),
    `TEST_LOCKED(1),
    `TEST_UNLOCKED(1),
    `TEST_LOCKED(0),
    `TEST_UNLOCKED(0),
    // RAW
    ZeroTokenIdx,          // -> SCRAP
    {4{InvalidTokenIdx}},  // -> RMA, PROD, PROD_END, DEV
    {8{RawUnlockTokenIdx,  // -> TEST_UNLOCKED0-7
       InvalidTokenIdx}}   // -> RAW, TEST_LOCKED0-6
  };

  // These macros are only used locally.
  `undef TEST_LOCKED
  `undef TEST_UNLOCKED

endpackage : lc_ctrl_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

package rom_ctrl_pkg;

  parameter int AlertFatal = 0;

  typedef struct packed {
    prim_mubi_pkg::mubi4_t done;
    prim_mubi_pkg::mubi4_t good;
  } pwrmgr_data_t;

  parameter pwrmgr_data_t PWRMGR_DATA_DEFAULT = '{
    done: prim_mubi_pkg::MuBi4True,
    good: prim_mubi_pkg::MuBi4True
  };

  typedef struct packed {
    logic [255:0] data;
    logic         valid;
  } keymgr_data_t;

  //
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 7 -n 6 -s 2 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (57.14%)
  //  4: ||||||||||||||| (42.86%)
  //  5: --
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4
  //
  // However, we glom on an extra 4 bits to hold a mubi4_t that encodes "state == Done". The idea is
  // that we can use them for the rom_select_bus_o signal without needing an intermediate 1-bit
  // signal which would need burying.

  typedef enum logic [9:0] {
    ReadingLow  = {6'b001100, prim_mubi_pkg::MuBi4False},
    ReadingHigh = {6'b001011, prim_mubi_pkg::MuBi4False},
    RomAhead    = {6'b111001, prim_mubi_pkg::MuBi4False},
    KmacAhead   = {6'b100111, prim_mubi_pkg::MuBi4False},
    Checking    = {6'b010101, prim_mubi_pkg::MuBi4False},
    Done        = {6'b100000, prim_mubi_pkg::MuBi4True},
    Invalid     = {6'b010010, prim_mubi_pkg::MuBi4False}
  } fsm_state_e;


endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package rom_ctrl_reg_pkg;

  // Param list
  parameter int NumAlerts = 1;

  // Address widths within the block
  parameter int RegsAw = 7;
  parameter int RomAw = 15;

  ///////////////////////////////////////////////
  // Typedefs for registers for regs interface //
  ///////////////////////////////////////////////

  typedef struct packed {
    logic        q;
    logic        qe;
  } rom_ctrl_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } rom_ctrl_reg2hw_digest_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } rom_ctrl_reg2hw_exp_digest_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } checker_error;
    struct packed {
      logic        d;
      logic        de;
    } integrity_error;
  } rom_ctrl_hw2reg_fatal_alert_cause_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } rom_ctrl_hw2reg_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } rom_ctrl_hw2reg_exp_digest_mreg_t;

  // Register -> HW type for regs interface
  typedef struct packed {
    rom_ctrl_reg2hw_alert_test_reg_t alert_test; // [513:512]
    rom_ctrl_reg2hw_digest_mreg_t [7:0] digest; // [511:256]
    rom_ctrl_reg2hw_exp_digest_mreg_t [7:0] exp_digest; // [255:0]
  } rom_ctrl_regs_reg2hw_t;

  // HW -> register type for regs interface
  typedef struct packed {
    rom_ctrl_hw2reg_fatal_alert_cause_reg_t fatal_alert_cause; // [531:528]
    rom_ctrl_hw2reg_digest_mreg_t [7:0] digest; // [527:264]
    rom_ctrl_hw2reg_exp_digest_mreg_t [7:0] exp_digest; // [263:0]
  } rom_ctrl_regs_hw2reg_t;

  // Register offsets for regs interface
  parameter logic [RegsAw-1:0] ROM_CTRL_ALERT_TEST_OFFSET = 7'h 0;
  parameter logic [RegsAw-1:0] ROM_CTRL_FATAL_ALERT_CAUSE_OFFSET = 7'h 4;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_0_OFFSET = 7'h 8;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_1_OFFSET = 7'h c;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_2_OFFSET = 7'h 10;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_3_OFFSET = 7'h 14;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_4_OFFSET = 7'h 18;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_5_OFFSET = 7'h 1c;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_6_OFFSET = 7'h 20;
  parameter logic [RegsAw-1:0] ROM_CTRL_DIGEST_7_OFFSET = 7'h 24;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_0_OFFSET = 7'h 28;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_1_OFFSET = 7'h 2c;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_2_OFFSET = 7'h 30;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_3_OFFSET = 7'h 34;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_4_OFFSET = 7'h 38;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_5_OFFSET = 7'h 3c;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_6_OFFSET = 7'h 40;
  parameter logic [RegsAw-1:0] ROM_CTRL_EXP_DIGEST_7_OFFSET = 7'h 44;

  // Reset values for hwext registers and their fields for regs interface
  parameter logic [0:0] ROM_CTRL_ALERT_TEST_RESVAL = 1'h 0;
  parameter logic [0:0] ROM_CTRL_ALERT_TEST_FATAL_RESVAL = 1'h 0;

  // Register index for regs interface
  typedef enum int {
    ROM_CTRL_ALERT_TEST,
    ROM_CTRL_FATAL_ALERT_CAUSE,
    ROM_CTRL_DIGEST_0,
    ROM_CTRL_DIGEST_1,
    ROM_CTRL_DIGEST_2,
    ROM_CTRL_DIGEST_3,
    ROM_CTRL_DIGEST_4,
    ROM_CTRL_DIGEST_5,
    ROM_CTRL_DIGEST_6,
    ROM_CTRL_DIGEST_7,
    ROM_CTRL_EXP_DIGEST_0,
    ROM_CTRL_EXP_DIGEST_1,
    ROM_CTRL_EXP_DIGEST_2,
    ROM_CTRL_EXP_DIGEST_3,
    ROM_CTRL_EXP_DIGEST_4,
    ROM_CTRL_EXP_DIGEST_5,
    ROM_CTRL_EXP_DIGEST_6,
    ROM_CTRL_EXP_DIGEST_7
  } rom_ctrl_regs_id_e;

  // Register width information to check illegal writes for regs interface
  parameter logic [3:0] ROM_CTRL_REGS_PERMIT [18] = '{
    4'b 0001, // index[ 0] ROM_CTRL_ALERT_TEST
    4'b 0001, // index[ 1] ROM_CTRL_FATAL_ALERT_CAUSE
    4'b 1111, // index[ 2] ROM_CTRL_DIGEST_0
    4'b 1111, // index[ 3] ROM_CTRL_DIGEST_1
    4'b 1111, // index[ 4] ROM_CTRL_DIGEST_2
    4'b 1111, // index[ 5] ROM_CTRL_DIGEST_3
    4'b 1111, // index[ 6] ROM_CTRL_DIGEST_4
    4'b 1111, // index[ 7] ROM_CTRL_DIGEST_5
    4'b 1111, // index[ 8] ROM_CTRL_DIGEST_6
    4'b 1111, // index[ 9] ROM_CTRL_DIGEST_7
    4'b 1111, // index[10] ROM_CTRL_EXP_DIGEST_0
    4'b 1111, // index[11] ROM_CTRL_EXP_DIGEST_1
    4'b 1111, // index[12] ROM_CTRL_EXP_DIGEST_2
    4'b 1111, // index[13] ROM_CTRL_EXP_DIGEST_3
    4'b 1111, // index[14] ROM_CTRL_EXP_DIGEST_4
    4'b 1111, // index[15] ROM_CTRL_EXP_DIGEST_5
    4'b 1111, // index[16] ROM_CTRL_EXP_DIGEST_6
    4'b 1111  // index[17] ROM_CTRL_EXP_DIGEST_7
  };

  // Window parameters for rom interface
  parameter logic [RomAw-1:0] ROM_CTRL_ROM_OFFSET = 15'h 0;
  parameter int unsigned      ROM_CTRL_ROM_SIZE   = 'h 4000;

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module decodes a differentially encoded signal and detects
// incorrectly encoded differential states.
//
// In case the differential pair crosses an asynchronous boundary, it has
// to be re-synchronized to the local clock. This can be achieved by
// setting the AsyncOn parameter to 1'b1. In that case, two additional
// input registers are added (to counteract metastability), and
// a pattern detector is instantiated that detects skewed level changes on
// the differential pair (i.e., when level changes on the diff pair are
// sampled one cycle apart due to a timing skew between the two wires).
//
// See also: prim_alert_sender, prim_alert_receiver, alert_handler

`include "prim_assert.sv"

module prim_diff_decode #(
  // enables additional synchronization logic
  parameter bit AsyncOn = 1'b0
) (
  input        clk_i,
  input        rst_ni,
  // input diff pair
  input        diff_pi,
  input        diff_ni,
  // logical level and
  // detected edges
  output logic level_o,
  output logic rise_o,
  output logic fall_o,
  // either rise or fall
  output logic event_o,
  //signal integrity issue detected
  output logic sigint_o
);

  logic level_d, level_q;

  ///////////////////////////////////////////////////////////////
  // synchronization regs for incoming diff pair (if required) //
  ///////////////////////////////////////////////////////////////
  if (AsyncOn) begin : gen_async

    typedef enum logic [1:0] {IsStd, IsSkewed, SigInt} state_e;
    state_e state_d, state_q;
    logic diff_p_edge, diff_n_edge, diff_check_ok, level;

    // 2 sync regs, one reg for edge detection
    logic diff_pq, diff_nq, diff_pd, diff_nd;

    prim_flop_2sync #(
      .Width(1),
      .ResetValue('0)
    ) i_sync_p (
      .clk_i,
      .rst_ni,
      .d_i(diff_pi),
      .q_o(diff_pd)
    );

    prim_flop_2sync #(
      .Width(1),
      .ResetValue(1'b1)
    ) i_sync_n (
      .clk_i,
      .rst_ni,
      .d_i(diff_ni),
      .q_o(diff_nd)
    );

    // detect level transitions
    assign diff_p_edge   = diff_pq ^ diff_pd;
    assign diff_n_edge   = diff_nq ^ diff_nd;

    // detect sigint issue
    assign diff_check_ok = diff_pd ^ diff_nd;

    // this is the current logical level
    assign level         = diff_pd;

    // outputs
    assign level_o  = level_d;
    assign event_o = rise_o | fall_o;

    // sigint detection is a bit more involved in async case since
    // we might have skew on the diff pair, which can result in a
    // one cycle sampling delay between the two wires
    // so we need a simple pattern matcher
    // the following waves are legal
    // clk    |   |   |   |   |   |   |   |
    //           _______     _______
    // p _______/        ...        \________
    //   _______                     ________
    // n        \_______ ... _______/
    //              ____     ___
    // p __________/     ...    \________
    //   _______                     ________
    // n        \_______ ... _______/
    //
    // i.e., level changes may be off by one cycle - which is permissible
    // as long as this condition is only one cycle long.


    always_comb begin : p_diff_fsm
      // default
      state_d  = state_q;
      level_d  = level_q;
      rise_o   = 1'b0;
      fall_o   = 1'b0;
      sigint_o = 1'b0;

      unique case (state_q)
        // we remain here as long as
        // the diff pair is correctly encoded
        IsStd: begin
          if (diff_check_ok) begin
            level_d = level;
            if (diff_p_edge && diff_n_edge) begin
              if (level) begin
                rise_o = 1'b1;
              end else begin
                fall_o = 1'b1;
              end
            end
          end else begin
            if (diff_p_edge || diff_n_edge) begin
              state_d = IsSkewed;
            end else begin
              state_d = SigInt;
              sigint_o = 1'b1;
            end
          end
        end
        // diff pair must be correctly encoded, otherwise we got a sigint
        IsSkewed: begin
          if (diff_check_ok) begin
            state_d = IsStd;
            level_d = level;
            if (level) rise_o = 1'b1;
            else       fall_o = 1'b1;
          end else begin
            state_d  = SigInt;
            sigint_o = 1'b1;
          end
        end
        // Signal integrity issue detected, remain here
        // until resolved
        SigInt: begin
          sigint_o = 1'b1;
          if (diff_check_ok) begin
            state_d  = IsStd;
            sigint_o = 1'b0;
          end
        end
        default : ;
      endcase
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin : p_sync_reg
      if (!rst_ni) begin
        state_q  <= IsStd;
        diff_pq  <= 1'b0;
        diff_nq  <= 1'b1;
        level_q  <= 1'b0;
      end else begin
        state_q  <= state_d;
        diff_pq  <= diff_pd;
        diff_nq  <= diff_nd;
        level_q  <= level_d;
      end
    end

  //////////////////////////////////////////////////////////
  // fully synchronous case, no skew present in this case //
  //////////////////////////////////////////////////////////
  end else begin : gen_no_async
    logic diff_pq, diff_pd;

    // one reg for edge detection
    assign diff_pd = diff_pi;

    // incorrect encoding -> signal integrity issue
    assign sigint_o = ~(diff_pi ^ diff_ni);

    assign level_o = (sigint_o) ? level_q : diff_pi;
    assign level_d = level_o;

    // detect level transitions
    assign rise_o  = (~diff_pq &  diff_pi) & ~sigint_o;
    assign fall_o  = ( diff_pq & ~diff_pi) & ~sigint_o;
    assign event_o = rise_o | fall_o;

    always_ff @(posedge clk_i or negedge rst_ni) begin : p_edge_reg
      if (!rst_ni) begin
        diff_pq  <= 1'b0;
        level_q  <= 1'b0;
      end else begin
        diff_pq  <= diff_pd;
        level_q  <= level_d;
      end
    end
  end

  ////////////////
  // assertions //
  ////////////////

  // shared assertions
  // sigint -> level stays the same during sigint
  // $isunknown is needed to avoid false assertion in first clock cycle
  `ASSERT(SigintLevelCheck_A, ##1 sigint_o |-> $stable(level_o))
  // sigint -> no additional events asserted at output
  `ASSERT(SigintEventCheck_A, sigint_o |-> !event_o)
  `ASSERT(SigintRiseCheck_A,  sigint_o |-> !rise_o)
  `ASSERT(SigintFallCheck_A,  sigint_o |-> !fall_o)

  if (AsyncOn) begin : gen_async_assert
    // assertions for asynchronous case
`ifdef INC_ASSERT
  `ifndef FPV_ALERT_NO_SIGINT_ERR
    // correctly detect sigint issue (only one transition cycle of permissible due to skew)
    `ASSERT(SigintCheck0_A, gen_async.diff_pd == gen_async.diff_nd [*2] |-> sigint_o)
    // the synchronizer adds 2 cycles of latency with respect to input signals.
    `ASSERT(SigintCheck1_A,
        ##1 (gen_async.diff_pd ^ gen_async.diff_nd) &&
        $stable(gen_async.diff_pd) && $stable(gen_async.diff_nd) ##1
        $rose(gen_async.diff_pd) && $stable(gen_async.diff_nd) ##1
        $stable(gen_async.diff_pd) && $fell(gen_async.diff_nd)
        |-> rise_o)
    `ASSERT(SigintCheck2_A,
        ##1 (gen_async.diff_pd ^ gen_async.diff_nd) &&
        $stable(gen_async.diff_pd) && $stable(gen_async.diff_nd) ##1
        $fell(gen_async.diff_pd) && $stable(gen_async.diff_nd) ##1
        $stable(gen_async.diff_pd) && $rose(gen_async.diff_nd)
        |-> fall_o)
    `ASSERT(SigintCheck3_A,
        ##1 (gen_async.diff_pd ^ gen_async.diff_nd) &&
        $stable(gen_async.diff_pd) && $stable(gen_async.diff_nd) ##1
        $rose(gen_async.diff_nd) && $stable(gen_async.diff_pd) ##1
        $stable(gen_async.diff_nd) && $fell(gen_async.diff_pd)
        |-> fall_o)
    `ASSERT(SigintCheck4_A,
        ##1 (gen_async.diff_pd ^ gen_async.diff_nd) &&
        $stable(gen_async.diff_pd) && $stable(gen_async.diff_nd) ##1
        $fell(gen_async.diff_nd) && $stable(gen_async.diff_pd) ##1
        $stable(gen_async.diff_nd) && $rose(gen_async.diff_pd)
        |-> rise_o)
  `endif

    // correctly detect edges
    `ASSERT(RiseCheck_A,
        !sigint_o ##1 $rose(gen_async.diff_pd) && (gen_async.diff_pd ^ gen_async.diff_nd) |->
        ##[0:1] rise_o,  clk_i, !rst_ni || sigint_o)
    `ASSERT(FallCheck_A,
        !sigint_o ##1 $fell(gen_async.diff_pd) && (gen_async.diff_pd ^ gen_async.diff_nd) |->
        ##[0:1] fall_o,  clk_i, !rst_ni || sigint_o)
    `ASSERT(EventCheck_A,
        !sigint_o ##1 $changed(gen_async.diff_pd) && (gen_async.diff_pd ^ gen_async.diff_nd) |->
        ##[0:1] event_o, clk_i, !rst_ni || sigint_o)
    // correctly detect level
    `ASSERT(LevelCheck0_A,
        !sigint_o && (gen_async.diff_pd ^ gen_async.diff_nd) [*2] |->
        gen_async.diff_pd == level_o,
        clk_i, !rst_ni || sigint_o)
`endif
  end else begin : gen_sync_assert
    // assertions for synchronous case

  `ifndef FPV_ALERT_NO_SIGINT_ERR
    // correctly detect sigint issue
    `ASSERT(SigintCheck_A, diff_pi == diff_ni |-> sigint_o)
  `endif

    // correctly detect edges
    `ASSERT(RiseCheck_A,  ##1 $rose(diff_pi)    && (diff_pi ^ diff_ni) |->  rise_o)
    `ASSERT(FallCheck_A,  ##1 $fell(diff_pi)    && (diff_pi ^ diff_ni) |->  fall_o)
    `ASSERT(EventCheck_A, ##1 $changed(diff_pi) && (diff_pi ^ diff_ni) |-> event_o)
    // correctly detect level
    `ASSERT(LevelCheck_A, (diff_pi ^ diff_ni) |-> diff_pi == level_o)
  end

endmodule : prim_diff_decode


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Edge Detector

module prim_edge_detector #(
  parameter int unsigned Width = 1,

  parameter logic [Width-1:0] ResetValue = '0,

  // EnSync
  //
  // Enable Synchronizer to the input signal.
  // It is assumed that the input signal is glitch free (registered input).
  parameter bit EnSync  = 1'b 1
) (
  input clk_i,
  input rst_ni,

  input        [Width-1:0] d_i,
  output logic [Width-1:0] q_sync_o,

  output logic [Width-1:0] q_posedge_pulse_o,
  output logic [Width-1:0] q_negedge_pulse_o
);

  logic [Width-1:0] q_sync_d, q_sync_q;

  if (EnSync) begin : g_sync
    prim_flop_2sync #(
      .Width (Width),
      .ResetValue (ResetValue)
    ) u_sync (
      .clk_i,
      .rst_ni,
      .d_i,
      .q_o (q_sync_d)
    );
  end : g_sync
  else begin : g_nosync
    assign q_sync_d = d_i;
  end : g_nosync

  assign q_sync_o = q_sync_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) q_sync_q <= ResetValue;
    else         q_sync_q <= q_sync_d;
  end

  assign q_posedge_pulse_o = q_sync_d & ~q_sync_q;
  assign q_negedge_pulse_o = ~q_sync_d & q_sync_q;

endmodule : prim_edge_detector


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Generic Asynchronous SRAM FIFO (Dual port SRAM)

`include "prim_assert.sv"

module prim_fifo_async_sram_adapter #(
  parameter int unsigned Width = 32,
  parameter int unsigned Depth = 16,

  // SRAM parameters
  parameter int unsigned       SramAw = 16,

  // If SramDw > Width, upper data bits are 0.
  parameter int unsigned       SramDw = 32,
  parameter logic [SramAw-1:0] SramBaseAddr = 'h 0,

  // derived
  localparam int unsigned DepthW = $clog2(Depth+1)
) (
  // Write port
  input                     clk_wr_i,
  input                     rst_wr_ni,
  input                     wvalid_i,
  output logic              wready_o,
  input        [Width-1:0]  wdata_i,
  output logic [DepthW-1:0] wdepth_o,

  // Read port
  input                     clk_rd_i,
  input                     rst_rd_ni,
  output logic              rvalid_o,
  input                     rready_i,
  output logic [Width-1:0]  rdata_o,
  output logic [DepthW-1:0] rdepth_o,

  output logic r_full_o,
  output logic r_notempty_o,

  output logic w_full_o,

  // TODO: watermark(threshold) ?

  // SRAM interface
  // Write SRAM port
  output logic              w_sram_req_o,
  input                     w_sram_gnt_i,
  output logic              w_sram_write_o,
  output logic [SramAw-1:0] w_sram_addr_o,
  output logic [SramDw-1:0] w_sram_wdata_o,
  output logic [SramDw-1:0] w_sram_wmask_o,
  input                     w_sram_rvalid_i, // not used
  input        [SramDw-1:0] w_sram_rdata_i,  // not used
  input        [1:0]        w_sram_rerror_i, // not used

  // Read SRAM port
  output logic              r_sram_req_o,
  input                     r_sram_gnt_i,
  output logic              r_sram_write_o,
  output logic [SramAw-1:0] r_sram_addr_o,
  output logic [SramDw-1:0] r_sram_wdata_o, // not used
  output logic [SramDw-1:0] r_sram_wmask_o, // not used
  input                     r_sram_rvalid_i,
  input        [SramDw-1:0] r_sram_rdata_i,
  input        [1:0]        r_sram_rerror_i
);

  ////////////////
  // Definition //
  ////////////////
  // w_: write clock domain signals
  // r_: read clock domain signals

  // PtrVW: Pointer Value (without msb, flip) width
  localparam int unsigned PtrVW = $clog2(Depth);
  // PtrW: Read/Write pointer with flip bit
  localparam int unsigned PtrW  = PtrVW+1;

  ////////////
  // Signal //
  ////////////

  logic [PtrW-1:0]  w_wptr_q, w_wptr_d, w_wptr_gray_d, w_wptr_gray_q;
  logic [PtrW-1:0]  r_wptr_gray, r_wptr;
  logic [PtrVW-1:0] w_wptr_v, r_wptr_v;
  logic             w_wptr_p, r_wptr_p; // phase

  logic [PtrW-1:0]  r_rptr_q, r_rptr_d, r_rptr_gray_d, r_rptr_gray_q;
  logic [PtrW-1:0]  w_rptr_gray, w_rptr;
  logic [PtrVW-1:0] r_rptr_v, w_rptr_v;
  logic             r_rptr_p, w_rptr_p; // phase

  logic w_wptr_inc, r_rptr_inc;

  logic w_full, r_full, r_empty;

  // SRAM response one clock delayed. So store the value into read clock
  // domain
  logic             stored;
  logic [Width-1:0] rdata_q, rdata_d;

  // SRAM has another read pointer (for address of SRAM req)
  // It is -1 of r_rptr if stored, else same to r_rptr
  logic            r_sram_rptr_inc;
  logic [PtrW-1:0] r_sram_rptr;

  // r_sram_rptr == r_wptr
  // Used to determine r_sram_req
  logic r_sramrptr_empty;

  logic rfifo_ack; // Used to check if FIFO read interface consumes a data
  logic rsram_ack;

  //////////////
  // Datapath //
  //////////////

  // Begin: Write pointer sync to read clock ========================
  assign w_wptr_inc = wvalid_i & wready_o;

  assign w_wptr_d = w_wptr_q + PtrW'(1);

  always_ff @(posedge clk_wr_i or negedge rst_wr_ni) begin
    if (!rst_wr_ni) begin
      w_wptr_q      <= PtrW'(0);
      w_wptr_gray_q <= PtrW'(0);
    end else if (w_wptr_inc) begin
      w_wptr_q      <= w_wptr_d;
      w_wptr_gray_q <= w_wptr_gray_d;
    end
  end

  assign w_wptr_v = w_wptr_q[0+:PtrVW];
  assign w_wptr_p = w_wptr_q[PtrW-1];

  assign w_wptr_gray_d = dec2gray(w_wptr_d);

  prim_flop_2sync #(
    .Width (PtrW)
  ) u_sync_wptr_gray (
    .clk_i  (clk_rd_i),
    .rst_ni (rst_rd_ni),
    .d_i    (w_wptr_gray_q),
    .q_o    (r_wptr_gray)
  );

  assign r_wptr   = gray2dec(r_wptr_gray);
  assign r_wptr_p = r_wptr[PtrW-1];
  assign r_wptr_v = r_wptr[0+:PtrVW];

  assign wdepth_o = (w_wptr_p == w_rptr_p)
                  ? DepthW'(w_wptr_v - w_rptr_v)
                  : DepthW'({1'b1, w_wptr_v} - {1'b 0, w_rptr_v});
  // End:   Write pointer sync to read clock ------------------------

  // Begin: Read pointer sync to write clock ========================
  //assign r_rptr_inc = rvalid_o & rready_i;
  //assign r_rptr_inc = r_sram_req_o && r_sram_gnt_i;
  // Increase the read pointer (crossing the clock domain) only when the
  // reader acked.
  assign r_rptr_inc = rfifo_ack;

  assign r_rptr_d = r_rptr_q + PtrW'(1);

  always_ff @(posedge clk_rd_i or negedge rst_rd_ni) begin
    if (!rst_rd_ni) begin
      r_rptr_q      <= PtrW'(0);
      r_rptr_gray_q <= PtrW'(0);
    end else if (r_rptr_inc) begin
      r_rptr_q      <= r_rptr_d;
      r_rptr_gray_q <= r_rptr_gray_d;
    end
  end

  assign r_rptr_v = r_rptr_q[0+:PtrVW];
  assign r_rptr_p = r_rptr_q[PtrW-1];

  assign r_rptr_gray_d = dec2gray(r_rptr_d);

  prim_flop_2sync #(
    .Width (PtrW)
  ) u_sync_rptr_gray (
    .clk_i  (clk_wr_i),
    .rst_ni (rst_wr_ni),
    .d_i    (r_rptr_gray_q),
    .q_o    (w_rptr_gray)
  );

  assign w_rptr = gray2dec(w_rptr_gray);
  assign w_rptr_p = w_rptr[PtrW-1];
  assign w_rptr_v = w_rptr[0+:PtrVW];

  assign rdepth_o = (r_wptr_p == r_rptr_p)
                  ? DepthW'(r_wptr_v - r_rptr_v)
                  : DepthW'({1'b1, r_wptr_v} - {1'b 0, r_rptr_v});
  // End:   Read pointer sync to write clock ------------------------

  // Begin: SRAM Read pointer
  assign r_sram_rptr_inc = rsram_ack;

  always_ff @(posedge clk_rd_i or negedge rst_rd_ni) begin
    if (!rst_rd_ni) begin
      r_sram_rptr <= PtrW'(0);
    end else if (r_sram_rptr_inc) begin
      r_sram_rptr <= r_sram_rptr + PtrW'(1);
    end
  end

  assign r_sramrptr_empty = (r_wptr == r_sram_rptr);
  // End:   SRAM Read pointer

  // Full/ Empty
  // Lint complains PtrW'(1) << (PtrW-1). So changed as below
  localparam logic [PtrW-1:0] XorMask = {1'b 1, {PtrW-1{1'b0}}};
  assign w_full  = (w_wptr_q == (w_rptr   ^ XorMask));
  assign r_full  = (r_wptr   == (r_rptr_q ^ XorMask));
  assign r_empty = (r_wptr   == r_rptr_q);

  logic  unused_r_empty;
  assign unused_r_empty = r_empty;

  assign r_full_o     = r_full;
  assign w_full_o     = w_full;

  // The notempty status !(wptr == rptr) assert one clock earlier than the
  // actual `rvalid` signals.
  //
  // The reason is due to the SRAM read latency. The module uses SRAM FIFO
  // interface. When the logic in producer domain pushes entries, the pointer
  // is increased. This triggers the FIFO logic in the consumer clock domain
  // fetches data from SRAM.
  //
  // The pointer crosses the clock boundary. It takes usually two cycles (in
  // the consumer side). Then, as the read and write pointer in the read clock
  // domain has a gap by 1, the FIFO not empty status is raised.
  //
  // At this time, the logic just sent the read request to the SRAM. The data
  // is not yet read. The `rvalid` asserts when it receives data from the
  // SRAM.
  //
  // So, if the consumer reads data at the same cycle when notempty status is
  // raised, it reads incorrect data.
  assign r_notempty_o = rvalid_o;

  assign rsram_ack = r_sram_req_o && r_sram_gnt_i;
  assign rfifo_ack = rvalid_o     && rready_i;

  // SRAM Write Request
  assign w_sram_req_o   = wvalid_i && !w_full;
  assign wready_o       = !w_full && w_sram_gnt_i;
  assign w_sram_write_o = 1'b 1; // Always write
  assign w_sram_addr_o  = SramBaseAddr + SramAw'(w_wptr_v);

  assign w_sram_wdata_o = SramDw'(wdata_i);
  assign w_sram_wmask_o = SramDw'({Width{1'b1}});

  logic unused_w_sram;
  assign unused_w_sram = ^{w_sram_rvalid_i, w_sram_rdata_i, w_sram_rerror_i};

  // SRAM Read Request
  // Request Scenario (!r_empty):
  //  - storage empty: Send request if
  //               !r_sram_rvalid_i || (rfifo_ack && r_sram_rvalid_i);
  //  - storage !empty: depends on the rfifo_ack:
  //    - r_rptr_inc: Can request more
  //    - !r_rptr_inc: Can't request
  always_comb begin : r_sram_req
    r_sram_req_o = 1'b 0;
    // Karnough Map (!empty): sram_req
    // {sram_rv, rfifo_ack} | 00 | 01          | 11 | 10
    // ----------------------------------------------------------
    // stored          | 0  |  1 |  impossible |  1 |  0
    //                 | 1  |  0 |  1          |  X |  impossible
    //
    // req_o = r_ptr_inc || (!stored && !r_sram_rvalid_i)

    if (stored) begin
      // storage has data. depends on rfifo_ack
      // rfifo_ack can be replaced to rready_i as `rvalid_o` is 1
      r_sram_req_o = !r_sramrptr_empty && rfifo_ack;
    end else begin
      // storage has no data.
      // Can send request only when the reader accept the request or no
      // previous request sent out.
      r_sram_req_o = !r_sramrptr_empty && !(r_sram_rvalid_i ^ rfifo_ack);
    end
  end : r_sram_req

  assign rvalid_o       = stored || r_sram_rvalid_i;
  assign r_sram_write_o = 1'b 0; // always read
  assign r_sram_wdata_o = '0;
  assign r_sram_wmask_o = '0;

  // Send SRAM request with sram read pointer.
  assign r_sram_addr_o  = SramBaseAddr + SramAw'(r_sram_rptr[0+:PtrVW]);

  assign rdata_d = (r_sram_rvalid_i) ? r_sram_rdata_i[0+:Width] : Width'(0);

  assign rdata_o = (stored) ? rdata_q : rdata_d;

  logic unused_rsram;
  assign unused_rsram = ^{r_sram_rerror_i};

  if (Width < SramDw) begin : g_unused_rdata
    logic unused_rdata;
    assign unused_rdata = ^r_sram_rdata_i[SramDw-1:Width];
  end : g_unused_rdata

  // read clock domain rdata storage
  logic store_en;

  // Karnough Map (r_sram_rvalid_i):
  // rfifo_ack   | 0 | 1 |
  // ---------------------
  // stored    0 | 1 | 0 |
  //           1 | 0 | 1 |
  //
  // stored = s.r.v && XNOR(stored, rptr_inc)
  assign store_en = r_sram_rvalid_i && !(stored ^ rfifo_ack);

  always_ff @(posedge clk_rd_i or negedge rst_rd_ni) begin
    if (!rst_rd_ni) begin
      stored <= 1'b 0;
      rdata_q <= Width'(0);
    end else if (store_en) begin
      stored <= 1'b 1;
      rdata_q <= rdata_d;
    end else if (!r_sram_rvalid_i && rfifo_ack) begin
      // No request sent, host reads the data
      stored <= 1'b 0;
      rdata_q <= Width'(0);
    end
  end

  //////////////
  // Function //
  //////////////

  // dec2gray / gray2dec copied from prim_fifo_async.sv
  function automatic [PtrW-1:0] dec2gray(input logic [PtrW-1:0] decval);
    logic [PtrW-1:0] decval_sub;
    logic [PtrW-1:0] decval_in;
    logic            unused_decval_msb;

    decval_sub = (PtrW)'(Depth) - {1'b0, decval[PtrW-2:0]} - 1'b1;

    decval_in = decval[PtrW-1] ? decval_sub : decval;

    // We do not care about the MSB, hence we mask it out
    unused_decval_msb = decval_in[PtrW-1];
    decval_in[PtrW-1] = 1'b0;

    // Perform the XOR conversion
    dec2gray = decval_in;
    dec2gray ^= (decval_in >> 1);

    // Override the MSB
    dec2gray[PtrW-1] = decval[PtrW-1];
  endfunction

  // Algorithm walks up from 0..N-1 then flips the upper bit and walks down from N-1 to 0.
  function automatic [PtrW-1:0] gray2dec(input logic [PtrW-1:0] grayval);
    logic [PtrW-1:0] dec_tmp, dec_tmp_sub;
    logic            unused_decsub_msb;

    dec_tmp = '0;
    for (int i = PtrW-2; i >= 0; i--) begin
      dec_tmp[i] = dec_tmp[i+1] ^ grayval[i];
    end
    dec_tmp_sub = (PtrW)'(Depth) - dec_tmp - 1'b1;
    if (grayval[PtrW-1]) begin
      gray2dec = dec_tmp_sub;
      // Override MSB
      gray2dec[PtrW-1] = 1'b1;
      unused_decsub_msb = dec_tmp_sub[PtrW-1];
    end else begin
      gray2dec = dec_tmp;
    end
  endfunction

  ///////////////
  // Assertion //
  ///////////////

  `ASSERT_INIT(ParamCheckDepth_A, (Depth == 2**$clog2(Depth)))

  // Use FF if less than 4.
  `ASSERT_INIT(MinDepth_A, Depth >= 4)

  // SramDw greather than or equal to Width
  `ASSERT_INIT(WidthMatch_A, SramDw >= Width)

  // Not stored, Not read valid, but rptr_inc case is impossible
  `ASSERT(RptrIncDataValid_A,
          r_rptr_inc |-> stored || r_sram_rvalid_i,
          clk_rd_i, !rst_rd_ni)
  `ASSERT(SramRvalid_A,
          r_sram_rvalid_i |-> !stored || r_rptr_inc,
          clk_rd_i, !rst_rd_ni)

  // FIFO interface
  `ASSERT(NoWAckInFull_A, w_wptr_inc |-> !w_full,
          clk_wr_i, !rst_wr_ni)

  `ASSERT(WptrIncrease_A,
          w_wptr_inc |=> w_wptr_v == PtrVW'($past(w_wptr_v,2) + 1),
          clk_wr_i, !rst_wr_ni)
  `ASSERT(WptrGrayOneBitAtATime_A,
          w_wptr_inc |=> $countones(w_wptr_gray_q ^ $past(w_wptr_gray_q,2)) == 1,
          clk_wr_i, !rst_wr_ni)

  `ASSERT(NoRAckInEmpty_A, r_rptr_inc |-> !r_empty,
          clk_rd_i, !rst_rd_ni)

  `ASSERT(RptrIncrease_A,
          r_rptr_inc |=> PtrVW'($past(r_rptr_v) + 1) == r_rptr_v,
          clk_rd_i, !rst_rd_ni)
  `ASSERT(RptrGrayOneBitAtATime_A,
          r_rptr_inc |=> $countones(r_rptr_gray_q ^ $past(r_rptr_gray_q)) == 1,
          clk_rd_i, !rst_rd_ni)

  // SRAM interface
  `ASSERT(WSramRvalid_A, !w_sram_rvalid_i, clk_wr_i, !rst_wr_ni)
  `ASSUME_FPV(WSramRdataError_M, w_sram_rdata_i == '0 && w_sram_rerror_i == '0,
              clk_wr_i, !rst_wr_ni)

  `ASSUME(RSramRvalidOneCycle_M,
          r_sram_req_o && r_sram_gnt_i |=> r_sram_rvalid_i,
          clk_rd_i, !rst_rd_ni)
  `ASSUME_FPV(RErrorTied_M, r_sram_rerror_i == '0,
              clk_rd_i, !rst_rd_ni)


  // FPV coverage
  `COVER_FPV(WFull_C, w_full, clk_wr_i, !rst_wr_ni)

endmodule : prim_fifo_async_sram_adapter


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

`include "prim_assert.sv"

module prim_fifo_async_simple #(
  parameter int unsigned Width  = 16,
  parameter bit          EnRstChks = 1'b0, // Enable reset-related assertion checks, disabled by
                                           // default.
  parameter bit          EnRzHs = 1'b0     // By Default, the faster NRZ handshake protocol
                                           // (EnRzHs = 0) is used. Enable the RZ handshake protocol
                                           // if the FSMs need to be partial-reset-safe.
) (
  // write port
  input  logic              clk_wr_i,
  input  logic              rst_wr_ni,
  input  logic              wvalid_i,
  output logic              wready_o,
  input  logic [Width-1:0]  wdata_i,

  // read port
  input  logic              clk_rd_i,
  input  logic              rst_rd_ni,
  output logic              rvalid_o,
  input  logic              rready_i,
  output logic [Width-1:0]  rdata_o
);

  ////////////////
  // FIFO logic //
  ////////////////

  // Convert ready/valid to req/ack
  logic wr_en;
  logic src_req, src_ack;
  logic pending_d, pending_q, not_in_reset_q;
  assign wready_o = !pending_q && not_in_reset_q;
  assign wr_en = wvalid_i && wready_o;
  assign src_req = pending_q || wvalid_i;

  assign pending_d = (src_ack)  ? 1'b0 :
                     (wr_en)    ? 1'b1 : pending_q;

  logic dst_req, dst_ack;
  assign rvalid_o = dst_req;
  assign dst_ack = dst_req && rready_i;

  always_ff @(posedge clk_wr_i or negedge rst_wr_ni) begin
    if (!rst_wr_ni) begin
      pending_q <= 1'b0;
      not_in_reset_q <= 1'b0;
    end else begin
      pending_q <= pending_d;
      not_in_reset_q <= 1'b1;
    end
  end

  ////////////////////////////////////
  // REQ/ACK synchronizer primitive //
  ////////////////////////////////////

  prim_sync_reqack #(
    .EnRstChks(EnRstChks),
    .EnRzHs(EnRzHs)
  ) u_prim_sync_reqack (
    .clk_src_i(clk_wr_i),
    .rst_src_ni(rst_wr_ni),
    .clk_dst_i(clk_rd_i),
    .rst_dst_ni(rst_rd_ni),
    .req_chk_i(1'b0),
    .src_req_i(src_req),
    .src_ack_o(src_ack),
    .dst_req_o(dst_req),
    .dst_ack_i(dst_ack)
  );

  //////////////////////
  // Data holding reg //
  //////////////////////

  logic [Width-1:0] data_q;
  always_ff @(posedge clk_wr_i) begin
    if (wr_en) begin
      data_q <= wdata_i;
    end
  end
  assign rdata_o = data_q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Generic asynchronous fifo for use in a variety of devices.

`include "prim_assert.sv"

module prim_fifo_async #(
  parameter  int unsigned Width  = 16,
  parameter  int unsigned Depth  = 4,
  parameter  bit OutputZeroIfEmpty = 1'b0, // if == 1 always output 0 when FIFO is empty
  parameter  bit OutputZeroIfInvalid = 1'b0, // if == 1 always output 0 when rvalid_o is low
  localparam int unsigned DepthW = $clog2(Depth+1) // derived parameter representing [0..Depth]
) (
  // write port
  input  logic              clk_wr_i,
  input  logic              rst_wr_ni,
  input  logic              wvalid_i,
  output logic              wready_o,
  input  logic [Width-1:0]  wdata_i,
  output logic [DepthW-1:0] wdepth_o,

  // read port
  input  logic              clk_rd_i,
  input  logic              rst_rd_ni,
  output logic              rvalid_o,
  input  logic              rready_i,
  output logic [Width-1:0]  rdata_o,
  output logic [DepthW-1:0] rdepth_o
);

  // Depth must be a power of 2 for the gray code pointers to work
  `ASSERT_INIT(ParamCheckDepth_A, (Depth == 2**$clog2(Depth)))

  localparam int unsigned PTRV_W    = (Depth == 1) ? 1 : $clog2(Depth);
  localparam int unsigned PTR_WIDTH = (Depth == 1) ? 1 : PTRV_W+1;

  logic [PTR_WIDTH-1:0] fifo_wptr_q, fifo_wptr_d;
  logic [PTR_WIDTH-1:0] fifo_rptr_q, fifo_rptr_d;
  logic [PTR_WIDTH-1:0] fifo_wptr_sync_combi, fifo_rptr_sync_combi;
  logic [PTR_WIDTH-1:0] fifo_wptr_gray_sync, fifo_rptr_gray_sync, fifo_rptr_sync_q;
  logic [PTR_WIDTH-1:0] fifo_wptr_gray_q, fifo_wptr_gray_d;
  logic [PTR_WIDTH-1:0] fifo_rptr_gray_q, fifo_rptr_gray_d;
  logic                 fifo_incr_wptr, fifo_incr_rptr;
  logic                 full_wclk, full_rclk, empty_rclk;
  logic [Width-1:0]     storage [Depth];

  ///////////////////
  // Write Pointer //
  ///////////////////

  assign fifo_incr_wptr = wvalid_i & wready_o;

  // decimal version
  assign fifo_wptr_d = fifo_wptr_q + PTR_WIDTH'(1'b1);

  always_ff @(posedge clk_wr_i or negedge rst_wr_ni) begin
    if (!rst_wr_ni) begin
      fifo_wptr_q <= '0;
    end else if (fifo_incr_wptr) begin
      fifo_wptr_q <= fifo_wptr_d;
    end
  end

  // gray-coded version
  always_ff @(posedge clk_wr_i or negedge rst_wr_ni) begin
    if (!rst_wr_ni) begin
      fifo_wptr_gray_q <= '0;
    end else if (fifo_incr_wptr) begin
      fifo_wptr_gray_q <= fifo_wptr_gray_d;
    end
  end

  // sync gray-coded pointer to read clk
  prim_flop_2sync #(.Width(PTR_WIDTH)) sync_wptr (
    .clk_i    (clk_rd_i),
    .rst_ni   (rst_rd_ni),
    .d_i      (fifo_wptr_gray_q),
    .q_o      (fifo_wptr_gray_sync));

  //////////////////
  // Read Pointer //
  //////////////////

  assign fifo_incr_rptr = rvalid_o & rready_i;

  // decimal version
  assign fifo_rptr_d = fifo_rptr_q + PTR_WIDTH'(1'b1);

  always_ff @(posedge clk_rd_i or negedge rst_rd_ni) begin
    if (!rst_rd_ni) begin
      fifo_rptr_q <= '0;
    end else if (fifo_incr_rptr) begin
      fifo_rptr_q <= fifo_rptr_d;
    end
  end

  // gray-coded version
  always_ff @(posedge clk_rd_i or negedge rst_rd_ni) begin
    if (!rst_rd_ni) begin
      fifo_rptr_gray_q <= '0;
    end else if (fifo_incr_rptr) begin
      fifo_rptr_gray_q <= fifo_rptr_gray_d;
    end
  end

  // sync gray-coded pointer to write clk
  prim_flop_2sync #(.Width(PTR_WIDTH)) sync_rptr (
    .clk_i    (clk_wr_i),
    .rst_ni   (rst_wr_ni),
    .d_i      (fifo_rptr_gray_q),
    .q_o      (fifo_rptr_gray_sync));

  // Registered version of synced read pointer
  always_ff @(posedge clk_wr_i or negedge rst_wr_ni) begin
    if (!rst_wr_ni) begin
      fifo_rptr_sync_q <= '0;
    end else begin
      fifo_rptr_sync_q <= fifo_rptr_sync_combi;
    end
  end

  //////////////////
  // Empty / Full //
  //////////////////

  logic [PTR_WIDTH-1:0] xor_mask;
  assign xor_mask   =  PTR_WIDTH'(1'b1) << (PTR_WIDTH-1);
  assign full_wclk  = (fifo_wptr_q == (fifo_rptr_sync_q ^ xor_mask));
  assign full_rclk  = (fifo_wptr_sync_combi == (fifo_rptr_q ^ xor_mask));
  assign empty_rclk = (fifo_wptr_sync_combi ==  fifo_rptr_q);

  if (Depth > 1) begin : g_depth_calc

    // Current depth in the write clock side
    logic               wptr_msb;
    logic               rptr_sync_msb;
    logic  [PTRV_W-1:0] wptr_value;
    logic  [PTRV_W-1:0] rptr_sync_value;

    assign wptr_msb        = fifo_wptr_q[PTR_WIDTH-1];
    assign rptr_sync_msb   = fifo_rptr_sync_q[PTR_WIDTH-1];
    assign wptr_value      = fifo_wptr_q[0+:PTRV_W];
    assign rptr_sync_value = fifo_rptr_sync_q[0+:PTRV_W];
    assign wdepth_o = (full_wclk) ? DepthW'(Depth) :
                      (wptr_msb == rptr_sync_msb) ? DepthW'(wptr_value) - DepthW'(rptr_sync_value) :
                      (DepthW'(Depth) - DepthW'(rptr_sync_value) + DepthW'(wptr_value)) ;

    // Current depth in the read clock side
    logic               rptr_msb;
    logic               wptr_sync_msb;
    logic  [PTRV_W-1:0] rptr_value;
    logic  [PTRV_W-1:0] wptr_sync_value;

    assign wptr_sync_msb   = fifo_wptr_sync_combi[PTR_WIDTH-1];
    assign rptr_msb        = fifo_rptr_q[PTR_WIDTH-1];
    assign wptr_sync_value = fifo_wptr_sync_combi[0+:PTRV_W];
    assign rptr_value      = fifo_rptr_q[0+:PTRV_W];
    assign rdepth_o = (full_rclk) ? DepthW'(Depth) :
                      (wptr_sync_msb == rptr_msb) ? DepthW'(wptr_sync_value) - DepthW'(rptr_value) :
                      (DepthW'(Depth) - DepthW'(rptr_value) + DepthW'(wptr_sync_value)) ;

  end else begin : g_no_depth_calc

    assign rdepth_o = full_rclk;
    assign wdepth_o = full_wclk;

  end

  assign wready_o = ~full_wclk;
  assign rvalid_o = ~empty_rclk;

  /////////////
  // Storage //
  /////////////

  logic [Width-1:0] rdata_int;
  if (Depth > 1) begin : g_storage_mux

    always_ff @(posedge clk_wr_i) begin
      if (fifo_incr_wptr) begin
        storage[fifo_wptr_q[PTRV_W-1:0]] <= wdata_i;
      end
    end

    assign rdata_int = storage[fifo_rptr_q[PTRV_W-1:0]];

  end else begin : g_storage_simple

    always_ff @(posedge clk_wr_i) begin
      if (fifo_incr_wptr) begin
        storage[0] <= wdata_i;
      end
    end

    assign rdata_int = storage[0];

  end

  // rdata_o is qualified with rvalid_o to avoid CDC error
  if (OutputZeroIfEmpty == 1'b1) begin : gen_output_zero
    if (OutputZeroIfInvalid  == 1'b1) begin : gen_invalid_zero
      assign rdata_o = empty_rclk ? '0 : (rvalid_o ? rdata_int : '0);
    end
    else begin : gen_invalid_non_zero
      assign rdata_o = empty_rclk ? '0 : rdata_int;
    end
  end else begin : gen_no_output_zero
    if (OutputZeroIfInvalid  == 1'b1) begin : gen_invalid_zero
        assign rdata_o = rvalid_o ? rdata_int : '0;
    end
    else begin : gen_invalid_non_zero
        assign rdata_o = rdata_int;
    end
  end

  //////////////////////////////////////
  // Decimal <-> Gray-code Conversion //
  //////////////////////////////////////

  // This code is all in a generate context to avoid lint errors when Depth <= 2
  if (Depth > 2) begin : g_full_gray_conversion

    function automatic [PTR_WIDTH-1:0] dec2gray(input logic [PTR_WIDTH-1:0] decval);
      logic [PTR_WIDTH-1:0] decval_sub;
      logic [PTR_WIDTH-1:0] decval_in;
      logic                 unused_decval_msb;

      decval_sub = (PTR_WIDTH)'(Depth) - {1'b0, decval[PTR_WIDTH-2:0]} - 1'b1;

      decval_in = decval[PTR_WIDTH-1] ? decval_sub : decval;

      // We do not care about the MSB, hence we mask it out
      unused_decval_msb = decval_in[PTR_WIDTH-1];
      decval_in[PTR_WIDTH-1] = 1'b0;

      // Perform the XOR conversion
      dec2gray = decval_in;
      dec2gray ^= (decval_in >> 1);

      // Override the MSB
      dec2gray[PTR_WIDTH-1] = decval[PTR_WIDTH-1];
    endfunction

    // Algorithm walks up from 0..N-1 then flips the upper bit and walks down from N-1 to 0.
    function automatic [PTR_WIDTH-1:0] gray2dec(input logic [PTR_WIDTH-1:0] grayval);
      logic [PTR_WIDTH-1:0] dec_tmp, dec_tmp_sub;
      logic                 unused_decsub_msb;

      dec_tmp = '0;
      for (int i = PTR_WIDTH-2; i >= 0; i--) begin
        dec_tmp[i] = dec_tmp[i+1] ^ grayval[i];
      end
      dec_tmp_sub = (PTR_WIDTH)'(Depth) - dec_tmp - 1'b1;
      if (grayval[PTR_WIDTH-1]) begin
        gray2dec = dec_tmp_sub;
        // Override MSB
        gray2dec[PTR_WIDTH-1] = 1'b1;
        unused_decsub_msb = dec_tmp_sub[PTR_WIDTH-1];
      end else begin
        gray2dec = dec_tmp;
      end
    endfunction

    // decimal version of read pointer in write domain
    assign fifo_rptr_sync_combi = gray2dec(fifo_rptr_gray_sync);
    // decimal version of write pointer in read domain
    assign fifo_wptr_sync_combi = gray2dec(fifo_wptr_gray_sync);

    assign fifo_rptr_gray_d = dec2gray(fifo_rptr_d);
    assign fifo_wptr_gray_d = dec2gray(fifo_wptr_d);

  end else if (Depth == 2) begin : g_simple_gray_conversion

    assign fifo_rptr_sync_combi = {fifo_rptr_gray_sync[PTR_WIDTH-1], ^fifo_rptr_gray_sync};
    assign fifo_wptr_sync_combi = {fifo_wptr_gray_sync[PTR_WIDTH-1], ^fifo_wptr_gray_sync};

    assign fifo_rptr_gray_d = {fifo_rptr_d[PTR_WIDTH-1], ^fifo_rptr_d};
    assign fifo_wptr_gray_d = {fifo_wptr_d[PTR_WIDTH-1], ^fifo_wptr_d};

  end else begin : g_no_gray_conversion

    assign fifo_rptr_sync_combi = fifo_rptr_gray_sync;
    assign fifo_wptr_sync_combi = fifo_wptr_gray_sync;

    assign fifo_rptr_gray_d = fifo_rptr_d;
    assign fifo_wptr_gray_d = fifo_wptr_d;

  end

  // TODO: assertions on full, empty
  `ASSERT(GrayWptr_A, ##1 $countones(fifo_wptr_gray_q ^ $past(fifo_wptr_gray_q)) <= 1,
          clk_wr_i, !rst_wr_ni)
  `ASSERT(GrayRptr_A, ##1 $countones(fifo_rptr_gray_q ^ $past(fifo_rptr_gray_q)) <= 1,
          clk_rd_i, !rst_rd_ni)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Generic synchronous fifo for use in a variety of devices.

`include "prim_assert.sv"

module prim_fifo_sync #(
  parameter int unsigned Width       = 16,
  parameter bit Pass                 = 1'b1, // if == 1 allow requests to pass through empty FIFO
  parameter int unsigned Depth       = 4,
  parameter bit OutputZeroIfEmpty    = 1'b1, // if == 1 always output 0 when FIFO is empty
  parameter bit Secure               = 1'b0, // use prim count for pointers
  // derived parameter
  localparam int          DepthW     = prim_util_pkg::vbits(Depth+1)
) (
  input                   clk_i,
  input                   rst_ni,
  // synchronous clear / flush port
  input                   clr_i,
  // write port
  input                   wvalid_i,
  output                  wready_o,
  input   [Width-1:0]     wdata_i,
  // read port
  output                  rvalid_o,
  input                   rready_i,
  output  [Width-1:0]     rdata_o,
  // occupancy
  output                  full_o,
  output  [DepthW-1:0]    depth_o,
  output                  err_o
);


  // FIFO is in complete passthrough mode
  if (Depth == 0) begin : gen_passthru_fifo
    `ASSERT_INIT(paramCheckPass, Pass == 1)

    assign depth_o = 1'b0; //output is meaningless

    // devie facing
    assign rvalid_o = wvalid_i;
    assign rdata_o = wdata_i;

    // host facing
    assign wready_o = rready_i;
    assign full_o = rready_i;

    // this avoids lint warnings
    logic unused_clr;
    assign unused_clr = clr_i;

    // No error
    assign err_o = 1'b 0;

  // Normal FIFO construction
  end else begin : gen_normal_fifo

    localparam int unsigned PTRV_W    = prim_util_pkg::vbits(Depth);
    localparam int unsigned PTR_WIDTH = PTRV_W+1;

    logic [PTR_WIDTH-1:0] fifo_wptr, fifo_rptr;
    logic                 fifo_incr_wptr, fifo_incr_rptr, fifo_empty;

    // module under reset flag
    logic under_rst;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        under_rst <= 1'b1;
      end else if (under_rst) begin
        under_rst <= ~under_rst;
      end
    end

    // create the write and read pointers
    logic  full, empty;
    logic  wptr_msb;
    logic  rptr_msb;
    logic  [PTRV_W-1:0] wptr_value;
    logic  [PTRV_W-1:0] rptr_value;

    assign wptr_msb = fifo_wptr[PTR_WIDTH-1];
    assign rptr_msb = fifo_rptr[PTR_WIDTH-1];
    assign wptr_value = fifo_wptr[0+:PTRV_W];
    assign rptr_value = fifo_rptr[0+:PTRV_W];
    assign depth_o = (full)                 ? DepthW'(Depth) :
                     (wptr_msb == rptr_msb) ? DepthW'(wptr_value) - DepthW'(rptr_value) :
                     (DepthW'(Depth) - DepthW'(rptr_value) + DepthW'(wptr_value)) ;

    assign fifo_incr_wptr = wvalid_i & wready_o & ~under_rst;
    assign fifo_incr_rptr = rvalid_o & rready_i & ~under_rst;

    // full and not ready for write are two different concepts.
    // The latter can be '0' when under reset, while the former is an indication that no more
    // entries can be written.
    assign wready_o = ~full & ~under_rst;
    assign full_o   = full;
    assign rvalid_o = ~empty & ~under_rst;

    prim_fifo_sync_cnt #(
      .Width(PTR_WIDTH),
      .Depth(Depth),
      .Secure(Secure)
    ) u_fifo_cnt (
      .clk_i,
      .rst_ni,
      .clr_i,
      .incr_wptr_i(fifo_incr_wptr),
      .incr_rptr_i(fifo_incr_rptr),
      .wptr_o(fifo_wptr),
      .rptr_o(fifo_rptr),
      .err_o
    );

    //always_ff @(posedge clk_i or negedge rst_ni) begin
    //  if (!rst_ni) begin
    //    fifo_wptr <= {(PTR_WIDTH){1'b0}};
    //  end else if (clr_i) begin
    //    fifo_wptr <= {(PTR_WIDTH){1'b0}};
    //  end else if (fifo_incr_wptr) begin
    //    if (fifo_wptr[PTR_WIDTH-2:0] == (PTR_WIDTH-1)'(Depth-1)) begin
    //      fifo_wptr <= {~fifo_wptr[PTR_WIDTH-1],{(PTR_WIDTH-1){1'b0}}};
    //    end else begin
    //      fifo_wptr <= fifo_wptr + {{(PTR_WIDTH-1){1'b0}},1'b1};
    //    end
    //  end
    //end
    //
    //always_ff @(posedge clk_i or negedge rst_ni) begin
    //  if (!rst_ni) begin
    //    fifo_rptr <= {(PTR_WIDTH){1'b0}};
    //  end else if (clr_i) begin
    //    fifo_rptr <= {(PTR_WIDTH){1'b0}};
    //  end else if (fifo_incr_rptr) begin
    //    if (fifo_rptr[PTR_WIDTH-2:0] == (PTR_WIDTH-1)'(Depth-1)) begin
    //      fifo_rptr <= {~fifo_rptr[PTR_WIDTH-1],{(PTR_WIDTH-1){1'b0}}};
    //    end else begin
    //      fifo_rptr <= fifo_rptr + {{(PTR_WIDTH-1){1'b0}},1'b1};
    //    end
    //  end
    //end

    assign  full       = (fifo_wptr == (fifo_rptr ^ {1'b1,{(PTR_WIDTH-1){1'b0}}}));
    assign  fifo_empty = (fifo_wptr ==  fifo_rptr);


    // the generate blocks below are needed to avoid lint errors due to array indexing
    // in the where the fifo only has one storage element
    logic [Depth-1:0][Width-1:0] storage;
    logic [Width-1:0] storage_rdata;
    if (Depth == 1) begin : gen_depth_eq1
      assign storage_rdata = storage[0];

      always_ff @(posedge clk_i)
        if (fifo_incr_wptr) begin
          storage[0] <= wdata_i;
        end
    // fifo with more than one storage element
    end else begin : gen_depth_gt1
      assign storage_rdata = storage[fifo_rptr[PTR_WIDTH-2:0]];

      always_ff @(posedge clk_i)
        if (fifo_incr_wptr) begin
          storage[fifo_wptr[PTR_WIDTH-2:0]] <= wdata_i;
        end
    end

    logic [Width-1:0] rdata_int;
    if (Pass == 1'b1) begin : gen_pass
      assign rdata_int = (fifo_empty && wvalid_i) ? wdata_i : storage_rdata;
      assign empty = fifo_empty & ~wvalid_i;
    end else begin : gen_nopass
      assign rdata_int = storage_rdata;
      assign empty = fifo_empty;
    end

    if (OutputZeroIfEmpty == 1'b1) begin : gen_output_zero
      assign rdata_o = empty ? 'b0 : rdata_int;
    end else begin : gen_no_output_zero
      assign rdata_o = rdata_int;
    end

    `ASSERT(depthShallNotExceedParamDepth, !empty |-> depth_o <= DepthW'(Depth))
  end // block: gen_normal_fifo


  //////////////////////
  // Known Assertions //
  //////////////////////

  `ASSERT(DataKnown_A, rvalid_o |-> !$isunknown(rdata_o))
  `ASSERT_KNOWN(DepthKnown_A, depth_o)
  `ASSERT_KNOWN(RvalidKnown_A, rvalid_o)
  `ASSERT_KNOWN(WreadyKnown_A, wready_o)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Generic synchronous fifo for use in a variety of devices.

`include "prim_assert.sv"

module prim_fifo_sync_cnt #(
  parameter int Depth = 4,
  parameter int Width = 16,
  parameter bit Secure = 1'b0
) (
  input clk_i,
  input rst_ni,
  input clr_i,
  input incr_wptr_i,
  input incr_rptr_i,
  output logic [Width-1:0] wptr_o,
  output logic [Width-1:0] rptr_o,
  output logic err_o
);

  logic wptr_wrap;
  logic [Width-1:0] wptr_wrap_cnt;
  logic rptr_wrap;
  logic [Width-1:0] rptr_wrap_cnt;

  assign wptr_wrap = incr_wptr_i & (wptr_o[Width-2:0] == unsigned'((Width-1)'(Depth-1)));
  assign rptr_wrap = incr_rptr_i & (rptr_o[Width-2:0] == unsigned'((Width-1)'(Depth-1)));

  assign wptr_wrap_cnt = {~wptr_o[Width-1],{(Width-1){1'b0}}};
  assign rptr_wrap_cnt = {~rptr_o[Width-1],{(Width-1){1'b0}}};

  if (Secure) begin : gen_secure_ptrs
    logic wptr_err;
    prim_count #(
      .Width(Width)
    ) u_wptr (
      .clk_i,
      .rst_ni,
      .clr_i,
      .set_i(wptr_wrap),
      .set_cnt_i(wptr_wrap_cnt),
      .incr_en_i(incr_wptr_i),
      .decr_en_i(1'b0),
      .step_i(Width'(1'b1)),
      .cnt_o(wptr_o),
      .cnt_next_o(),
      .err_o(wptr_err)
    );

    logic rptr_err;
    prim_count #(
      .Width(Width)
    ) u_rptr (
      .clk_i,
      .rst_ni,
      .clr_i,
      .set_i(rptr_wrap),
      .set_cnt_i(rptr_wrap_cnt),
      .incr_en_i(incr_rptr_i),
      .decr_en_i(1'b0),
      .step_i(Width'(1'b1)),
      .cnt_o(rptr_o),
      .cnt_next_o(),
      .err_o(rptr_err)
    );

    assign err_o = wptr_err | rptr_err;

  end else begin : gen_normal_ptrs
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        wptr_o <= {(Width){1'b0}};
      end else if (clr_i) begin
        wptr_o <= {(Width){1'b0}};
      end else if (wptr_wrap) begin
        wptr_o <= wptr_wrap_cnt;
      end else if (incr_wptr_i) begin
        wptr_o <= wptr_o + {{(Width-1){1'b0}},1'b1};
      end
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        rptr_o <= {(Width){1'b0}};
      end else if (clr_i) begin
        rptr_o <= {(Width){1'b0}};
      end else if (rptr_wrap) begin
         rptr_o <= rptr_wrap_cnt;
      end else if (incr_rptr_i) begin
         rptr_o <= rptr_o + {{(Width-1){1'b0}},1'b1};
      end
    end

    assign err_o = '0;
  end



endmodule // prim_fifo_sync_cnt


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Single-Port SRAM Wrapper
//
// Supported configurations:
// - ECC for 32b and 64b wide memories with no write mask
//   (Width == 32 or Width == 64, DataBitsPerMask is ignored).
// - Byte parity if Width is a multiple of 8 bit and write masks have Byte
//   granularity (DataBitsPerMask == 8).
//
// Note that the write mask needs to be per Byte if parity is enabled. If ECC is enabled, the write
// mask cannot be used and has to be tied to {Width{1'b1}}.

`include "prim_assert.sv"

module prim_ram_1p_adv import prim_ram_1p_pkg::*; #(
  parameter  int Depth                = 512,
  parameter  int Width                = 32,
  parameter  int DataBitsPerMask      = 1,  // Number of data bits per bit of write mask
  parameter      MemInitFile          = "", // VMEM file to initialize the memory with

  // Configurations
  parameter  bit EnableECC            = 0, // Enables per-word ECC
  parameter  bit EnableParity         = 0, // Enables per-Byte Parity
  parameter  bit EnableInputPipeline  = 0, // Adds an input register (read latency +1)
  parameter  bit EnableOutputPipeline = 0, // Adds an output register (read latency +1)

  // This switch allows to switch to standard Hamming ECC instead of the HSIAO ECC.
  // It is recommended to leave this parameter at its default setting (HSIAO),
  // since this results in a more compact and faster implementation.
  parameter bit HammingECC            = 0,

  localparam int Aw                   = prim_util_pkg::vbits(Depth)
) (
  input clk_i,
  input rst_ni,

  input                      req_i,
  input                      write_i,
  input        [Aw-1:0]      addr_i,
  input        [Width-1:0]   wdata_i,
  input        [Width-1:0]   wmask_i,
  output logic [Width-1:0]   rdata_o,
  output logic               rvalid_o, // read response (rdata_o) is valid
  output logic [1:0]         rerror_o, // Bit1: Uncorrectable, Bit0: Correctable

  // config
  input ram_1p_cfg_t         cfg_i
);


  `ASSERT_INIT(CannotHaveEccAndParity_A, !(EnableParity && EnableECC))

  // Calculate ECC width
  localparam int ParWidth  = (EnableParity) ? Width/8 :
                             (!EnableECC)   ? 0 :
                             (Width <=   4) ? 4 :
                             (Width <=  11) ? 5 :
                             (Width <=  26) ? 6 :
                             (Width <=  57) ? 7 :
                             (Width <= 120) ? 8 : 8 ;
  localparam int TotalWidth = Width + ParWidth;

  // If byte parity is enabled, the write enable bits are used to write memory colums
  // with 8 + 1 = 9 bit width (data plus corresponding parity bit).
  // If ECC is enabled, the DataBitsPerMask is ignored.
  localparam int LocalDataBitsPerMask = (EnableParity) ? 9          :
                                        (EnableECC)    ? TotalWidth :
                                                         DataBitsPerMask;

  ////////////////////////////
  // RAM Primitive Instance //
  ////////////////////////////

  logic                    req_q,    req_d ;
  logic                    write_q,  write_d ;
  logic [Aw-1:0]           addr_q,   addr_d ;
  logic [TotalWidth-1:0]   wdata_q,  wdata_d ;
  logic [TotalWidth-1:0]   wmask_q,  wmask_d ;
  logic                    rvalid_q, rvalid_d, rvalid_sram_q ;
  logic [Width-1:0]        rdata_q,  rdata_d ;
  logic [TotalWidth-1:0]   rdata_sram ;
  logic [1:0]              rerror_q, rerror_d ;

  prim_ram_1p #(
    .MemInitFile     (MemInitFile),

    .Width           (TotalWidth),
    .Depth           (Depth),
    .DataBitsPerMask (LocalDataBitsPerMask)
  ) u_mem (
    .clk_i,

    .req_i    (req_q),
    .write_i  (write_q),
    .addr_i   (addr_q),
    .wdata_i  (wdata_q),
    .wmask_i  (wmask_q),
    .rdata_o  (rdata_sram),
    .cfg_i
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rvalid_sram_q <= 1'b0;
    end else begin
      rvalid_sram_q <= req_q & ~write_q;
    end
  end

  assign req_d              = req_i;
  assign write_d            = write_i;
  assign addr_d             = addr_i;
  assign rvalid_o           = rvalid_q;
  assign rdata_o            = rdata_q;
  assign rerror_o           = rerror_q;

  /////////////////////////////
  // ECC / Parity Generation //
  /////////////////////////////

  if (EnableParity == 0 && EnableECC) begin : gen_secded
    logic unused_wmask;
    assign unused_wmask = ^wmask_i;

    // check supported widths
    `ASSERT_INIT(SecDecWidth_A, Width inside {16, 32})

    // the wmask is constantly set to 1 in this case
    `ASSERT(OnlyWordWritePossibleWithEccPortA_A, req_i |->
          wmask_i == {Width{1'b1}})

    assign wmask_d = {TotalWidth{1'b1}};

    if (Width == 16) begin : gen_secded_22_16
      if (HammingECC) begin : gen_hamming
        prim_secded_inv_hamming_22_16_enc u_enc (
          .data_i(wdata_i),
          .data_o(wdata_d)
        );
        prim_secded_inv_hamming_22_16_dec u_dec (
          .data_i     (rdata_sram),
          .data_o     (rdata_d[0+:Width]),
          .syndrome_o ( ),
          .err_o      (rerror_d)
        );
      end else begin : gen_hsiao
        prim_secded_inv_22_16_enc u_enc (
          .data_i(wdata_i),
          .data_o(wdata_d)
        );
        prim_secded_inv_22_16_dec u_dec (
          .data_i     (rdata_sram),
          .data_o     (rdata_d[0+:Width]),
          .syndrome_o ( ),
          .err_o      (rerror_d)
        );
      end
    end else if (Width == 32) begin : gen_secded_39_32
      if (HammingECC) begin : gen_hamming
        prim_secded_inv_hamming_39_32_enc u_enc (
          .data_i(wdata_i),
          .data_o(wdata_d)
        );
        prim_secded_inv_hamming_39_32_dec u_dec (
          .data_i     (rdata_sram),
          .data_o     (rdata_d[0+:Width]),
          .syndrome_o ( ),
          .err_o      (rerror_d)
        );
      end else begin : gen_hsiao
        prim_secded_inv_39_32_enc u_enc (
          .data_i(wdata_i),
          .data_o(wdata_d)
        );
        prim_secded_inv_39_32_dec u_dec (
          .data_i     (rdata_sram),
          .data_o     (rdata_d[0+:Width]),
          .syndrome_o ( ),
          .err_o      (rerror_d)
        );
      end
    end

  end else if (EnableParity) begin : gen_byte_parity

    `ASSERT_INIT(WidthNeedsToBeByteAligned_A, Width % 8 == 0)
    `ASSERT_INIT(ParityNeedsByteWriteMask_A, DataBitsPerMask == 8)

    always_comb begin : p_parity
      rerror_d = '0;
      for (int i = 0; i < Width/8; i ++) begin
        // Data mapping. We have to make 8+1 = 9 bit groups
        // that have the same write enable such that FPGA tools
        // can map this correctly to BRAM resources.
        wmask_d[i*9 +: 8] = wmask_i[i*8 +: 8];
        wdata_d[i*9 +: 8] = wdata_i[i*8 +: 8];
        rdata_d[i*8 +: 8] = rdata_sram[i*9 +: 8];

        // parity generation (odd parity)
        wdata_d[i*9 + 8] = ~(^wdata_i[i*8 +: 8]);
        wmask_d[i*9 + 8] = &wmask_i[i*8 +: 8];
        // parity decoding (errors are always uncorrectable)
        rerror_d[1] |= ~(^{rdata_sram[i*9 +: 8], rdata_sram[i*9 + 8]});
      end
    end
  end else begin : gen_nosecded_noparity
    assign wmask_d = wmask_i;
    assign wdata_d = wdata_i;

    assign rdata_d  = rdata_sram[0+:Width];
    assign rerror_d = '0;
  end

  assign rvalid_d = rvalid_sram_q;

  /////////////////////////////////////
  // Input/Output Pipeline Registers //
  /////////////////////////////////////

  if (EnableInputPipeline) begin : gen_regslice_input
    // Put the register slices between ECC encoding to SRAM port
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        req_q   <= '0;
        write_q <= '0;
        addr_q  <= '0;
        wdata_q <= '0;
        wmask_q <= '0;
      end else begin
        req_q   <= req_d;
        write_q <= write_d;
        addr_q  <= addr_d;
        wdata_q <= wdata_d;
        wmask_q <= wmask_d;
      end
    end
  end else begin : gen_dirconnect_input
    assign req_q   = req_d;
    assign write_q = write_d;
    assign addr_q  = addr_d;
    assign wdata_q = wdata_d;
    assign wmask_q = wmask_d;
  end

  if (EnableOutputPipeline) begin : gen_regslice_output
    // Put the register slices between ECC decoding to output
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        rvalid_q <= '0;
        rdata_q  <= '0;
        rerror_q <= '0;
      end else begin
        rvalid_q <= rvalid_d;
        rdata_q  <= rdata_d;
        // tie to zero if the read data is not valid
        rerror_q <= rerror_d & {2{rvalid_d}};
      end
    end
  end else begin : gen_dirconnect_output
    assign rvalid_q = rvalid_d;
    assign rdata_q  = rdata_d;
    // tie to zero if the read data is not valid
    assign rerror_q = rerror_d & {2{rvalid_d}};
  end

endmodule : prim_ram_1p_adv


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ROM wrapper with rvalid register

`include "prim_assert.sv"

module prim_rom_adv import prim_rom_pkg::*; #(
  // Parameters passed on the ROM primitive.
  parameter  int Width       = 32,
  parameter  int Depth       = 2048, // 8kB default
  parameter      MemInitFile = "", // VMEM file to initialize the memory with

  localparam int Aw          = $clog2(Depth)
) (
  input  logic             clk_i,
  input  logic             rst_ni,
  input  logic             req_i,
  input  logic [Aw-1:0]    addr_i,
  output logic             rvalid_o,
  output logic [Width-1:0] rdata_o,

  input rom_cfg_t          cfg_i
);

  prim_rom #(
    .Width(Width),
    .Depth(Depth),
    .MemInitFile(MemInitFile)
  ) u_prim_rom (
    .clk_i,
    .req_i,
    .addr_i,
    .rdata_o,
    .cfg_i
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rvalid_o <= 1'b0;
    end else begin
      rvalid_o <= req_i;
    end
  end

  ////////////////
  // ASSERTIONS //
  ////////////////

  // Control Signals should never be X
  `ASSERT(noXOnCsI, !$isunknown(req_i), clk_i, '0)
endmodule : prim_rom_adv


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Reset synchronizer
/** Conventional 2FF async assert sync de-assert reset synchronizer
 *
 */

module prim_rst_sync #(
  // ActiveHigh should be 0 if the input reset is active low reset
  parameter bit ActiveHigh = 1'b 0,

  // In certain case, Scan may be inserted at the following reset chain.
  // Set SkipScan to 1'b 1 in that case.
  parameter bit SkipScan   = 1'b 0
) (
  input        clk_i,
  input        d_i, // raw reset (not synched to clk_i)
  output logic q_o, // reset synched to clk_i

  // Scan chain
  input                        scan_rst_ni,
  input prim_mubi_pkg::mubi4_t scanmode_i
);

  logic async_rst_n, scan_rst;
  logic rst_sync;

  // TODO: Check if 2FF set can be used.
  if (ActiveHigh == 1'b 1) begin : g_rst_inv
    assign async_rst_n = ~d_i;
    assign scan_rst    = ~scan_rst_ni;
  end else begin : g_rst_direct
    assign async_rst_n = d_i;
    assign scan_rst    = scan_rst_ni;
  end

  prim_flop_2sync #(
    .Width        (1),
    .ResetValue   (ActiveHigh)
  ) u_sync (
    .clk_i,
    .rst_ni (async_rst_n),
    .d_i    (!ActiveHigh), // reset release value
    .q_o    (rst_sync   )
  );

  if (SkipScan) begin : g_skip_scan
    logic  unused_scan;
    assign unused_scan = ^{scan_rst, scanmode_i};

    assign q_o = rst_sync;
  end else begin : g_scan_mux
    prim_clock_mux2 #(
      .NoFpgaBufG(1'b1)
    ) u_scan_mux (
      .clk0_i(rst_sync                                         ),
      .clk1_i(scan_rst                                         ),
      .sel_i (prim_mubi_pkg::mubi4_test_true_strict(scanmode_i)),
      .clk_o (q_o                                              )
    );
  end

endmodule : prim_rst_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package tlul_pkg;

  // this can be either PPC or BINTREE
  // there is no functional difference, but timing and area behavior is different
  // between the two instances. PPC can result in smaller implementations when timing
  // is not critical, whereas BINTREE is favorable when timing pressure is high (but this
  // may also result in a larger implementation). on FPGA targets, BINTREE is favorable
  // both in terms of area and timing.
  parameter ArbiterImpl = "PPC";

  typedef enum logic [2:0] {
    PutFullData    = 3'h 0,
    PutPartialData = 3'h 1,
    Get            = 3'h 4
  } tl_a_op_e;

  typedef enum logic [2:0] {
    AccessAck     = 3'h 0,
    AccessAckData = 3'h 1
  } tl_d_op_e;

  parameter int H2DCmdMaxWidth  = 57;
  parameter int H2DCmdIntgWidth = 7;
  parameter int H2DCmdFullWidth = H2DCmdMaxWidth + H2DCmdIntgWidth;
  parameter int D2HRspMaxWidth  = 57;
  parameter int D2HRspIntgWidth = 7;
  parameter int D2HRspFullWidth = D2HRspMaxWidth + D2HRspIntgWidth;
  parameter int DataMaxWidth    = 32;
  parameter int DataIntgWidth   = 7;
  parameter int DataFullWidth   = DataMaxWidth + DataIntgWidth;

  // Data that is returned upon an a TL-UL error belonging to an instruction fetch.
  // Note that this data will be returned with the correct bus integrity value.
  parameter logic [top_pkg::TL_DW-1:0] DataWhenInstrError = '0;
  // Data that is returned upon an a TL-UL error not belonging to an instruction fetch.
  // Note that this data will be returned with the correct bus integrity value.
  parameter logic [top_pkg::TL_DW-1:0] DataWhenError      = {top_pkg::TL_DW{1'b1}};

  typedef struct packed {
    logic [4:0]                 rsvd;
    prim_mubi_pkg::mubi4_t      instr_type;
    logic [H2DCmdIntgWidth-1:0] cmd_intg;
    logic [DataIntgWidth-1:0]   data_intg;
  } tl_a_user_t;

  parameter tl_a_user_t TL_A_USER_DEFAULT = '{
    rsvd: '0,
    instr_type: prim_mubi_pkg::MuBi4False,
    cmd_intg:  {H2DCmdIntgWidth{1'b1}},
    data_intg: {DataIntgWidth{1'b1}}
  };

  typedef struct packed {
    prim_mubi_pkg::mubi4_t        instr_type;
    logic   [top_pkg::TL_AW-1:0]  addr;
    tl_a_op_e                     opcode;
    logic  [top_pkg::TL_DBW-1:0]  mask;
  } tl_h2d_cmd_intg_t;

  typedef struct packed {
    logic                         a_valid;
    tl_a_op_e                     a_opcode;
    logic                  [2:0]  a_param;
    logic  [top_pkg::TL_SZW-1:0]  a_size;
    logic  [top_pkg::TL_AIW-1:0]  a_source;
    logic   [top_pkg::TL_AW-1:0]  a_address;
    logic  [top_pkg::TL_DBW-1:0]  a_mask;
    logic   [top_pkg::TL_DW-1:0]  a_data;
    tl_a_user_t                   a_user;

    logic                         d_ready;
  } tl_h2d_t;

  typedef struct packed {
    logic                         a_valid;
    tl_a_op_e                     a_opcode;
    logic                  [2:0]  a_param;
    logic  [top_pkg::TL_SZW64-1:0]  a_size;
    logic  [top_pkg::TL_AIW-1:0]  a_source;
    logic   [top_pkg::TL_AW-1:0]  a_address;
    logic  [top_pkg::TL_DBW64-1:0]  a_mask;
    logic   [top_pkg::TL_DW64-1:0]  a_data;
    tl_a_user_t                   a_user;

    logic                         d_ready;
  } tl_h2d_t64;

  // The choice of all 1's as the blanked value is deliberate.
  // It is assumed that most security features of the design are opt-in instead
  // of opt-out.
  // Given the opt-in nature, if a 0 were to propagate, the feature would be turned
  // off.  Whereas if a 1 were to propagate, it would either stay on or be turned on.
  // There is however no perfect value for this purpose.
  localparam logic [top_pkg::TL_DW-1:0] BlankedAData = {top_pkg::TL_DW{1'b1}};

  localparam tl_h2d_t TL_H2D_DEFAULT = '{
    d_ready:  1'b1,
    a_opcode: tl_a_op_e'('0),
    a_user:   TL_A_USER_DEFAULT,
    a_data:   BlankedAData,
    default:  '0
  };

  typedef struct packed {
    logic [D2HRspIntgWidth-1:0]    rsp_intg;
    logic [DataIntgWidth-1:0]      data_intg;
  } tl_d_user_t;

  parameter tl_d_user_t TL_D_USER_DEFAULT = '{
    rsp_intg: {D2HRspIntgWidth{1'b1}},
    data_intg: {DataIntgWidth{1'b1}}
  };

  typedef struct packed {
    logic                         d_valid;
    tl_d_op_e                     d_opcode;
    logic                  [2:0]  d_param;
    logic  [top_pkg::TL_SZW-1:0]  d_size;   // Bouncing back a_size
    logic  [top_pkg::TL_AIW-1:0]  d_source;
    logic  [top_pkg::TL_DIW-1:0]  d_sink;
    logic   [top_pkg::TL_DW-1:0]  d_data;
    tl_d_user_t                   d_user;
    logic                         d_error;

    logic                         a_ready;

  } tl_d2h_t;

  typedef struct packed {
    logic                         d_valid;
    tl_d_op_e                     d_opcode;
    logic                  [2:0]  d_param;
    logic  [top_pkg::TL_SZW64-1:0]  d_size;   // Bouncing back a_size
    logic  [top_pkg::TL_AIW-1:0]  d_source;
    logic  [top_pkg::TL_DIW-1:0]  d_sink;
    logic   [top_pkg::TL_DW64-1:0]  d_data;
    tl_d_user_t                   d_user;
    logic                         d_error;

    logic                         a_ready;

  } tl_d2h_t64;

  typedef struct packed {
    tl_d_op_e                     opcode;
    logic  [top_pkg::TL_SZW-1:0]  size;
    // Temporarily removed because source changes throughout the fabric
    // and thus cannot be used for end-to-end checking.
    // A different PR will propose a work-around (a hoaky one) to see if
    // it gets the job done.
    //logic  [top_pkg::TL_AIW-1:0]  source;
    logic                         error;
  } tl_d2h_rsp_intg_t;

  localparam tl_d2h_t TL_D2H_DEFAULT = '{
    a_ready:  1'b1,
    d_opcode: tl_d_op_e'('0),
    d_user:   TL_D_USER_DEFAULT,
    default:  '0
  };

  // Check user for unsupported values
  function automatic logic tl_a_user_chk(tl_a_user_t user);
    logic malformed_err;
    logic unused_user;
    unused_user = |user;
    malformed_err = prim_mubi_pkg::mubi4_test_invalid(user.instr_type);
    return malformed_err;
  endfunction // tl_a_user_chk

  // extract variables used for command checking
  function automatic tl_h2d_cmd_intg_t extract_h2d_cmd_intg(tl_h2d_t tl);
    tl_h2d_cmd_intg_t payload;
    logic unused_tlul;
    unused_tlul = ^tl;
    payload.addr = tl.a_address;
    payload.opcode = tl.a_opcode;
    payload.mask = tl.a_mask;
    payload.instr_type = tl.a_user.instr_type;
    return payload;
  endfunction // extract_h2d_payload

  // extract variables used for response checking
  function automatic tl_d2h_rsp_intg_t extract_d2h_rsp_intg(tl_d2h_t tl);
    tl_d2h_rsp_intg_t payload;
    logic unused_tlul;
    unused_tlul = ^tl;
    payload.opcode = tl.d_opcode;
    payload.size   = tl.d_size;
    //payload.source = tl.d_source;
    payload.error  = tl.d_error;
    return payload;
  endfunction // extract_d2h_rsp_intg

  // calculate ecc for command checking
  function automatic logic [H2DCmdIntgWidth-1:0] get_cmd_intg(tl_h2d_t tl);
    logic [H2DCmdIntgWidth-1:0] cmd_intg;
    logic [H2DCmdMaxWidth-1:0] unused_cmd_payload;
    tl_h2d_cmd_intg_t cmd;
    cmd = extract_h2d_cmd_intg(tl);
    {cmd_intg, unused_cmd_payload} =
        prim_secded_pkg::prim_secded_inv_64_57_enc(H2DCmdMaxWidth'(cmd));
   return cmd_intg;
  endfunction  // get_cmd_intg

  // calculate ecc for data checking
  function automatic logic [DataIntgWidth-1:0] get_data_intg(logic [top_pkg::TL_DW-1:0] data);
    logic [DataIntgWidth-1:0] data_intg;
    logic [top_pkg::TL_DW-1:0] unused_data;
    logic [DataIntgWidth + top_pkg::TL_DW - 1 : 0] enc_data;
    enc_data = prim_secded_pkg::prim_secded_inv_39_32_enc(data);
    data_intg = enc_data[DataIntgWidth + top_pkg::TL_DW - 1 : top_pkg::TL_DW];
    unused_data = enc_data[top_pkg::TL_DW - 1 : 0];
    return data_intg;
  endfunction  // get_data_intg

  // return inverted integrity for command payload
  function automatic logic [H2DCmdIntgWidth-1:0] get_bad_cmd_intg(tl_h2d_t tl);
    logic [H2DCmdIntgWidth-1:0] cmd_intg;
    cmd_intg = get_cmd_intg(tl);
    return ~cmd_intg;
  endfunction // get_bad_cmd_intg

  // return inverted integrity for data payload
  function automatic logic [H2DCmdIntgWidth-1:0] get_bad_data_intg(logic [top_pkg::TL_DW-1:0] data);
    logic [H2DCmdIntgWidth-1:0] data_intg;
    data_intg = get_data_intg(data);
    return ~data_intg;
  endfunction // get_bad_data_intg

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package otp_ctrl_pkg;

  import prim_util_pkg::vbits;
  import otp_ctrl_reg_pkg::*;

  ////////////////////////
  // General Parameters //
  ////////////////////////

  // Number of vendor-specific test CSR bits coming from and going to
  // the life cycle TAP registers.
  parameter int OtpTestCtrlWidth   = 32;
  parameter int OtpTestStatusWidth = 32;
  parameter int OtpTestVectWidth   = 8;

  // Width of entropy input
  parameter int EdnDataWidth = 64;

  parameter int NumPartWidth = vbits(NumPart);

  parameter int SwWindowAddrWidth = vbits(NumSwCfgWindowWords);

  // Background check timer LFSR width.
  parameter int LfsrWidth = 40;
  // The LFSR will be reseeded once LfsrUsageThreshold
  // values have been drawn from it.
  parameter int LfsrUsageThreshold = 16;

  // Redundantly encoded and complementary values are used to for signalling to the partition
  // controller FSMs and the DAI whether a partition is locked or not. Any other value than
  // "Mubi8Lo" is interpreted as "Locked" in those FSMs.
  typedef struct packed {
    prim_mubi_pkg::mubi8_t read_lock;
    prim_mubi_pkg::mubi8_t write_lock;
  } part_access_t;

  parameter int DaiCmdWidth = 3;
  typedef enum logic [DaiCmdWidth-1:0] {
    DaiRead   = 3'b001,
    DaiWrite  = 3'b010,
    DaiDigest = 3'b100
  } dai_cmd_e;

  parameter int DeviceIdWidth = 256;
  typedef logic [DeviceIdWidth-1:0] otp_device_id_t;

  parameter int ManufStateWidth = 256;
  typedef logic [ManufStateWidth-1:0] otp_manuf_state_t;

  //////////////////////////////////////
  // Typedefs for OTP Macro Interface //
  //////////////////////////////////////

  // OTP-macro specific
  parameter int OtpWidth         = 16;
  parameter int OtpAddrWidth     = OtpByteAddrWidth - $clog2(OtpWidth/8);
  parameter int OtpDepth         = 2**OtpAddrWidth;
  parameter int OtpSizeWidth     = 2; // Allows to transfer up to 4 native OTP words at once.
  parameter int OtpErrWidth      = 3;
  parameter int OtpPwrSeqWidth   = 2;
  parameter int OtpIfWidth       = 2**OtpSizeWidth*OtpWidth;
  // Number of Byte address bits to cut off in order to get the native OTP word address.
  parameter int OtpAddrShift     = OtpByteAddrWidth - OtpAddrWidth;

  typedef enum logic [OtpErrWidth-1:0] {
    NoError              = 3'h0,
    MacroError           = 3'h1,
    MacroEccCorrError    = 3'h2,
    MacroEccUncorrError  = 3'h3,
    MacroWriteBlankError = 3'h4,
    AccessError          = 3'h5,
    CheckFailError       = 3'h6,
    FsmStateError        = 3'h7
  } otp_err_e;

  /////////////////////////////////
  // Typedefs for OTP Scrambling //
  /////////////////////////////////

  parameter int ScrmblKeyWidth   = 128;
  parameter int ScrmblBlockWidth = 64;

  parameter int NumPresentRounds = 31;
  parameter int ScrmblBlockHalfWords = ScrmblBlockWidth / OtpWidth;

  typedef enum logic [2:0] {
    Decrypt,
    Encrypt,
    LoadShadow,
    Digest,
    DigestInit,
    DigestFinalize
  } otp_scrmbl_cmd_e;

  ///////////////////////////////
  // Typedefs for LC Interface //
  ///////////////////////////////

  // The tokens below are all hash post-images
  typedef struct packed {
    logic                            valid;
    logic                            error;
    // Use lc_state_t and lc_cnt_t here as very wide enumerations ( > 64 bits )
    // are not supported for virtual interfaces by Excelium yet
    // https://github.com/lowRISC/opentitan/issues/8884 (Cadence issue: cds_46570160)
    // The enumeration types lc_state_e and lc_cnt_e are still ok in other circumstances
    lc_ctrl_state_pkg::lc_state_t    state;
    lc_ctrl_state_pkg::lc_cnt_t      count;
    // This is set to "On" if the partition containing the
    // root secrets have been locked. In that case, the device
    // is considered "personalized".
    lc_ctrl_pkg::lc_tx_t             secrets_valid;
    // This is set to "On" if the partition containing the
    // test tokens has been locked.
    lc_ctrl_pkg::lc_tx_t             test_tokens_valid;
    lc_ctrl_state_pkg::lc_token_t    test_unlock_token;
    lc_ctrl_state_pkg::lc_token_t    test_exit_token;
    // This is set to "On" if the partition containing the
    // rma token has been locked.
    lc_ctrl_pkg::lc_tx_t             rma_token_valid;
    lc_ctrl_state_pkg::lc_token_t    rma_token;
  } otp_lc_data_t;

  // Default for dangling connection.
  // Note that we put the life cycle into
  // TEST_UNLOCKED0 by default such that top levels without
  // the OTP controller can still function.
  parameter otp_lc_data_t OTP_LC_DATA_DEFAULT = '{
    valid: 1'b1,
    error: 1'b0,
    state: lc_ctrl_state_pkg::LcStTestUnlocked0,
    count: lc_ctrl_state_pkg::LcCnt1,
    secrets_valid: lc_ctrl_pkg::Off,
    test_tokens_valid: lc_ctrl_pkg::Off,
    test_unlock_token: '0,
    test_exit_token: '0,
    rma_token_valid: lc_ctrl_pkg::Off,
    rma_token: '0
  };

  typedef struct packed {
    logic req;
    lc_ctrl_state_pkg::lc_state_e state;
    lc_ctrl_state_pkg::lc_cnt_e   count;
  } lc_otp_program_req_t;

  typedef struct packed {
    logic err;
    logic ack;
  } lc_otp_program_rsp_t;

  // RAW unlock token hashing request.
  typedef struct packed {
    logic req;
    lc_ctrl_state_pkg::lc_token_t token_input;
  } lc_otp_token_req_t;

  typedef struct packed {
    logic ack;
    lc_ctrl_state_pkg::lc_token_t hashed_token;
  } lc_otp_token_rsp_t;

  typedef struct packed {
    logic [OtpTestCtrlWidth-1:0] ctrl;
  } lc_otp_vendor_test_req_t;

  typedef struct packed {
    logic [OtpTestStatusWidth-1:0] status;
  } lc_otp_vendor_test_rsp_t;

  ////////////////////////////////
  // Typedefs for Key Broadcast //
  ////////////////////////////////

  parameter int FlashKeySeedWidth = 256;
  parameter int SramKeySeedWidth  = 128;
  parameter int KeyMgrKeyWidth    = 256;
  parameter int FlashKeyWidth     = 128;
  parameter int SramKeyWidth      = 128;
  parameter int SramNonceWidth    = 128;
  parameter int OtbnKeyWidth      = 128;
  parameter int OtbnNonceWidth    = 64;

  typedef logic [SramKeyWidth-1:0]   sram_key_t;
  typedef logic [SramNonceWidth-1:0] sram_nonce_t;
  typedef logic [OtbnKeyWidth-1:0]   otbn_key_t;
  typedef logic [OtbnNonceWidth-1:0] otbn_nonce_t;

  localparam int OtbnNonceSel  = OtbnNonceWidth / ScrmblBlockWidth;
  localparam int FlashNonceSel = FlashKeyWidth / ScrmblBlockWidth;
  localparam int SramNonceSel  = SramNonceWidth / ScrmblBlockWidth;

  // Get maximum nonce width
  localparam int NumNonceChunks =
    (OtbnNonceWidth > FlashKeyWidth) ?
    ((OtbnNonceWidth > SramNonceSel) ? OtbnNonceSel : SramNonceSel) :
    ((FlashKeyWidth > SramNonceSel)  ? FlashNonceSel  : SramNonceSel);

  typedef struct packed {
    logic valid;
    logic [KeyMgrKeyWidth-1:0] key_share0;
    logic [KeyMgrKeyWidth-1:0] key_share1;
  } otp_keymgr_key_t;

  parameter otp_keymgr_key_t OTP_KEYMGR_KEY_DEFAULT = '{
    valid: 1'b1,
    key_share0: 256'hefb7ea7ee90093cf4affd9aaa2d6c0ec446cfdf5f2d5a0bfd7e2d93edc63a102,
    key_share1: 256'h56d24a00181de99e0f690b447a8dde2a1ffb8bc306707107aa6e2410f15cfc37
  };

  typedef struct packed {
    logic data_req; // Requests static key for data scrambling.
    logic addr_req; // Requests static key for address scrambling.
  } flash_otp_key_req_t;

  typedef struct packed {
    logic req; // Requests ephemeral scrambling key and nonce.
  } sram_otp_key_req_t;

  typedef struct packed {
    logic req; // Requests ephemeral scrambling key and nonce.
  } otbn_otp_key_req_t;

  typedef struct packed {
    logic data_ack;                    // Ack for data key.
    logic addr_ack;                    // Ack for address key.
    logic [FlashKeyWidth-1:0] key;     // 128bit static scrambling key.
    logic [FlashKeyWidth-1:0] rand_key;
    logic seed_valid;                  // Set to 1 if the key seed has been provisioned and is
                                       // valid.
  } flash_otp_key_rsp_t;

  // Default for dangling connection
  parameter flash_otp_key_rsp_t FLASH_OTP_KEY_RSP_DEFAULT = '{
    data_ack: 1'b1,
    addr_ack: 1'b1,
    key: '0,
    rand_key: '0,
    seed_valid: 1'b1
  };

  typedef struct packed {
    logic        ack;        // Ack for key.
    sram_key_t   key;        // 128bit ephemeral scrambling key.
    sram_nonce_t nonce;      // 128bit nonce.
    logic        seed_valid; // Set to 1 if the key seed has been provisioned and is valid.
  } sram_otp_key_rsp_t;

  // Default for dangling connection
  parameter sram_otp_key_rsp_t SRAM_OTP_KEY_RSP_DEFAULT = '{
    ack: 1'b1,
    key: '0,
    nonce: '0,
    seed_valid: 1'b1
  };

  typedef struct packed {
    logic        ack;        // Ack for key.
    otbn_key_t   key;        // 128bit ephemeral scrambling key.
    otbn_nonce_t nonce;      // 256bit nonce.
    logic        seed_valid; // Set to 1 if the key seed has been provisioned and is valid.
  } otbn_otp_key_rsp_t;

  ////////////////////////////////
  // Power/Reset Ctrl Interface //
  ////////////////////////////////

  typedef struct packed {
    logic init;
  } pwr_otp_init_req_t;

  typedef struct packed {
    logic done;
  } pwr_otp_init_rsp_t;

  typedef struct packed {
    logic idle;
  } otp_pwr_state_t;


  ///////////////////
  // AST Interface //
  ///////////////////

  typedef struct packed {
    logic [OtpPwrSeqWidth-1:0] pwr_seq;
  } otp_ast_req_t;

  typedef struct packed {
    logic [OtpPwrSeqWidth-1:0] pwr_seq_h;
  } otp_ast_rsp_t;

  ///////////////////////////////////////////
  // Defaults for random netlist constants //
  ///////////////////////////////////////////

  // These LFSR parameters have been generated with
  // $ util/design/gen-lfsr-seed.py --width 40 --seed 4247488366
  typedef logic [LfsrWidth-1:0]                        lfsr_seed_t;
  typedef logic [LfsrWidth-1:0][$clog2(LfsrWidth)-1:0] lfsr_perm_t;
  localparam lfsr_seed_t RndCnstLfsrSeedDefault = 40'h453d28ea98;
  localparam lfsr_perm_t RndCnstLfsrPermDefault =
      240'h4235171482c225f79289b32181a0163a760355d3447063d16661e44c12a5;

  typedef struct packed {
    sram_key_t   key;
    sram_nonce_t nonce;
  } scrmbl_key_init_t;
  localparam scrmbl_key_init_t RndCnstScrmblKeyInitDefault =
      256'hcebeb96ffe0eced795f8b2cfe23c1e519e4fa08047a6bcfb811b04f0a479006e;

endpackage : otp_ctrl_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package csrng_reg_pkg;

  // Param list
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 7;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } cs_cmd_req_done;
    struct packed {
      logic        q;
    } cs_entropy_req;
    struct packed {
      logic        q;
    } cs_hw_inst_exc;
    struct packed {
      logic        q;
    } cs_fatal_err;
  } csrng_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } cs_cmd_req_done;
    struct packed {
      logic        q;
    } cs_entropy_req;
    struct packed {
      logic        q;
    } cs_hw_inst_exc;
    struct packed {
      logic        q;
    } cs_fatal_err;
  } csrng_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } cs_cmd_req_done;
    struct packed {
      logic        q;
      logic        qe;
    } cs_entropy_req;
    struct packed {
      logic        q;
      logic        qe;
    } cs_hw_inst_exc;
    struct packed {
      logic        q;
      logic        qe;
    } cs_fatal_err;
  } csrng_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_alert;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_alert;
  } csrng_reg2hw_alert_test_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } enable;
    struct packed {
      logic [3:0]  q;
    } sw_app_enable;
    struct packed {
      logic [3:0]  q;
    } read_int_state;
  } csrng_reg2hw_ctrl_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } csrng_reg2hw_cmd_req_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        re;
  } csrng_reg2hw_genbits_reg_t;

  typedef struct packed {
    logic [3:0]  q;
    logic        qe;
  } csrng_reg2hw_int_state_num_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        re;
  } csrng_reg2hw_int_state_val_reg_t;

  typedef struct packed {
    logic [4:0]  q;
    logic        qe;
  } csrng_reg2hw_err_code_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } cs_cmd_req_done;
    struct packed {
      logic        d;
      logic        de;
    } cs_entropy_req;
    struct packed {
      logic        d;
      logic        de;
    } cs_hw_inst_exc;
    struct packed {
      logic        d;
      logic        de;
    } cs_fatal_err;
  } csrng_hw2reg_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } cmd_rdy;
    struct packed {
      logic        d;
      logic        de;
    } cmd_sts;
  } csrng_hw2reg_sw_cmd_sts_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } genbits_vld;
    struct packed {
      logic        d;
    } genbits_fips;
  } csrng_hw2reg_genbits_vld_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } csrng_hw2reg_genbits_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } csrng_hw2reg_int_state_val_reg_t;

  typedef struct packed {
    logic [15:0] d;
    logic        de;
  } csrng_hw2reg_hw_exc_sts_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } enable_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } sw_app_enable_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } read_int_state_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } acmd_flag0_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } cs_bus_cmp_alert;
    struct packed {
      logic        d;
      logic        de;
    } cs_main_sm_alert;
  } csrng_hw2reg_recov_alert_sts_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } sfifo_cmd_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_genbits_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_cmdreq_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_rcstage_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_keyvrc_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_updreq_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_bencreq_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_bencack_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_pdata_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_final_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_gbencack_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_grcstage_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_ggenreq_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_gadstage_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_ggenbits_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_blkenc_err;
    struct packed {
      logic        d;
      logic        de;
    } cmd_stage_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } main_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } drbg_gen_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } drbg_updbe_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } drbg_updob_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } aes_cipher_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } cmd_gen_cnt_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_write_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_read_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_state_err;
  } csrng_hw2reg_err_code_reg_t;

  typedef struct packed {
    logic [7:0]  d;
    logic        de;
  } csrng_hw2reg_main_sm_state_reg_t;

  // Register -> HW type
  typedef struct packed {
    csrng_reg2hw_intr_state_reg_t intr_state; // [141:138]
    csrng_reg2hw_intr_enable_reg_t intr_enable; // [137:134]
    csrng_reg2hw_intr_test_reg_t intr_test; // [133:126]
    csrng_reg2hw_alert_test_reg_t alert_test; // [125:122]
    csrng_reg2hw_ctrl_reg_t ctrl; // [121:110]
    csrng_reg2hw_cmd_req_reg_t cmd_req; // [109:77]
    csrng_reg2hw_genbits_reg_t genbits; // [76:44]
    csrng_reg2hw_int_state_num_reg_t int_state_num; // [43:39]
    csrng_reg2hw_int_state_val_reg_t int_state_val; // [38:6]
    csrng_reg2hw_err_code_test_reg_t err_code_test; // [5:0]
  } csrng_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    csrng_hw2reg_intr_state_reg_t intr_state; // [167:160]
    csrng_hw2reg_sw_cmd_sts_reg_t sw_cmd_sts; // [159:156]
    csrng_hw2reg_genbits_vld_reg_t genbits_vld; // [155:154]
    csrng_hw2reg_genbits_reg_t genbits; // [153:122]
    csrng_hw2reg_int_state_val_reg_t int_state_val; // [121:90]
    csrng_hw2reg_hw_exc_sts_reg_t hw_exc_sts; // [89:73]
    csrng_hw2reg_recov_alert_sts_reg_t recov_alert_sts; // [72:61]
    csrng_hw2reg_err_code_reg_t err_code; // [60:9]
    csrng_hw2reg_main_sm_state_reg_t main_sm_state; // [8:0]
  } csrng_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] CSRNG_INTR_STATE_OFFSET = 7'h 0;
  parameter logic [BlockAw-1:0] CSRNG_INTR_ENABLE_OFFSET = 7'h 4;
  parameter logic [BlockAw-1:0] CSRNG_INTR_TEST_OFFSET = 7'h 8;
  parameter logic [BlockAw-1:0] CSRNG_ALERT_TEST_OFFSET = 7'h c;
  parameter logic [BlockAw-1:0] CSRNG_REGWEN_OFFSET = 7'h 10;
  parameter logic [BlockAw-1:0] CSRNG_CTRL_OFFSET = 7'h 14;
  parameter logic [BlockAw-1:0] CSRNG_CMD_REQ_OFFSET = 7'h 18;
  parameter logic [BlockAw-1:0] CSRNG_SW_CMD_STS_OFFSET = 7'h 1c;
  parameter logic [BlockAw-1:0] CSRNG_GENBITS_VLD_OFFSET = 7'h 20;
  parameter logic [BlockAw-1:0] CSRNG_GENBITS_OFFSET = 7'h 24;
  parameter logic [BlockAw-1:0] CSRNG_INT_STATE_NUM_OFFSET = 7'h 28;
  parameter logic [BlockAw-1:0] CSRNG_INT_STATE_VAL_OFFSET = 7'h 2c;
  parameter logic [BlockAw-1:0] CSRNG_HW_EXC_STS_OFFSET = 7'h 30;
  parameter logic [BlockAw-1:0] CSRNG_RECOV_ALERT_STS_OFFSET = 7'h 34;
  parameter logic [BlockAw-1:0] CSRNG_ERR_CODE_OFFSET = 7'h 38;
  parameter logic [BlockAw-1:0] CSRNG_ERR_CODE_TEST_OFFSET = 7'h 3c;
  parameter logic [BlockAw-1:0] CSRNG_MAIN_SM_STATE_OFFSET = 7'h 40;

  // Reset values for hwext registers and their fields
  parameter logic [3:0] CSRNG_INTR_TEST_RESVAL = 4'h 0;
  parameter logic [0:0] CSRNG_INTR_TEST_CS_CMD_REQ_DONE_RESVAL = 1'h 0;
  parameter logic [0:0] CSRNG_INTR_TEST_CS_ENTROPY_REQ_RESVAL = 1'h 0;
  parameter logic [0:0] CSRNG_INTR_TEST_CS_HW_INST_EXC_RESVAL = 1'h 0;
  parameter logic [0:0] CSRNG_INTR_TEST_CS_FATAL_ERR_RESVAL = 1'h 0;
  parameter logic [1:0] CSRNG_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] CSRNG_ALERT_TEST_RECOV_ALERT_RESVAL = 1'h 0;
  parameter logic [0:0] CSRNG_ALERT_TEST_FATAL_ALERT_RESVAL = 1'h 0;
  parameter logic [1:0] CSRNG_GENBITS_VLD_RESVAL = 2'h 0;
  parameter logic [31:0] CSRNG_GENBITS_RESVAL = 32'h 0;
  parameter logic [31:0] CSRNG_INT_STATE_VAL_RESVAL = 32'h 0;

  // Register index
  typedef enum int {
    CSRNG_INTR_STATE,
    CSRNG_INTR_ENABLE,
    CSRNG_INTR_TEST,
    CSRNG_ALERT_TEST,
    CSRNG_REGWEN,
    CSRNG_CTRL,
    CSRNG_CMD_REQ,
    CSRNG_SW_CMD_STS,
    CSRNG_GENBITS_VLD,
    CSRNG_GENBITS,
    CSRNG_INT_STATE_NUM,
    CSRNG_INT_STATE_VAL,
    CSRNG_HW_EXC_STS,
    CSRNG_RECOV_ALERT_STS,
    CSRNG_ERR_CODE,
    CSRNG_ERR_CODE_TEST,
    CSRNG_MAIN_SM_STATE
  } csrng_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] CSRNG_PERMIT [17] = '{
    4'b 0001, // index[ 0] CSRNG_INTR_STATE
    4'b 0001, // index[ 1] CSRNG_INTR_ENABLE
    4'b 0001, // index[ 2] CSRNG_INTR_TEST
    4'b 0001, // index[ 3] CSRNG_ALERT_TEST
    4'b 0001, // index[ 4] CSRNG_REGWEN
    4'b 0011, // index[ 5] CSRNG_CTRL
    4'b 1111, // index[ 6] CSRNG_CMD_REQ
    4'b 0001, // index[ 7] CSRNG_SW_CMD_STS
    4'b 0001, // index[ 8] CSRNG_GENBITS_VLD
    4'b 1111, // index[ 9] CSRNG_GENBITS
    4'b 0001, // index[10] CSRNG_INT_STATE_NUM
    4'b 1111, // index[11] CSRNG_INT_STATE_VAL
    4'b 0011, // index[12] CSRNG_HW_EXC_STS
    4'b 0011, // index[13] CSRNG_RECOV_ALERT_STS
    4'b 1111, // index[14] CSRNG_ERR_CODE
    4'b 0001, // index[15] CSRNG_ERR_CODE_TEST
    4'b 0001  // index[16] CSRNG_MAIN_SM_STATE
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package csrng_pkg;

  //-------------------------
  // Application Interfaces
  //-------------------------

  parameter int unsigned GENBITS_BUS_WIDTH = 128;
  parameter int unsigned CSRNG_CMD_WIDTH = 32;
  parameter int unsigned FIPS_GENBITS_BUS_WIDTH = entropy_src_pkg::FIPS_BUS_WIDTH +
                         GENBITS_BUS_WIDTH;
  parameter int unsigned MainSmStateWidth = 8;

  // instantiation interface
  typedef struct packed {
    logic                       csrng_req_valid;
    logic [CSRNG_CMD_WIDTH-1:0] csrng_req_bus;
    logic                       genbits_ready;
  } csrng_req_t;

  typedef struct packed {
    logic                         csrng_req_ready;
    logic                         csrng_rsp_ack;
    logic                         csrng_rsp_sts;
    logic                         genbits_valid;
    logic                         genbits_fips;
    logic [GENBITS_BUS_WIDTH-1:0] genbits_bus;
  } csrng_rsp_t;

  parameter csrng_req_t CSRNG_REQ_DEFAULT = '{default: '0};
  parameter csrng_rsp_t CSRNG_RSP_DEFAULT = '{default: '0};

  typedef enum logic [2:0] {
    INV  = 3'h0,
    INS  = 3'h1,
    RES  = 3'h2,
    GEN  = 3'h3,
    UPD  = 3'h4,
    UNI  = 3'h5,
    GENB = 3'h6,
    GENU = 3'h7
  } acmd_e;


  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 15 -n 8 \
  //      -s 1300573258 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||| (32.38%)
  //  4: |||||||||||||||||||| (35.24%)
  //  5: |||||||| (15.24%)
  //  6: |||||| (11.43%)
  //  7: ||| (5.71%)
  //  8: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 7
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 7
  //
  typedef    enum logic [MainSmStateWidth-1:0] {
    MainSmIdle          = 8'b01001110, // idle
    MainSmParseCmd      = 8'b10111011, // parse the cmd
    MainSmInstantPrep   = 8'b11000001, // instantiate prep
    MainSmInstantReq    = 8'b01010100, // instantiate request (takes adata or entropy)
    MainSmReseedPrep    = 8'b11011101, // reseed prep
    MainSmReseedReq     = 8'b01011011, // reseed request (takes adata and entropy and Key,V,RC)
    MainSmGeneratePrep  = 8'b11101111, // generate request (takes adata? and Key,V,RC)
    MainSmGenerateReq   = 8'b00100100, // generate request (takes adata? and Key,V,RC)
    MainSmUpdatePrep    = 8'b00110001, // update prep
    MainSmUpdateReq     = 8'b10010000, // update request (takes adata and Key,V,RC)
    MainSmUninstantPrep = 8'b11110110, // uninstantiate prep
    MainSmUninstantReq  = 8'b01100011, // uninstantiate request
    MainSmClrAData      = 8'b00000010, // clear out the additional data packer fifo
    MainSmCmdCompWait   = 8'b10111100, // wait for command to complete
    MainSmError         = 8'b01111000  // error state, results in fatal alert
  } main_sm_state_e;

  parameter int CsKeymgrDivWidth = 384;
  typedef logic [CsKeymgrDivWidth-1:0] cs_keymgr_div_t;

endpackage : csrng_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package prim_alert_pkg;

  typedef struct packed {
    logic alert_p;
    logic alert_n;
  } alert_tx_t;

  typedef struct packed {
    logic ping_p;
    logic ping_n;
    logic ack_p;
    logic ack_n;
  } alert_rx_t;

  parameter alert_tx_t ALERT_TX_DEFAULT = '{alert_p:  1'b0,
                                            alert_n:  1'b1};

  parameter alert_rx_t ALERT_RX_DEFAULT = '{ping_p: 1'b0,
                                            ping_n: 1'b1,
                                            ack_p: 1'b0,
                                            ack_n: 1'b1};

endpackage : prim_alert_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// The alert receiver primitive decodes alerts that have been differentially
// encoded and transmitted via a handshake protocol on alert_p/n and
// ack_p/n. In case an alert handshake is initiated, the output alert_o will
// immediately be asserted (even before completion of the handshake).
//
// In case the differential input is not correctly encoded, this module will
// raise an error by asserting integ_fail_o.
//
// Further, the module supports ping testing of the alert diff pair. In order to
// initiate a ping test, ping_req_i shall be set to 1'b1 until ping_ok_o is
// asserted for one cycle. The signal may be de-asserted (e.g. after a long)
// timeout period. However note that all ping responses that come in after
// deasserting ping_req_i will be treated as native alerts.
//
// The protocol works in both asynchronous and synchronous cases. In the
// asynchronous case, the parameter AsyncOn must be set to 1'b1 in order to
// instantiate additional synchronization logic. Further, it must be ensured
// that the timing skew between all diff pairs is smaller than the shortest
// clock period of the involved clocks.
//
// Note that in case of synchronous operation, alerts on the diffpair are
// decoded combinationally and forwarded on alert_o within the same cycle.
//
// See also: prim_alert_sender, prim_diff_decode, alert_handler

`include "prim_assert.sv"

module prim_alert_receiver
  import prim_alert_pkg::*;
  import prim_mubi_pkg::mubi4_t;
#(
  // enables additional synchronization logic
  parameter bit AsyncOn = 1'b0
) (
  input             clk_i,
  input             rst_ni,
  // if set to lc_ctrl_pkg::On, this triggers the in-band alert channel
  // reset, which resets both the sender and receiver FSMs into IDLE.
  input mubi4_t     init_trig_i,
  // this triggers a ping test. keep asserted
  // until ping_ok_o is asserted.
  input             ping_req_i,
  output logic      ping_ok_o,
  // asserted if signal integrity issue detected
  output logic      integ_fail_o,
  // alert output (pulsed high) if a handshake is initiated
  // on alert_p/n and no ping request is outstanding
  output logic      alert_o,
  // ping input diff pair and ack diff pair
  output alert_rx_t alert_rx_o,
  // alert output diff pair
  input alert_tx_t  alert_tx_i
);

  import prim_mubi_pkg::mubi4_test_true_strict;

  /////////////////////////////////
  // decode differential signals //
  /////////////////////////////////
  logic alert_level, alert_sigint, alert_p, alert_n;

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_buf #(
    .Width(2)
  ) u_prim_buf_in (
    .in_i({alert_tx_i.alert_n,
           alert_tx_i.alert_p}),
    .out_o({alert_n,
            alert_p})
  );

  prim_diff_decode #(
    .AsyncOn(AsyncOn)
  ) u_decode_alert (
    .clk_i,
    .rst_ni,
    .diff_pi  ( alert_p            ),
    .diff_ni  ( alert_n            ),
    .level_o  ( alert_level        ),
    .rise_o   (                    ),
    .fall_o   (                    ),
    .event_o  (                    ),
    .sigint_o ( alert_sigint       )
  );

  /////////////////////////////////////////////////////
  //  main protocol FSM that drives the diff outputs //
  /////////////////////////////////////////////////////
  typedef enum logic [2:0] {Idle, HsAckWait, Pause0, Pause1, InitReq, InitAckWait} state_e;
  state_e state_d, state_q;
  logic ping_rise;
  logic ping_tog_pd, ping_tog_pq, ping_tog_dn, ping_tog_nq;
  logic ack_pd, ack_pq, ack_dn, ack_nq;
  logic ping_req_d, ping_req_q;
  logic ping_pending_d, ping_pending_q;
  logic send_init;
  logic send_ping;

  // signal ping request upon positive transition on ping_req_i
  // signalling is performed by a level change event on the diff output
  assign ping_req_d  = ping_req_i;
  assign ping_rise   = ping_req_d && !ping_req_q;
  assign ping_tog_pd = (send_init) ? 1'b0         :
                       (send_ping) ? ~ping_tog_pq : ping_tog_pq;

  // in-band reset is performed by sending out an integrity error on purpose.
  assign ack_dn      = (send_init) ? ack_pd : ~ack_pd;
  assign ping_tog_dn = ~ping_tog_pd;

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_flop #(
    .Width     (2),
    .ResetValue(2'b10)
  ) u_prim_generic_flop_ack (
    .clk_i,
    .rst_ni,
    .d_i({ack_dn,
          ack_pd}),
    .q_o({ack_nq,
          ack_pq})
  );

  prim_sec_anchor_flop #(
    .Width     (2),
    .ResetValue(2'b10)
  ) u_prim_generic_flop_ping (
    .clk_i,
    .rst_ni,
    .d_i({ping_tog_dn,
          ping_tog_pd}),
    .q_o({ping_tog_nq,
          ping_tog_pq})
  );

  // the ping pending signal is used in the FSM to distinguish whether the
  // incoming handshake shall be treated as an alert or a ping response.
  // it is important that this is only set on a rising ping_en level change, since
  // otherwise the ping enable signal could be abused to "mask" all native alerts
  // as ping responses by constantly tying it to 1.
  assign ping_pending_d = ping_rise | ((~ping_ok_o) & ping_req_i & ping_pending_q);

  // diff pair outputs
  assign alert_rx_o.ack_p = ack_pq;
  assign alert_rx_o.ack_n = ack_nq;

  assign alert_rx_o.ping_p = ping_tog_pq;
  assign alert_rx_o.ping_n = ping_tog_nq;

  // this FSM receives the four phase handshakes from the alert receiver
  // note that the latency of the alert_p/n input diff pair is at least one
  // cycle until it enters the receiver FSM. the same holds for the ack_* diff
  // pair outputs.
  always_comb begin : p_fsm
    // default
    state_d      = state_q;
    ack_pd       = 1'b0;
    ping_ok_o    = 1'b0;
    integ_fail_o = 1'b0;
    alert_o      = 1'b0;
    send_init    = 1'b0;
    // by default, a ping request leads to a toogle on the differential ping pair
    send_ping    = ping_rise;

    unique case (state_q)
      Idle: begin
        // wait for handshake to be initiated
        if (alert_level) begin
          state_d = HsAckWait;
          ack_pd  = 1'b1;
          // signal either an alert or ping received on the output
          if (ping_pending_q) begin
            ping_ok_o = 1'b1;
          end else begin
            alert_o   = 1'b1;
          end
        end
      end
      // waiting for deassertion of alert to complete HS
      HsAckWait: begin
        if (!alert_level) begin
          state_d  = Pause0;
        end else begin
          ack_pd = 1'b1;
        end
      end
      // pause cycles between back-to-back handshakes
      Pause0: state_d = Pause1;
      Pause1: state_d = Idle;
      // this state is only reached if an in-band reset is
      // requested via the low-power logic.
      InitReq: begin
        // we deliberately place a sigint error on the ack and ping lines in this case.
        send_init = 1'b1;
        // suppress any toggles on the ping line while we are in the init phase.
        send_ping = 1'b0;
        // As long as init req is asserted, we remain in this state and acknowledge all incoming
        // ping requests. As soon as the init request is dropped however, ping requests are not
        // acked anymore such that the ping mechanism can also flag alert channels that got stuck
        // in the initialization sequence.
        if (mubi4_test_true_strict(init_trig_i)) begin
          ping_ok_o = ping_pending_q;
        // the sender will respond to the sigint error above with a sigint error on the alert lines.
        // hence we treat the alert_sigint like an acknowledgement in this case.
        end else if (alert_sigint) begin
          state_d = InitAckWait;
        end
      end
      // We get here if the sender has responded with alert_sigint, and init_trig_i==lc_ctrl_pkg::On
      // has been deasserted. At this point, we need to wait for the alert_sigint to drop again
      // before resuming normal operation.
      InitAckWait: begin
        // suppress any toggles on the ping line while we are in the init phase.
        send_ping = 1'b0;
        if (!alert_sigint) begin
          state_d = Pause0;
          // If we get a ping request in this cycle, or if we realize that there is an unhandled
          // ping request that came in during initialization (but after init_trig_i has been
          // deasserted), we signal this to the alert sender by toggling the request line.
          send_ping = ping_rise || ping_pending_q;
        end
      end
      default: state_d = Idle;
    endcase

    // once the initialization sequence has been triggered,
    // overrides are not allowed anymore until the initialization has been completed.
    if (!(state_q inside {InitReq, InitAckWait})) begin
      // in this case, abort and jump into the initialization sequence
      if (mubi4_test_true_strict(init_trig_i)) begin
        state_d      = InitReq;
        ack_pd       = 1'b0;
        ping_ok_o    = 1'b0;
        integ_fail_o = 1'b0;
        alert_o      = 1'b0;
        send_init    = 1'b1;
      // if we're not busy with an init request, we clamp down all outputs
      // and indicate an integrity failure.
      end else if (alert_sigint) begin
        state_d      = Idle;
        ack_pd       = 1'b0;
        ping_ok_o    = 1'b0;
        integ_fail_o = 1'b1;
        alert_o      = 1'b0;
      end
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_reg
    if (!rst_ni) begin
      // Reset into the init request so that an alert handler reset implicitly
      // triggers an in-band reset of all alert channels.
      state_q        <= InitReq;
      ping_req_q     <= 1'b0;
      ping_pending_q <= 1'b0;
    end else begin
      state_q        <= state_d;
      ping_req_q     <= ping_req_d;
      ping_pending_q <= ping_pending_d;
    end
  end


  ////////////////
  // assertions //
  ////////////////

`ifdef INC_ASSERT
  import prim_mubi_pkg::mubi4_test_false_loose;
`endif

  // check whether all outputs have a good known state after reset
  `ASSERT_KNOWN(PingOkKnownO_A, ping_ok_o)
  `ASSERT_KNOWN(IntegFailKnownO_A, integ_fail_o)
  `ASSERT_KNOWN(AlertKnownO_A, alert_o)
  `ASSERT_KNOWN(PingPKnownO_A, alert_rx_o)

  // check encoding of outgoing diffpairs. note that during init, the outgoing diffpairs are
  // supposed to be incorrectly encoded on purpose.
  // shift sequence two cycles to the right to avoid reset effects.
  `ASSERT(PingDiffOk_A, alert_rx_o.ping_p ^ alert_rx_o.ping_n)
  `ASSERT(AckDiffOk_A, ##2 $past(send_init) ^ alert_rx_o.ack_p ^ alert_rx_o.ack_n)
  `ASSERT(InitReq_A, mubi4_test_true_strict(init_trig_i) &&
          !(state_q inside {InitReq, InitAckWait}) |=> send_init)

  // ping request at input -> need to see encoded ping request
  `ASSERT(PingRequest0_A, ##1 $rose(ping_req_i) && !state_q inside {InitReq, InitAckWait}
      |=> $changed(alert_rx_o.ping_p))
  // ping response implies it has been requested
  `ASSERT(PingResponse0_A, ping_ok_o |-> ping_pending_q)
  // correctly latch ping request
  `ASSERT(PingPending_A, ##1 $rose(ping_req_i) |=> ping_pending_q)

  if (AsyncOn) begin : gen_async_assert
    // signal integrity check propagation
    `ASSERT(SigInt_A,
        alert_tx_i.alert_p == alert_tx_i.alert_n [*2] ##2
        !(state_q inside {InitReq, InitAckWait}) &&
        mubi4_test_false_loose(init_trig_i)
        |->
        ##[0:1] integ_fail_o)
    `ASSERT(PingResponse1_A,
        ##1 $rose(alert_tx_i.alert_p) &&
        (alert_tx_i.alert_p ^ alert_tx_i.alert_n) ##2
        state_q == Idle && ping_pending_q
        |->
        ##[0:1] ping_ok_o,
        clk_i, !rst_ni || integ_fail_o || mubi4_test_true_strict(init_trig_i))
    // alert
    `ASSERT(Alert_A,
        ##1 $rose(alert_tx_i.alert_p) &&
        (alert_tx_i.alert_p ^ alert_tx_i.alert_n) ##2
        state_q == Idle &&
        !ping_pending_q
        |->
        ##[0:1] alert_o,
        clk_i, !rst_ni || integ_fail_o || mubi4_test_true_strict(init_trig_i))
  end else begin : gen_sync_assert
    // signal integrity check propagation
    `ASSERT(SigInt_A,
        alert_tx_i.alert_p == alert_tx_i.alert_n &&
        !(state_q inside {InitReq, InitAckWait}) &&
        mubi4_test_false_loose(init_trig_i)
        |->
        integ_fail_o)
    // ping response
    `ASSERT(PingResponse1_A,
        ##1 $rose(alert_tx_i.alert_p) &&
        state_q == Idle &&
        ping_pending_q
        |->
        ping_ok_o,
        clk_i, !rst_ni || integ_fail_o || mubi4_test_true_strict(init_trig_i))
    // alert
    `ASSERT(Alert_A,
        ##1 $rose(alert_tx_i.alert_p) &&
        state_q == Idle &&
        !ping_pending_q
        |->
        alert_o,
        clk_i, !rst_ni || integ_fail_o || mubi4_test_true_strict(init_trig_i))
  end

  // check in-band init request is always accepted
  `ASSERT(InBandInitRequest_A,
      mubi4_test_true_strict(init_trig_i) &&
      state_q != InitAckWait
      |=>
      state_q == InitReq)
  // check in-band init sequence moves FSM into IDLE state
  `ASSERT(InBandInitSequence_A,
      (state_q == InitReq &&
      mubi4_test_true_strict(init_trig_i)) ##1
      (alert_sigint &&
      mubi4_test_false_loose(init_trig_i)) [*1:$] ##1
      (!alert_sigint &&
      mubi4_test_false_loose(init_trig_i)) [*3]
      |=>
      state_q == Idle)
  // check there are no spurious alerts during init
  `ASSERT(NoSpuriousAlertsDuringInit_A,
      mubi4_test_true_strict(init_trig_i) ||
      (state_q inside {InitReq, InitAckWait})
      |->
      !alert_o)
  // check that there are no spurious ping OKs
  `ASSERT(NoSpuriousPingOksDuringInit_A,
      (mubi4_test_true_strict(init_trig_i) ||
      (state_q inside {InitReq, InitAckWait})) &&
      !ping_pending_q
      |->
      !ping_ok_o)
  // check ping request is bypassed when in init state
  `ASSERT(PingOkBypassDuringInit_A,
      $rose(ping_req_i) ##1
      state_q == InitReq &&
      mubi4_test_true_strict(init_trig_i)
      |->
      ping_ok_o)

endmodule : prim_alert_receiver


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// The alert sender primitive module differentially encodes and transmits an
// alert signal to the prim_alert_receiver module. An alert will be signalled
// by a full handshake on alert_p/n and ack_p/n. The alert_req_i signal may
// be continuously asserted, in which case the alert signalling handshake
// will be repeatedly initiated.
//
// The alert_req_i signal may also be used as part of req/ack. The parent module
// can keep alert_req_i asserted until it has been ack'd (transferred to the alert
// receiver).  The parent module is not required to use this.
//
// In case the alert sender parameter IsFatal is set to 1, an incoming alert
// alert_req_i is latched in a local register until the next reset, causing the
// alert sender to behave as if alert_req_i were continously asserted.
// The alert_state_o output reflects the state of this internal latching register.
//
// The alert sender also exposes an alert test input, which can be used to trigger
// single alert handshakes. This input behaves exactly the same way as the
// alert_req_i input with IsFatal set to 0. Test alerts do not cause alert_ack_o
// to be asserted, nor are they latched until reset (regardless of the value of the
// IsFatal parameter).
//
// Further, this module supports in-band ping testing, which means that a level
// change on the ping_p/n diff pair will result in a full-handshake response
// on alert_p/n and ack_p/n.
//
// The protocol works in both asynchronous and synchronous cases. In the
// asynchronous case, the parameter AsyncOn must be set to 1'b1 in order to
// instantiate additional synchronization logic. Further, it must be ensured
// that the timing skew between all diff pairs is smaller than the shortest
// clock period of the involved clocks.
//
// Incorrectly encoded diff inputs can be detected and will be signalled
// to the receiver by placing an inconsistent diff value on the differential
// output (and continuously toggling it).
//
// See also: prim_alert_receiver, prim_diff_decode, alert_handler

`include "prim_assert.sv"

module prim_alert_sender
  import prim_alert_pkg::*;
#(
  // enables additional synchronization logic
  parameter bit AsyncOn = 1'b1,
  // alert sender will latch the incoming alert event permanently and
  // keep on sending alert events until the next reset.
  parameter bit IsFatal = 1'b0
) (
  input             clk_i,
  input             rst_ni,
  // alert test trigger (this will never be latched, even if IsFatal == 1)
  input             alert_test_i,
  // native alert from the peripheral
  input             alert_req_i,
  output logic      alert_ack_o,
  // state of the alert latching register
  output logic      alert_state_o,
  // ping input diff pair and ack diff pair
  input alert_rx_t  alert_rx_i,
  // alert output diff pair
  output alert_tx_t alert_tx_o
);


  /////////////////////////////////
  // decode differential signals //
  /////////////////////////////////
  logic ping_sigint, ping_event, ping_n, ping_p;

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_buf #(
    .Width(2)
  ) u_prim_buf_ping (
    .in_i({alert_rx_i.ping_n,
           alert_rx_i.ping_p}),
    .out_o({ping_n,
            ping_p})
  );

  prim_diff_decode #(
    .AsyncOn(AsyncOn)
  ) u_decode_ping (
    .clk_i,
    .rst_ni,
    .diff_pi  ( ping_p      ),
    .diff_ni  ( ping_n      ),
    .level_o  (             ),
    .rise_o   (             ),
    .fall_o   (             ),
    .event_o  ( ping_event  ),
    .sigint_o ( ping_sigint )
  );

  logic ack_sigint, ack_level, ack_n, ack_p;

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_buf #(
    .Width(2)
  ) u_prim_buf_ack (
    .in_i({alert_rx_i.ack_n,
           alert_rx_i.ack_p}),
    .out_o({ack_n,
            ack_p})
  );

  prim_diff_decode #(
    .AsyncOn(AsyncOn)
  ) u_decode_ack (
    .clk_i,
    .rst_ni,
    .diff_pi  ( ack_p      ),
    .diff_ni  ( ack_n      ),
    .level_o  ( ack_level  ),
    .rise_o   (            ),
    .fall_o   (            ),
    .event_o  (            ),
    .sigint_o ( ack_sigint )
  );


  ///////////////////////////////////////////////////
  // main protocol FSM that drives the diff output //
  ///////////////////////////////////////////////////
  typedef enum logic [2:0] {
    Idle,
    AlertHsPhase1,
    AlertHsPhase2,
    PingHsPhase1,
    PingHsPhase2,
    Pause0,
    Pause1
    } state_e;
  state_e state_d, state_q;
  logic alert_pq, alert_nq, alert_pd, alert_nd;
  logic sigint_detected;

  assign sigint_detected = ack_sigint | ping_sigint;


  // diff pair output
  assign alert_tx_o.alert_p = alert_pq;
  assign alert_tx_o.alert_n = alert_nq;

  // alert and ping set regs
  logic alert_set_d, alert_set_q, alert_clr;
  logic alert_test_set_d, alert_test_set_q;
  logic ping_set_d, ping_set_q, ping_clr;
  logic alert_req_trigger, alert_test_trigger, ping_trigger;

  // if handshake is ongoing, capture additional alert requests.
  logic alert_req;
  prim_sec_anchor_buf #(
    .Width(1)
  ) u_prim_buf_in_req (
    .in_i(alert_req_i),
    .out_o(alert_req)
  );

  assign alert_req_trigger = alert_req | alert_set_q;
  if (IsFatal) begin : gen_fatal
    assign alert_set_d = alert_req_trigger;
  end else begin : gen_recov
    assign alert_set_d = (alert_clr) ? 1'b0 : alert_req_trigger;
  end

  // the alert test request is always cleared.
  assign alert_test_trigger = alert_test_i | alert_test_set_q;
  assign alert_test_set_d = (alert_clr) ? 1'b0 : alert_test_trigger;

  logic alert_trigger;
  assign alert_trigger = alert_req_trigger | alert_test_trigger;

  assign ping_trigger = ping_set_q | ping_event;
  assign ping_set_d  = (ping_clr) ? 1'b0 : ping_trigger;


  // alert event acknowledge and state (not affected by alert_test_i)
  assign alert_ack_o = alert_clr & alert_set_q;
  assign alert_state_o = alert_set_q;

  // this FSM performs a full four phase handshake upon a ping or alert trigger.
  // note that the latency of the alert_p/n diff pair is at least one cycle
  // until it enters the receiver FSM. the same holds for the ack_* diff pair
  // input. in case a signal integrity issue is detected, the FSM bails out,
  // sets the alert_p/n diff pair to the same value and toggles it in order to
  // signal that condition over to the receiver.
  always_comb begin : p_fsm
    // default
    state_d   = state_q;
    alert_pd  = 1'b0;
    alert_nd  = 1'b1;
    ping_clr  = 1'b0;
    alert_clr = 1'b0;

    unique case (state_q)
      Idle: begin
        // alert always takes precedence
        if (alert_trigger || ping_trigger) begin
          state_d = (alert_trigger) ? AlertHsPhase1 : PingHsPhase1;
          alert_pd = 1'b1;
          alert_nd = 1'b0;
        end
      end
      // waiting for ack from receiver
      AlertHsPhase1: begin
        if (ack_level) begin
          state_d  = AlertHsPhase2;
        end else begin
          alert_pd = 1'b1;
          alert_nd = 1'b0;
        end
      end
      // wait for deassertion of ack
      AlertHsPhase2: begin
        if (!ack_level) begin
          state_d = Pause0;
          alert_clr = 1'b1;
        end
      end
      // waiting for ack from receiver
      PingHsPhase1: begin
        if (ack_level) begin
          state_d  = PingHsPhase2;
        end else begin
          alert_pd = 1'b1;
          alert_nd = 1'b0;
        end
      end
      // wait for deassertion of ack
      PingHsPhase2: begin
        if (!ack_level) begin
          ping_clr = 1'b1;
          state_d = Pause0;
        end
      end
      // pause cycles between back-to-back handshakes
      Pause0: begin
        state_d = Pause1;
      end
      // clear and ack alert request if it was set
      Pause1: begin
        state_d = Idle;
      end
      // catch parasitic states
      default : state_d = Idle;
    endcase

    // we have a signal integrity issue at one of the incoming diff pairs. this condition is
    // signalled by setting the output diffpair to zero. If the sigint has disappeared, we clear
    // the ping request state of this sender and go back to idle.
    if (sigint_detected) begin
      state_d   = Idle;
      alert_pd  = 1'b0;
      alert_nd  = 1'b0;
      ping_clr  = 1'b1;
      alert_clr = 1'b0;
    end
  end

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_flop #(
    .Width     (2),
    .ResetValue(2'b10)
  ) u_prim_flop_alert (
    .clk_i,
    .rst_ni,
    .d_i({alert_nd, alert_pd}),
    .q_o({alert_nq, alert_pq})
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_reg
    if (!rst_ni) begin
      state_q          <= Idle;
      alert_set_q      <= 1'b0;
      alert_test_set_q <= 1'b0;
      ping_set_q       <= 1'b0;
    end else begin
      state_q          <= state_d;
      alert_set_q      <= alert_set_d;
      alert_test_set_q <= alert_test_set_d;
      ping_set_q       <= ping_set_d;
    end
  end


  ////////////////
  // assertions //
  ////////////////

// however, since we use sequence constructs below, we need to wrap the entire block again.
// typically, the ASSERT macros already contain this INC_ASSERT macro.
`ifdef INC_ASSERT
  // check whether all outputs have a good known state after reset
  `ASSERT_KNOWN(AlertPKnownO_A, alert_tx_o)

  if (AsyncOn) begin : gen_async_assert
    sequence PingSigInt_S;
      alert_rx_i.ping_p == alert_rx_i.ping_n [*2];
    endsequence
    sequence AckSigInt_S;
      alert_rx_i.ping_p == alert_rx_i.ping_n [*2];
    endsequence

  `ifndef FPV_ALERT_NO_SIGINT_ERR
    // check propagation of sigint issues to output within three cycles, or four due to CDC
    // shift sequence to the right to avoid reset effects.
    `ASSERT(SigIntPing_A, ##1 PingSigInt_S |->
        ##[3:4] alert_tx_o.alert_p == alert_tx_o.alert_n)
    `ASSERT(SigIntAck_A, ##1 AckSigInt_S |->
        ##[3:4] alert_tx_o.alert_p == alert_tx_o.alert_n)
  `endif

    // Test in-band FSM reset request (via signal integrity error)
    `ASSERT(InBandInitFsm_A, PingSigInt_S or AckSigInt_S |-> ##[3:4] state_q == Idle)
    `ASSERT(InBandInitPing_A, PingSigInt_S or AckSigInt_S |-> ##[3:4] !ping_set_q)
    // output must be driven diff unless sigint issue detected
    `ASSERT(DiffEncoding_A, (alert_rx_i.ack_p ^ alert_rx_i.ack_n) &&
        (alert_rx_i.ping_p ^ alert_rx_i.ping_n) |->
        ##[3:5] alert_tx_o.alert_p ^ alert_tx_o.alert_n)

    // handshakes can take indefinite time if blocked due to sigint on outgoing
    // lines (which is not visible here). thus, we only check whether the
    // handshake is correctly initiated and defer the full handshake checking to the testbench.
    `ASSERT(PingHs_A, ##1 $changed(alert_rx_i.ping_p) &&
        (alert_rx_i.ping_p ^ alert_rx_i.ping_n) ##2 state_q == Idle |=>
        ##[0:1] $rose(alert_tx_o.alert_p), clk_i,
        !rst_ni || (alert_tx_o.alert_p == alert_tx_o.alert_n))
  end else begin : gen_sync_assert
    sequence PingSigInt_S;
      alert_rx_i.ping_p == alert_rx_i.ping_n;
    endsequence
    sequence AckSigInt_S;
      alert_rx_i.ping_p == alert_rx_i.ping_n;
    endsequence

  `ifndef FPV_ALERT_NO_SIGINT_ERR
    // check propagation of sigint issues to output within one cycle
    `ASSERT(SigIntPing_A, PingSigInt_S |=>
        alert_tx_o.alert_p == alert_tx_o.alert_n)
    `ASSERT(SigIntAck_A,  AckSigInt_S |=>
        alert_tx_o.alert_p == alert_tx_o.alert_n)
  `endif

    // Test in-band FSM reset request (via signal integrity error)
    `ASSERT(InBandInitFsm_A, PingSigInt_S or AckSigInt_S |=> state_q == Idle)
    `ASSERT(InBandInitPing_A, PingSigInt_S or AckSigInt_S |=> !ping_set_q)
    // output must be driven diff unless sigint issue detected
    `ASSERT(DiffEncoding_A, (alert_rx_i.ack_p ^ alert_rx_i.ack_n) &&
        (alert_rx_i.ping_p ^ alert_rx_i.ping_n) |=> alert_tx_o.alert_p ^ alert_tx_o.alert_n)
    // handshakes can take indefinite time if blocked due to sigint on outgoing
    // lines (which is not visible here). thus, we only check whether the handshake
    // is correctly initiated and defer the full handshake checking to the testbench.
    `ASSERT(PingHs_A, ##1 $changed(alert_rx_i.ping_p) && state_q == Idle |=>
        $rose(alert_tx_o.alert_p), clk_i, !rst_ni || (alert_tx_o.alert_p == alert_tx_o.alert_n))
  end

  // Test the alert state output.
  `ASSERT(AlertState0_A, alert_set_q === alert_state_o)

  if (IsFatal) begin : gen_fatal_assert
    `ASSERT(AlertState1_A, alert_req_i |=> alert_state_o)
    `ASSERT(AlertState2_A, alert_state_o |=> $stable(alert_state_o))
    `ASSERT(AlertState3_A, alert_ack_o |=> alert_state_o)
  end else begin : gen_recov_assert
    `ASSERT(AlertState1_A, alert_req_i && !alert_clr |=> alert_state_o)
    `ASSERT(AlertState2_A, alert_req_i && alert_ack_o |=> !alert_state_o)
  end

  // The alert test input should not set the alert state register.
  `ASSERT(AlertTest1_A, alert_test_i && !alert_req_i && !alert_state_o |=> $stable(alert_state_o))

  // if alert_req_i is true, handshakes should be continuously repeated
  `ASSERT(AlertHs_A, alert_req_i && state_q == Idle |=> $rose(alert_tx_o.alert_p),
      clk_i, !rst_ni || (alert_tx_o.alert_p == alert_tx_o.alert_n))

  // if alert_test_i is true, handshakes should be continuously repeated
  `ASSERT(AlertTestHs_A, alert_test_i && state_q == Idle |=> $rose(alert_tx_o.alert_p),
      clk_i, !rst_ni || (alert_tx_o.alert_p == alert_tx_o.alert_n))
`endif

`ifdef FPV_ALERT_NO_SIGINT_ERR
  // Assumptions for FPV security countermeasures to ensure the alert protocol functions collectly.
  `ASSUME_FPV(AckPFollowsAlertP_S, alert_rx_i.ack_p == $past(alert_tx_o.alert_p))
  `ASSUME_FPV(AckNFollowsAlertN_S, alert_rx_i.ack_n == $past(alert_tx_o.alert_n))
  `ASSUME_FPV(TriggerAlertInit_S, $stable(rst_ni) == 0 |=> alert_rx_i.ping_p == alert_rx_i.ping_n)
  `ASSUME_FPV(PingDiffPair_S, ##2 alert_rx_i.ping_p != alert_rx_i.ping_n)
`endif
endmodule : prim_alert_sender


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package prim_esc_pkg;

  typedef struct packed {
    logic esc_p;
    logic esc_n;
  } esc_tx_t;

  typedef struct packed {
    logic resp_p;
    logic resp_n;
  } esc_rx_t;

  parameter esc_tx_t ESC_TX_DEFAULT = '{esc_p:  1'b0,
                                        esc_n:  1'b1};

  parameter esc_rx_t ESC_RX_DEFAULT = '{resp_p: 1'b0,
                                        resp_n: 1'b1};

endpackage : prim_esc_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module decodes escalation enable pulses that have been encoded using
// the prim_esc_sender module.
//
// The module supports in-band ping testing of the escalation
// wires. This is accomplished by the sender module that places a single-cycle,
// differentially encoded pulse on esc_p/n which will be interpreted as a ping
// request by the receiver module. The receiver module responds by sending back
// the response pattern "1010".
//
// Native escalation enable pulses are differentiated from ping
// requests by making sure that these pulses are always longer than 1 cycle.
//
// See also: prim_esc_sender, prim_diff_decode, alert_handler

`include "prim_assert.sv"

module prim_esc_receiver
  import prim_esc_pkg::*;
#(
  // The number of escalation severities. Should be set to the Alert Handler's N_ESC_SEV when this
  // primitive is instantiated.
  parameter int N_ESC_SEV = 4,

  // The width of the Alert Handler's ping counter. Should be set to the Alert Handler's PING_CNT_DW
  // when this primitive is instantiated.
  parameter int PING_CNT_DW = 16,

  // This counter monitors incoming ping requests and auto-escalates if the alert handler
  // ceases to send them regularly. The maximum number of cycles between subsequent ping requests
  // is N_ESC_SEV x (2 x 2 x 2**PING_CNT_DW), see also implementation of the ping timer
  // (alert_handler_ping_timer.sv). The timeout counter below uses a timeout that is 4x larger than
  // that in order to incorporate some margin.
  //
  // Do NOT modify this counter value, when instantiating it in the design. It is only exposed to
  // reduce the state space in the FPV testbench.
  localparam int MarginFactor = 4,
  localparam int NumWaitCounts = 2,
  localparam int NumTimeoutCounts = 2,
  parameter int TimeoutCntDw = $clog2(MarginFactor) +
                               $clog2(N_ESC_SEV) +
                               $clog2(NumWaitCounts) +
                               $clog2(NumTimeoutCounts) +
                               PING_CNT_DW
) (
  input           clk_i,
  input           rst_ni,
  // escalation enable
  output logic    esc_req_o,
  // escalation / ping response
  output esc_rx_t esc_rx_o,
  // escalation output diff pair
  input esc_tx_t  esc_tx_i
);

  /////////////////////////////////
  // decode differential signals //
  /////////////////////////////////

  logic esc_level, esc_p, esc_n, sigint_detected;

  // This prevents further tool optimizations of the differential signal.
  prim_buf #(
    .Width(2)
  ) u_prim_buf_esc (
    .in_i({esc_tx_i.esc_n,
           esc_tx_i.esc_p}),
    .out_o({esc_n,
            esc_p})
  );

  prim_diff_decode #(
    .AsyncOn(1'b0)
  ) u_decode_esc (
    .clk_i,
    .rst_ni,
    .diff_pi  ( esc_p           ),
    .diff_ni  ( esc_n           ),
    .level_o  ( esc_level       ),
    .rise_o   (                 ),
    .fall_o   (                 ),
    .event_o  (                 ),
    .sigint_o ( sigint_detected )
  );

  ////////////////////////////////////////////
  // Ping Monitor Counter / Auto Escalation //
  ////////////////////////////////////////////

  // The timeout counter is kicked off when the first ping occurs, and subsequent pings reset
  // the counter to 1. The counter keeps on counting when it is nonzero, and saturates when it
  // has reached its maximum (this state is terminal).
  logic ping_en, timeout_cnt_error;
  logic timeout_cnt_set, timeout_cnt_en;
  logic [TimeoutCntDw-1:0] timeout_cnt;
  assign timeout_cnt_set = (ping_en && !(&timeout_cnt));
  assign timeout_cnt_en = ((timeout_cnt > '0) && !(&timeout_cnt));

  prim_count #(
    .Width(TimeoutCntDw),
    // The escalation receiver behaves differently than other comportable IP. I.e., instead of
    // sending out an alert signal, this condition is handled internally in the alert handler.
    .EnableAlertTriggerSVA(0)
  ) u_prim_count (
    .clk_i,
    .rst_ni,
    .clr_i(1'b0),
    .set_i(timeout_cnt_set),
    .set_cnt_i(TimeoutCntDw'(1)),
    .incr_en_i(timeout_cnt_en),
    .decr_en_i(1'b0),
    .step_i(TimeoutCntDw'(1)),
    .cnt_o(timeout_cnt),
    .cnt_next_o(),
    .err_o(timeout_cnt_error)
  );

  // Escalation is asserted if
  // - requested via the escalation sender/receiver path,
  // - the ping monitor timeout is reached,
  // - the two ping monitor counters are in an inconsistent state.
  logic esc_req;
  prim_sec_anchor_buf #(
    .Width(1)
  ) u_prim_buf_esc_req (
    .in_i(esc_req || (&timeout_cnt) || timeout_cnt_error),
    .out_o(esc_req_o)
  );

  /////////////////
  // RX/TX Logic //
  /////////////////

  typedef enum logic [2:0] {Idle, Check, PingResp, EscResp, SigInt} state_e;
  state_e state_d, state_q;
  logic resp_pd, resp_pq;
  logic resp_nd, resp_nq;

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_flop #(
    .Width(2),
    .ResetValue(2'b10)
  ) u_prim_flop_esc (
    .clk_i,
    .rst_ni,
    .d_i({resp_nd, resp_pd}),
    .q_o({resp_nq, resp_pq})
  );

  assign esc_rx_o.resp_p = resp_pq;
  assign esc_rx_o.resp_n = resp_nq;

  always_comb begin : p_fsm
    // default
    state_d = state_q;
    resp_pd = 1'b0;
    resp_nd = 1'b1;
    esc_req = 1'b0;
    ping_en = 1'b0;

    unique case (state_q)
      // wait for the esc_p/n diff pair
      Idle: begin
        if (esc_level) begin
          state_d = Check;
          resp_pd = ~resp_pq;
          resp_nd = resp_pq;
        end
      end
      // we decide here whether this is only a ping request or
      // whether this is an escalation enable
      Check: begin
        state_d = PingResp;
        resp_pd = ~resp_pq;
        resp_nd = resp_pq;
        if (esc_level) begin
          state_d = EscResp;
          esc_req = 1'b1;
        end
      end
      // finish ping response. in case esc_level is again asserted,
      // we got an escalation signal (pings cannot occur back to back)
      PingResp: begin
        state_d = Idle;
        resp_pd = ~resp_pq;
        resp_nd = resp_pq;
        ping_en = 1'b1;
        if (esc_level) begin
          state_d = EscResp;
          esc_req = 1'b1;
        end
      end
      // we have got an escalation enable pulse,
      // keep on toggling the outputs
      EscResp: begin
        state_d = Idle;
        if (esc_level) begin
          state_d = EscResp;
          resp_pd = ~resp_pq;
          resp_nd = resp_pq;
          esc_req = 1'b1;
        end
      end
      // we have a signal integrity issue at one of
      // the incoming diff pairs. this condition is
      // signalled to the sender by setting the resp
      // diffpair to the same value and continuously
      // toggling them.
      SigInt: begin
        state_d = Idle;
        esc_req = 1'b1;
        if (sigint_detected) begin
          state_d = SigInt;
          resp_pd = ~resp_pq;
          resp_nd = ~resp_pq;
        end
      end
      default: state_d = Idle;
    endcase

    // bail out if a signal integrity issue has been detected
    if (sigint_detected && (state_q != SigInt)) begin
      state_d = SigInt;
      resp_pd = 1'b0;
      resp_nd = 1'b0;
    end
  end


  ///////////////
  // Registers //
  ///////////////

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if (!rst_ni) begin
      state_q <= Idle;
    end else begin
      state_q <= state_d;
    end
  end

  ////////////////
  // assertions //
  ////////////////

  // check whether all outputs have a good known state after reset
  `ASSERT_KNOWN(EscEnKnownO_A, esc_req_o)
  `ASSERT_KNOWN(RespPKnownO_A, esc_rx_o)

  `ASSERT(SigIntCheck0_A, esc_tx_i.esc_p == esc_tx_i.esc_n |=> esc_rx_o.resp_p == esc_rx_o.resp_n)
  `ASSERT(SigIntCheck1_A, esc_tx_i.esc_p == esc_tx_i.esc_n |=> state_q == SigInt)
  // auto-escalate in case of signal integrity issue
  `ASSERT(SigIntCheck2_A, esc_tx_i.esc_p == esc_tx_i.esc_n |=> esc_req_o)
  // correct diff encoding
  `ASSERT(DiffEncCheck_A, esc_tx_i.esc_p ^ esc_tx_i.esc_n |=> esc_rx_o.resp_p ^ esc_rx_o.resp_n)
  // disable in case of signal integrity issue
  `ASSERT(PingRespCheck_A, state_q == Idle ##1 $rose(esc_tx_i.esc_p) ##1 $fell(esc_tx_i.esc_p) |->
      $rose(esc_rx_o.resp_p) ##1 $fell(esc_rx_o.resp_p),
      clk_i, !rst_ni || (esc_tx_i.esc_p == esc_tx_i.esc_n))
  // escalation response needs to continuously toggle
  `ASSERT(EscRespCheck_A, ##1 esc_tx_i.esc_p && $past(esc_tx_i.esc_p) &&
      (esc_tx_i.esc_p ^ esc_tx_i.esc_n) && $past(esc_tx_i.esc_p ^ esc_tx_i.esc_n)
      |=> esc_rx_o.resp_p != $past(esc_rx_o.resp_p))
  // detect escalation pulse
  `ASSERT(EscEnCheck_A,
          esc_tx_i.esc_p && (esc_tx_i.esc_p ^ esc_tx_i.esc_n) && state_q != SigInt
      ##1 esc_tx_i.esc_p && (esc_tx_i.esc_p ^ esc_tx_i.esc_n) |-> esc_req_o)
  // make sure the counter does not wrap around
  `ASSERT(EscCntWrap_A, &timeout_cnt |=> timeout_cnt != 0)
  // if the counter expires, escalation should be asserted
  `ASSERT(EscCntEsc_A, &timeout_cnt |-> esc_req_o)

endmodule : prim_esc_receiver


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module differentially encodes an escalation enable pulse
// of arbitrary width.
//
// The module supports in-band ping testing of the escalation
// wires. This is accomplished by sending out a single, differentially
// encoded pulse on esc_p/n which will be interpreted as a ping
// request by the escalation receiver. Note that ping_req_i shall
// be held high until either ping_ok_o or integ_fail_o is asserted.
//
// Native escalation enable pulses are differentiated from ping
// requests by making sure that these pulses are always longer than 1 cycle.
//
// If there is a differential encoding error, integ_fail_o
// will be asserted.
//
// See also: prim_esc_receiver, prim_diff_decode, alert_handler

`include "prim_assert.sv"

module prim_esc_sender
  import prim_esc_pkg::*;
(
  input           clk_i,
  input           rst_ni,
  // this triggers a ping test. keep asserted until ping_ok_o is pulsed high.
  input           ping_req_i,
  output logic    ping_ok_o,
  // asserted if signal integrity issue detected
  output logic    integ_fail_o,
  // escalation request signal
  input           esc_req_i,
  // escalation / ping response
  input esc_rx_t  esc_rx_i,
  // escalation output diff pair
  output esc_tx_t esc_tx_o
);

  /////////////////////////////////
  // decode differential signals //
  /////////////////////////////////

  logic resp, resp_n, resp_p, sigint_detected;

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_buf #(
    .Width(2)
  ) u_prim_buf_resp (
    .in_i({esc_rx_i.resp_n,
           esc_rx_i.resp_p}),
    .out_o({resp_n,
            resp_p})
  );

  prim_diff_decode #(
    .AsyncOn(1'b0)
  ) u_decode_resp (
    .clk_i,
    .rst_ni,
    .diff_pi  ( resp_p          ),
    .diff_ni  ( resp_n          ),
    .level_o  ( resp            ),
    .rise_o   (                 ),
    .fall_o   (                 ),
    .event_o  (                 ),
    .sigint_o ( sigint_detected )
  );

  //////////////
  // TX Logic //
  //////////////

  logic ping_req_d, ping_req_q;
  logic esc_req_d, esc_req_q, esc_req_q1;

  assign ping_req_d = ping_req_i;
  assign esc_req_d  = esc_req_i;

  // ping enable is 1 cycle pulse
  // escalation pulse is always longer than 2 cycles
  logic esc_p;
  assign esc_p = esc_req_i | esc_req_q | (ping_req_d & ~ping_req_q);

  // This prevents further tool optimizations of the differential signal.
  prim_sec_anchor_buf #(
    .Width(2)
  ) u_prim_buf_esc (
    .in_i({~esc_p,
           esc_p}),
    .out_o({esc_tx_o.esc_n,
            esc_tx_o.esc_p})
  );

  //////////////
  // RX Logic //
  //////////////

  typedef enum logic [2:0] {Idle, CheckEscRespLo, CheckEscRespHi,
    CheckPingResp0, CheckPingResp1, CheckPingResp2, CheckPingResp3} fsm_e;

  fsm_e state_d, state_q;

  always_comb begin : p_fsm
    // default
    state_d      = state_q;
    ping_ok_o    = 1'b0;
    integ_fail_o = sigint_detected;

    unique case (state_q)
      // wait for ping or escalation enable
      Idle: begin
        if (esc_req_i) begin
          state_d = CheckEscRespHi;
        end else if (ping_req_d & ~ping_req_q) begin
          state_d = CheckPingResp0;
        end
        // any assertion of the response signal
        // signal here will trigger a sigint error
        if (resp) begin
          integ_fail_o = 1'b1;
        end
      end
      // check whether response is 0
      CheckEscRespLo: begin
        state_d      = CheckEscRespHi;
        if (!esc_tx_o.esc_p || resp) begin
          state_d = Idle;
          integ_fail_o = sigint_detected | resp;
        end
      end
      // check whether response is 1
      CheckEscRespHi: begin
        state_d = CheckEscRespLo;
        if (!esc_tx_o.esc_p || !resp) begin
          state_d = Idle;
          integ_fail_o = sigint_detected | ~resp;
        end
      end
      // start of ping response sequence
      // we expect the sequence "1010"
      CheckPingResp0: begin
        state_d = CheckPingResp1;
        // abort sequence immediately if escalation is signalled,
        // jump to escalation response checking (lo state)
        if (esc_req_i) begin
          state_d = CheckEscRespLo;
        // abort if response is wrong
        end else if (!resp) begin
          state_d = Idle;
          integ_fail_o = 1'b1;
        end
      end
      CheckPingResp1: begin
        state_d = CheckPingResp2;
        // abort sequence immediately if escalation is signalled,
        // jump to escalation response checking (hi state)
        if (esc_req_i) begin
          state_d = CheckEscRespHi;
        // abort if response is wrong
        end else if (resp) begin
          state_d = Idle;
          integ_fail_o = 1'b1;
        end
      end
      CheckPingResp2: begin
        state_d = CheckPingResp3;
        // abort sequence immediately if escalation is signalled,
        // jump to escalation response checking (lo state)
        if (esc_req_i) begin
          state_d = CheckEscRespLo;
        // abort if response is wrong
        end else if (!resp) begin
          state_d = Idle;
          integ_fail_o = 1'b1;
        end
      end
      CheckPingResp3: begin
        state_d = Idle;
        // abort sequence immediately if escalation is signalled,
        // jump to escalation response checking (hi state)
        if (esc_req_i) begin
          state_d = CheckEscRespHi;
        // abort if response is wrong
        end else if (resp) begin
          integ_fail_o = 1'b1;
        end else begin
          ping_ok_o = ping_req_i;
        end
      end
      default : state_d = Idle;
    endcase

    // a sigint error will reset the state machine
    // and have it pause for two cycles to let the
    // receiver recover
    if (sigint_detected) begin
      ping_ok_o = 1'b0;
      state_d = Idle;
    end

    // escalation takes precedence,
    // immediately return ok in that case
    if ((esc_req_i || esc_req_q || esc_req_q1) && ping_req_i) begin
      ping_ok_o = 1'b1;
    end
  end

  ///////////////
  // Registers //
  ///////////////

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if (!rst_ni) begin
      state_q   <= Idle;
      esc_req_q  <= 1'b0;
      esc_req_q1 <= 1'b0;
      ping_req_q <= 1'b0;
    end else begin
      state_q   <= state_d;
      esc_req_q  <= esc_req_d;
      esc_req_q1 <= esc_req_q;
      ping_req_q <= ping_req_d;
    end
  end

  ////////////////
  // assertions //
  ////////////////

  // check whether all outputs have a good known state after reset
  `ASSERT_KNOWN(PingOkKnownO_A, ping_ok_o)
  `ASSERT_KNOWN(IntegFailKnownO_A, integ_fail_o)
  `ASSERT_KNOWN(EscPKnownO_A, esc_tx_o)

  // diff encoding of output
  `ASSERT(DiffEncCheck_A, esc_tx_o.esc_p ^ esc_tx_o.esc_n)
  // signal integrity check propagation
  `ASSERT(SigIntCheck0_A, esc_rx_i.resp_p == esc_rx_i.resp_n  |-> integ_fail_o)
  // this happens in case we did not get a correct escalation response
  `ASSERT(SigIntCheck1_A, ##1 $rose(esc_req_i) &&
      state_q inside {Idle, CheckPingResp1, CheckPingResp3} ##1 !esc_rx_i.resp_p |->
      integ_fail_o, clk_i, !rst_ni || (esc_rx_i.resp_p == esc_rx_i.resp_n) ||
      (state_q == Idle && resp))
  `ASSERT(SigIntCheck2_A, ##1 $rose(esc_req_i) &&
      state_q inside {CheckPingResp0, CheckPingResp2} ##1 esc_rx_i.resp_p |->
      integ_fail_o, clk_i, !rst_ni || (esc_rx_i.resp_p == esc_rx_i.resp_n) ||
      (state_q == Idle && resp))
  // unexpected response
  `ASSERT(SigIntCheck3_A, state_q == Idle && resp |-> integ_fail_o)
  // signal_int_backward_check
  `ASSERT(SigIntBackCheck_A, integ_fail_o |-> (esc_rx_i.resp_p == esc_rx_i.resp_n) ||
      (esc_rx_i.resp_p && !(state_q == CheckEscRespHi)) ||
      (!esc_rx_i.resp_p && !(state_q == CheckEscRespLo)))
  // state machine CheckEscRespLo and Hi as they are ideal resp signals
  `ASSERT(StateEscRespHiCheck_A, state_q == CheckEscRespLo && esc_tx_o.esc_p && !integ_fail_o |=>
      state_q == CheckEscRespHi)
  `ASSERT(StateEscRespLoCheck_A, state_q == CheckEscRespHi && esc_tx_o.esc_p && !integ_fail_o |=>
      state_q == CheckEscRespLo)
  `ASSERT(StateEscRespHiBackCheck_A, state_q == CheckEscRespHi |-> $past(esc_tx_o.esc_p))
  `ASSERT(StateEscRespLoBackCheck_A, state_q == CheckEscRespLo |-> $past(esc_tx_o.esc_p))
  // check that escalation signal is at least 2 cycles high
  `ASSERT(EscCheck_A, esc_req_i |-> esc_tx_o.esc_p [*2] )
  // escalation / ping collision
  `ASSERT(EscPingCheck_A, esc_req_i && ping_req_i |-> ping_ok_o)
  // check that ping request results in only a single cycle pulse
  `ASSERT(PingCheck_A, ##1 $rose(ping_req_i) |-> esc_tx_o.esc_p ##1 !esc_tx_o.esc_p , clk_i,
      !rst_ni || esc_req_i || integ_fail_o)

endmodule : prim_esc_sender


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Double-synchronizer flop for life cycle control signals with additional
// output buffers and life-cycle specific assertions.
//
// Should be used exactly as recommended in the life cycle controller spec:
// https://docs.opentitan.org/hw/ip/lc_ctrl/doc/index.html#control-signal-propagation

`include "prim_assert.sv"

module prim_lc_sync #(
  // Number of separately buffered output signals.
  // The buffer cells have a don't touch constraint
  // on them such that synthesis tools won't collapse
  // all copies into one signal.
  parameter int NumCopies = 1,
  // This instantiates the synchronizer flops if set to 1.
  // In special cases where the receiver is in the same clock domain as the sender,
  // this can be set to 0. However, it is recommended to leave this at 1.
  parameter bit AsyncOn = 1,
  // 0: reset value is lc_ctrl_pkg::Off
  // 1: reset value is lc_ctrl_pkg::On
  parameter bit ResetValueIsOn = 0
) (
  input                                       clk_i,
  input                                       rst_ni,
  input  lc_ctrl_pkg::lc_tx_t                 lc_en_i,
  output lc_ctrl_pkg::lc_tx_t [NumCopies-1:0] lc_en_o
);

  localparam lc_ctrl_pkg::lc_tx_t LcResetValue = (ResetValueIsOn) ? lc_ctrl_pkg::On :
                                                                  lc_ctrl_pkg::Off;

  `ASSERT_INIT(NumCopiesMustBeGreaterZero_A, NumCopies > 0)

  logic [lc_ctrl_pkg::TxWidth-1:0] lc_en;
  if (AsyncOn) begin : gen_flops
    prim_flop_2sync #(
      .Width(lc_ctrl_pkg::TxWidth),
      .ResetValue(lc_ctrl_pkg::TxWidth'(LcResetValue))
    ) u_prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(lc_en_i),
      .q_o(lc_en)
    );

// Note regarding SVA below:
//
// 1) Without the sampled rst_ni pre-condition, this may cause false assertion failures right after
// a reset release, since the "disable iff" condition with the rst_ni is sampled in the "observed"
// SV scheduler region after all assignments have been evaluated (see also LRM section 16.12, page
// 423). This is a simulation artifact due to reset synchronization in RTL, which releases rst_ni
// on the active clock edge. This causes the assertion to evaluate although the reset was actually
// 0 when entering this simulation cycle.
//
// 2) Similarly to 1) there can be sampling mismatches of the lc_en_i signal since that signal may
// originate from a different clock domain. I.e., in cases where the lc_en_i signal changes exactly
// at the same time that the clk_i signal rises, the SVA will not pick up that change in that clock
// cycle, whereas RTL will because SVAs sample values in the "preponed" region. To that end we make
// use of an RTL helper variable to sample the lc_en_i signal, hence ensuring that there are no
// sampling mismatches.
`ifdef INC_ASSERT
      lc_ctrl_pkg::lc_tx_t lc_en_in_sva_q;
      always_ff @(posedge clk_i) begin
        lc_en_in_sva_q <= lc_en_i;
      end
    `ASSERT(OutputDelay_A,
            rst_ni |-> ##3 lc_en_o == {NumCopies{$past(lc_en_in_sva_q, 2)}} ||
                           ($past(lc_en_in_sva_q, 2) != $past(lc_en_in_sva_q, 1)))
`endif
  end else begin : gen_no_flops
    //VCS coverage off
    // pragma coverage off

    // This unused companion logic helps remove lint errors
    // for modules where clock and reset are used for assertions only
    // or nothing at all.
    // This logic will be removed for sythesis since it is unloaded.
    lc_ctrl_pkg::lc_tx_t unused_logic;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
         unused_logic <= lc_ctrl_pkg::Off;
      end else begin
         unused_logic <= lc_en_i;
      end
    end
    //VCS coverage on
    // pragma coverage on

    assign lc_en = lc_en_i;

    `ASSERT(OutputDelay_A, lc_en_o == {NumCopies{lc_en_i}})
  end

  for (genvar j = 0; j < NumCopies; j++) begin : gen_buffs
    logic [lc_ctrl_pkg::TxWidth-1:0] lc_en_out;
    for (genvar k = 0; k < lc_ctrl_pkg::TxWidth; k++) begin : gen_bits
      prim_sec_anchor_buf u_prim_buf (
        .in_i(lc_en[k]),
        .out_o(lc_en_out[k])
      );
    end
    assign lc_en_o[j] = lc_ctrl_pkg::lc_tx_t'(lc_en_out);
  end

  ////////////////
  // Assertions //
  ////////////////

  // The outputs should be known at all times.
  `ASSERT_KNOWN(OutputsKnown_A, lc_en_o)

endmodule : prim_lc_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This is a draft implementation of a low-latency memory scrambling mechanism.
//
// The module is implemented as a primitive, in the same spirit as similar prim_ram_1p_adv wrappers.
// Hence, it can be conveniently instantiated by comportable IPs (such as OTBN) or in top_earlgrey
// for the main system memory.
//
// The currently implemented architecture uses a reduced-round PRINCE cipher primitive in CTR mode
// in order to (weakly) scramble the data written to the memory macro. Plain CTR mode does not
// diffuse the data since the keystream is just XOR'ed onto it, hence we also we perform byte-wise
// diffusion using a (shallow) substitution/permutation network layers in order to provide a limited
// avalanche effect within a byte.
//
// In order to break the linear addressing space, the address is passed through a bijective
// scrambling function constructed using a (shallow) substitution/permutation and a nonce. Due to
// that nonce, the address mapping is not fully baked into RTL and can be changed at runtime as
// well.
//
// See also: prim_cipher_pkg, prim_prince

`include "prim_assert.sv"

module prim_ram_1p_scr import prim_ram_1p_pkg::*; #(
  parameter  int Depth               = 16*1024, // Needs to be a power of 2 if NumAddrScrRounds > 0.
  parameter  int Width               = 32, // Needs to be byte aligned if byte parity is enabled.
  parameter  int DataBitsPerMask     = 8, // Needs to be set to 8 in case of byte parity.
  parameter  bit EnableParity        = 1, // Enable byte parity.

  // Scrambling parameters. Note that this needs to be low-latency, hence we have to keep the
  // amount of cipher rounds low. PRINCE has 5 half rounds in its original form, which corresponds
  // to 2*5 + 1 effective rounds. Setting this to 2 halves this to approximately 5 effective rounds.
  // Number of PRINCE half rounds, can be [1..5]
  parameter  int NumPrinceRoundsHalf = 2,
  // Number of extra diffusion rounds. Setting this to 0 to disable diffusion.
  parameter  int NumDiffRounds       = 2,
  // This parameter governs the block-width of additional diffusion layers.
  // For intra-byte diffusion, set this parameter to 8.
  parameter  int DiffWidth           = DataBitsPerMask,
  // Number of address scrambling rounds. Setting this to 0 disables address scrambling.
  parameter  int NumAddrScrRounds    = 2,
  // If set to 1, the same 64bit key stream is replicated if the data port is wider than 64bit.
  // If set to 0, the cipher primitive is replicated, and together with a wider nonce input,
  // a unique keystream is generated for the full data width.
  parameter  bit ReplicateKeyStream  = 1'b0,
  // Derived parameters
  localparam int AddrWidth           = prim_util_pkg::vbits(Depth),
  // Depending on the data width, we need to instantiate multiple parallel cipher primitives to
  // create a keystream that is wide enough (PRINCE has a block size of 64bit)
  localparam int NumParScr           = (ReplicateKeyStream) ? 1 : (Width + 63) / 64,
  localparam int NumParKeystr        = (ReplicateKeyStream) ? (Width + 63) / 64 : 1,
  // This is given by the PRINCE cipher primitive. All parallel cipher modules
  // use the same key, but they use a different IV
  localparam int DataKeyWidth        = 128,
  // Each 64 bit scrambling primitive requires a 64bit IV
  localparam int NonceWidth          = 64 * NumParScr
) (
  input                             clk_i,
  input                             rst_ni,

  // Key interface. Memory requests will not be granted if key_valid is set to 0.
  input                             key_valid_i,
  input        [DataKeyWidth-1:0]   key_i,
  input        [NonceWidth-1:0]     nonce_i,

  // Interface to TL-UL SRAM adapter
  input                             req_i,
  output logic                      gnt_o,
  input                             write_i,
  input        [AddrWidth-1:0]      addr_i,
  input        [Width-1:0]          wdata_i,
  input        [Width-1:0]          wmask_i,  // Needs to be byte-aligned for parity
  // On integrity errors, the primitive surpresses any real transaction to the memory.
  input                             intg_error_i,
  output logic [Width-1:0]          rdata_o,
  output logic                      rvalid_o, // Read response (rdata_o) is valid
  output logic [1:0]                rerror_o, // Bit1: Uncorrectable, Bit0: Correctable
  output logic [31:0]               raddr_o,  // Read address for error reporting.

  // config
  input ram_1p_cfg_t                cfg_i
);

  //////////////////////
  // Parameter Checks //
  //////////////////////

  // The depth needs to be a power of 2 in case address scrambling is turned on
  `ASSERT_INIT(DepthPow2Check_A, NumAddrScrRounds <= '0 || 2**$clog2(Depth) == Depth)
  `ASSERT_INIT(DiffWidthMinimum_A, DiffWidth >= 4)
  `ASSERT_INIT(DiffWidthWithParity_A, EnableParity && (DiffWidth == 8) || !EnableParity)

  /////////////////////////////////////////
  // Pending Write and Address Registers //
  /////////////////////////////////////////

  // Writes are delayed by one cycle, such the same keystream generation primitive (prim_prince) can
  // be reused among reads and writes. Note however that with this arrangement, we have to introduce
  // a mechanism to hold a pending write transaction in cases where that transaction is immediately
  // followed by a read. The pending write transaction is written to memory as soon as there is no
  // new read transaction incoming. The latter can be a special case if the incoming read goes to
  // the same address as the pending write. To that end, we detect the address collision and return
  // the data from the write holding register.

  // Read / write strobes
  logic read_en, write_en_d, write_en_q;
  assign gnt_o = req_i & key_valid_i;

  assign read_en = gnt_o & ~write_i;
  assign write_en_d = gnt_o & write_i;

  logic write_pending_q;
  logic addr_collision_d, addr_collision_q;
  logic [AddrWidth-1:0] addr_scr;
  logic [AddrWidth-1:0] waddr_scr_q;
  assign addr_collision_d = read_en & (write_en_q | write_pending_q) & (addr_scr == waddr_scr_q);

  // Macro requests and write strobe
  // The macro operation is silenced if an integrity error is seen
  logic intg_error_buf, intg_error_w_q;
  prim_buf u_intg_error (
    .in_i(intg_error_i),
    .out_o(intg_error_buf)
  );
  logic macro_req;
  assign macro_req   = ~intg_error_w_q & ~intg_error_buf & (read_en | write_en_q | write_pending_q);
  // We are allowed to write a pending write transaction to the memory if there is no incoming read.
  logic macro_write;
  assign macro_write = (write_en_q | write_pending_q) & ~read_en & ~intg_error_w_q;
  // New read write collision
  logic rw_collision;
  assign rw_collision = write_en_q & read_en;

  ////////////////////////
  // Address Scrambling //
  ////////////////////////

  // We only select the pending write address in case there is no incoming read transaction.
  logic [AddrWidth-1:0] addr_mux;
  assign addr_mux = (read_en) ? addr_scr : waddr_scr_q;

  // This creates a bijective address mapping using a substitution / permutation network.
  if (NumAddrScrRounds > 0) begin : gen_addr_scr
    logic [AddrWidth-1:0] addr_scr_nonce;
    assign addr_scr_nonce = nonce_i[NonceWidth - AddrWidth +: AddrWidth];

    prim_subst_perm #(
      .DataWidth ( AddrWidth        ),
      .NumRounds ( NumAddrScrRounds ),
      .Decrypt   ( 0                )
    ) u_prim_subst_perm (
      .data_i ( addr_i         ),
      // Since the counter mode concatenates {nonce_i[NonceWidth-1-AddrWidth:0], addr} to form
      // the IV, the upper AddrWidth bits of the nonce are not used and can be used for address
      // scrambling. In cases where N parallel PRINCE blocks are used due to a data
      // width > 64bit, N*AddrWidth nonce bits are left dangling.
      .key_i  ( addr_scr_nonce ),
      .data_o ( addr_scr       )
    );
  end else begin : gen_no_addr_scr
    assign addr_scr = addr_i;
  end

  // We latch the non-scrambled address for error reporting.
  logic [AddrWidth-1:0] raddr_q;
  assign raddr_o = 32'(raddr_q);

  //////////////////////////////////////////////
  // Keystream Generation for Data Scrambling //
  //////////////////////////////////////////////

  // This encrypts the IV consisting of the nonce and address using the key provided in order to
  // generate the keystream for the data. Note that we instantiate a register halfway within this
  // primitive to balance the delay between request and response side.
  localparam int DataNonceWidth = 64 - AddrWidth;
  logic [NumParScr*64-1:0] keystream;
  logic [NumParScr-1:0][DataNonceWidth-1:0] data_scr_nonce;
  for (genvar k = 0; k < NumParScr; k++) begin : gen_par_scr
    assign data_scr_nonce[k] = nonce_i[k * DataNonceWidth +: DataNonceWidth];

    prim_prince #(
      .DataWidth      (64),
      .KeyWidth       (128),
      .NumRoundsHalf  (NumPrinceRoundsHalf),
      .UseOldKeySched (1'b0),
      .HalfwayDataReg (1'b1), // instantiate a register halfway in the primitive
      .HalfwayKeyReg  (1'b0)  // no need to instantiate a key register as the key remains static
    ) u_prim_prince (
      .clk_i,
      .rst_ni,
      .valid_i ( gnt_o ),
      // The IV is composed of a nonce and the row address
      //.data_i  ( {nonce_i[k * (64 - AddrWidth) +: (64 - AddrWidth)], addr} ),
      .data_i  ( {data_scr_nonce[k], addr_i} ),
      // All parallel scramblers use the same key
      .key_i,
      // Since we operate in counter mode, this can always be set to encryption mode
      .dec_i   ( 1'b0 ),
      // Output keystream to be XOR'ed
      .data_o  ( keystream[k * 64 +: 64] ),
      .valid_o ( )
    );

    // Unread unused bits from keystream
    if (k == NumParKeystr-1 && (Width % 64) > 0) begin : gen_unread_last
      localparam int UnusedWidth = 64 - (Width % 64);
      logic [UnusedWidth-1:0] unused_keystream;
      assign unused_keystream = keystream[(k+1) * 64 - 1 -: UnusedWidth];
    end
  end

  // Replicate keystream if needed
  logic [Width-1:0] keystream_repl;
  assign keystream_repl = Width'({NumParKeystr{keystream}});

  /////////////////////
  // Data Scrambling //
  /////////////////////

  // Data scrambling is a two step process. First, we XOR the write data with the keystream obtained
  // by operating a reduced-round PRINCE cipher in CTR-mode. Then, we diffuse data within each byte
  // in order to get a limited "avalanche" behavior in case parts of the bytes are flipped as a
  // result of a malicious attempt to tamper with the data in memory. We perform the diffusion only
  // within bytes in order to maintain the ability to write individual bytes. Note that the
  // keystream XOR is performed first for the write path such that it can be performed last for the
  // read path. This allows us to hide a part of the combinational delay of the PRINCE primitive
  // behind the propagation delay of the SRAM macro and the per-byte diffusion step.

  logic [Width-1:0] rdata_scr, rdata;
  logic [Width-1:0] wdata_scr_d, wdata_scr_q, wdata_q;
  for (genvar k = 0; k < (Width + DiffWidth - 1) / DiffWidth; k++) begin : gen_diffuse_data
    // If the Width is not divisible by DiffWidth, we need to adjust the width of the last slice.
    localparam int LocalWidth = (Width - k * DiffWidth >= DiffWidth) ? DiffWidth :
                                                                       (Width - k * DiffWidth);

    // Write path. Note that since this does not fan out into the interconnect, the write path is
    // not as critical as the read path below in terms of timing.
    // Apply the keystream first
    logic [LocalWidth-1:0] wdata_xor;
    assign wdata_xor = wdata_q[k*DiffWidth +: LocalWidth] ^
                       keystream_repl[k*DiffWidth +: LocalWidth];

    // Byte aligned diffusion using a substitution / permutation network
    prim_subst_perm #(
      .DataWidth ( LocalWidth       ),
      .NumRounds ( NumDiffRounds ),
      .Decrypt   ( 0                )
    ) u_prim_subst_perm_enc (
      .data_i ( wdata_xor ),
      .key_i  ( '0        ),
      .data_o ( wdata_scr_d[k*DiffWidth +: LocalWidth] )
    );

    // Read path. This is timing critical. The keystream XOR operation is performed last in order to
    // hide the combinational delay of the PRINCE primitive behind the propagation delay of the
    // SRAM and the byte diffusion.
    // Reverse diffusion first
    logic [LocalWidth-1:0] rdata_xor;
    prim_subst_perm #(
      .DataWidth ( LocalWidth       ),
      .NumRounds ( NumDiffRounds ),
      .Decrypt   ( 1                )
    ) u_prim_subst_perm_dec (
      .data_i ( rdata_scr[k*DiffWidth +: LocalWidth] ),
      .key_i  ( '0        ),
      .data_o ( rdata_xor )
    );

    // Apply Keystream, replicate it if needed
    assign rdata[k*DiffWidth +: LocalWidth] = rdata_xor ^
                                              keystream_repl[k*DiffWidth +: LocalWidth];
  end

  ////////////////////////////////////////////////
  // Scrambled data register and forwarding mux //
  ////////////////////////////////////////////////

  // This is the scrambled data holding register for pending writes. This is needed in order to make
  // back to back patterns of the form WR -> RD -> WR work:
  //
  // cycle:          0   |  1   | 2   | 3   |
  // incoming op:    WR0 |  RD  | WR1 | -   |
  // prince:         -   |  WR0 | RD  | WR1 |
  // memory op:      -   |  RD  | WR0 | WR1 |
  //
  // The read transaction in cycle 1 interrupts the first write transaction which has already used
  // the PRINCE primitive for scrambling. If this sequence is followed by another write back-to-back
  // in cycle 2, we cannot use the PRINCE primitive a second time for the first write, and hence
  // need an additional holding register that can buffer the scrambled data of the first write in
  // cycle 1.

  // Clear this if we can write the memory in this cycle. Set only if the current write cannot
  // proceed due to an incoming read operation.
  logic write_scr_pending_d;
  assign write_scr_pending_d = (macro_write)  ? 1'b0 :
                               (rw_collision) ? 1'b1 :
                                                write_pending_q;

  // Select the correct scrambled word to be written, based on whether the word in the scrambled
  // data holding register is valid or not. Note that the write_scr_q register could in theory be
  // combined with the wdata_q register. We don't do that here for timing reasons, since that would
  // require another read data mux to inject the scrambled data into the read descrambling path.
  logic [Width-1:0] wdata_scr;
  assign wdata_scr = (write_pending_q) ? wdata_scr_q : wdata_scr_d;

  logic rvalid_q;
  logic intg_error_r_q;
  logic [Width-1:0] wmask_q;
  always_comb begin : p_forward_mux
    rdata_o = '0;
    rvalid_o = 1'b0;
    // Kill the read response in case an integrity error was seen.
    if (!intg_error_r_q && rvalid_q) begin
      rvalid_o = 1'b1;
      // In case of a collision, we forward the valid bytes of the write data from the unscrambled
      // holding register.
      if (addr_collision_q) begin
        for (int k = 0; k < Width; k++) begin
          if (wmask_q[k]) begin
            rdata_o[k] = wdata_q[k];
          end else begin
            rdata_o[k] = rdata[k];
          end
        end
      // regular reads. note that we just return zero in case
      // an integrity error was signalled.
      end else begin
        rdata_o = rdata;
      end
    end
  end

  ///////////////
  // Registers //
  ///////////////

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_wdata_buf
    if (!rst_ni) begin
      write_pending_q     <= 1'b0;
      addr_collision_q    <= 1'b0;
      rvalid_q            <= 1'b0;
      write_en_q          <= 1'b0;
      intg_error_r_q      <= 1'b0;
      intg_error_w_q      <= 1'b0;
      raddr_q             <= '0;
      waddr_scr_q         <= '0;
      wmask_q             <= '0;
      wdata_q             <= '0;
      wdata_scr_q         <= '0;
    end else begin
      write_pending_q     <= write_scr_pending_d;
      addr_collision_q    <= addr_collision_d;
      rvalid_q            <= read_en;
      write_en_q          <= write_en_d;
      intg_error_r_q      <= intg_error_buf;

      if (read_en) begin
        raddr_q <= addr_i;
      end
      if (write_en_d) begin
        waddr_scr_q    <= addr_scr;
        wmask_q        <= wmask_i;
        wdata_q        <= wdata_i;
        intg_error_w_q <= intg_error_buf;
      end
      if (rw_collision) begin
        wdata_scr_q <= wdata_scr_d;
      end
    end
  end

  //////////////////
  // Memory Macro //
  //////////////////

  prim_ram_1p_adv #(
    .Depth(Depth),
    .Width(Width),
    .DataBitsPerMask(DataBitsPerMask),
    .EnableECC(1'b0),
    .EnableParity(EnableParity),
    .EnableInputPipeline(1'b0),
    .EnableOutputPipeline(1'b0)
  ) u_prim_ram_1p_adv (
    .clk_i,
    .rst_ni,
    .req_i    ( macro_req   ),
    .write_i  ( macro_write ),
    .addr_i   ( addr_mux    ),
    .wdata_i  ( wdata_scr   ),
    .wmask_i  ( wmask_q     ),
    .rdata_o  ( rdata_scr   ),
    .rvalid_o ( ),
    .rerror_o,
    .cfg_i
  );

  `include "prim_util_get_scramble_params.svh"

endmodule : prim_ram_1p_scr


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Data integrity encoder for bus integrity scheme
 */

module tlul_data_integ_enc import tlul_pkg::*; (
  // TL-UL interface
  input        [DataMaxWidth-1:0]               data_i,
  output logic [DataMaxWidth+DataIntgWidth-1:0] data_intg_o
);

  prim_secded_inv_39_32_enc u_data_gen (
    .data_i,
    .data_o(data_intg_o)
  );

endmodule : tlul_data_integ_enc


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Data integrity decoder for bus integrity scheme
 */

module tlul_data_integ_dec import tlul_pkg::*; (
  // TL-UL interface
  input        [DataMaxWidth+DataIntgWidth-1:0] data_intg_i,
  output logic                                  data_err_o
);

  logic [1:0] data_err;
  prim_secded_inv_39_32_dec u_data_chk (
    .data_i(data_intg_i),
    .data_o(),
    .syndrome_o(),
    .err_o(data_err)
  );

  assign data_err_o = |data_err;

endmodule : tlul_data_integ_dec


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL command integrity generator
 */

module tlul_cmd_intg_gen import tlul_pkg::*; #(
  parameter bit EnableDataIntgGen = 1'b1
) (
  // TL-UL interface
  input  tl_h2d_t tl_i,
  output tl_h2d_t tl_o
);

  tl_h2d_cmd_intg_t cmd;
  assign cmd = extract_h2d_cmd_intg(tl_i);
  logic [H2DCmdMaxWidth-1:0] unused_cmd_payload;

  logic [H2DCmdIntgWidth-1:0] cmd_intg;
  prim_secded_inv_64_57_enc u_cmd_gen (
    .data_i(H2DCmdMaxWidth'(cmd)),
    .data_o({cmd_intg, unused_cmd_payload})
  );

  logic [top_pkg::TL_DW-1:0] data_final;
  logic [DataIntgWidth-1:0] data_intg;

  if (EnableDataIntgGen) begin : gen_data_intg
    assign data_final = tl_i.a_data;

    logic [DataMaxWidth-1:0] unused_data;
    prim_secded_inv_39_32_enc u_data_gen (
      .data_i(DataMaxWidth'(data_final)),
      .data_o({data_intg, unused_data})
    );
  end else begin : gen_passthrough_data_intg
    assign data_final = tl_i.a_data;
    assign data_intg = tl_i.a_user.data_intg;
  end

  always_comb begin
    tl_o = tl_i;
    tl_o.a_data = data_final;
    tl_o.a_user.cmd_intg = cmd_intg;
    tl_o.a_user.data_intg = data_intg;
  end


  logic unused_tl;
  assign unused_tl = ^tl_i;

  `ASSERT_INIT(PayMaxWidthCheck_A, $bits(tl_h2d_cmd_intg_t) <= H2DCmdMaxWidth)

endmodule : tlul_cmd_intg_gen


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL command integrity check
 */

module tlul_cmd_intg_chk import tlul_pkg::*; (
  // TL-UL interface
  input  tl_h2d_t tl_i,

  // error output
  output logic err_o
);

  logic [1:0] err;
  logic data_err;
  tl_h2d_cmd_intg_t cmd;
  assign cmd = extract_h2d_cmd_intg(tl_i);

  prim_secded_inv_64_57_dec u_chk (
    .data_i({tl_i.a_user.cmd_intg, H2DCmdMaxWidth'(cmd)}),
    .data_o(),
    .syndrome_o(),
    .err_o(err)
  );

  tlul_data_integ_dec u_tlul_data_integ_dec (
    .data_intg_i({tl_i.a_user.data_intg, DataMaxWidth'(tl_i.a_data)}),
    .data_err_o(data_err)
  );

  // error output is transactional, it is up to the instantiating module
  // to determine if a permanent latch is feasible
  // [LOWRISC] err and data_err is unknown when a_valid is low, so we can't cover
  // the condition coverage - (|err | (|data_err)) == 0/1, when a_valid = 0, which is
  // fine as driving unknown is better. `err_o` is used as a condition in other places,
  // which needs to be covered with 0 and 1, so it's OK to disable the entire coverage.
  //VCS coverage off
  // pragma coverage off
  // assign err_o = tl_i.a_valid & (|err | (|data_err));
  //zdr
  assign err_o = 1'b0;
  //VCS coverage on
  // pragma coverage on

  logic unused_tl;
  assign unused_tl = |tl_i;

  `ASSERT_INIT(PayLoadWidthCheck, $bits(tl_h2d_cmd_intg_t) <= H2DCmdMaxWidth)

endmodule // tlul_payload_chk


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL response integrity generator
 */

module tlul_rsp_intg_gen import tlul_pkg::*; #(
  parameter bit EnableRspIntgGen = 1'b1,
  parameter bit EnableDataIntgGen = 1'b1
) (
  // TL-UL interface
  input  tl_d2h_t tl_i,
  output tl_d2h_t tl_o
);

  logic [D2HRspIntgWidth-1:0] rsp_intg;
  if (EnableRspIntgGen) begin : gen_rsp_intg
    tl_d2h_rsp_intg_t rsp;
    logic [D2HRspMaxWidth-1:0] unused_payload;

    assign rsp = extract_d2h_rsp_intg(tl_i);

    prim_secded_inv_64_57_enc u_rsp_gen (
      .data_i(D2HRspMaxWidth'(rsp)),
      .data_o({rsp_intg, unused_payload})
    );
  end else begin : gen_passthrough_rsp_intg
    assign rsp_intg = tl_i.d_user.rsp_intg;
  end

  logic [DataIntgWidth-1:0] data_intg;
  if (EnableDataIntgGen) begin : gen_data_intg
    logic [DataMaxWidth-1:0] unused_data;
    tlul_data_integ_enc u_tlul_data_integ_enc (
      .data_i(DataMaxWidth'(tl_i.d_data)),
      .data_intg_o({data_intg, unused_data})
    );
  end else begin : gen_passthrough_data_intg
    assign data_intg = tl_i.d_user.data_intg;
  end

  always_comb begin
    tl_o = tl_i;
    tl_o.d_user.rsp_intg = rsp_intg;
    tl_o.d_user.data_intg = data_intg;
  end

  logic unused_tl;
  assign unused_tl = ^tl_i;


  `ASSERT_INIT(PayLoadWidthCheck, $bits(tl_d2h_rsp_intg_t) <= D2HRspMaxWidth)
  `ASSERT_INIT(DataWidthCheck_A, $bits(tl_i.d_data) <= DataMaxWidth)

endmodule // tlul_rsp_intg_gen


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL response integrity check
 */

module tlul_rsp_intg_chk import tlul_pkg::*; #(
  parameter bit EnableRspDataIntgCheck = 0
) (
  // TL-UL interface
  input  tl_d2h_t tl_i,

  // error output
  output logic err_o
);

  logic [1:0] rsp_err;
  tl_d2h_rsp_intg_t rsp;
  assign rsp = extract_d2h_rsp_intg(tl_i);

  prim_secded_inv_64_57_dec u_chk (
    .data_i({tl_i.d_user.rsp_intg, D2HRspMaxWidth'(rsp)}),
    .data_o(),
    .syndrome_o(),
    .err_o(rsp_err)
  );

  logic rsp_data_err;
  if (EnableRspDataIntgCheck) begin : gen_rsp_data_intg_check
    tlul_data_integ_dec u_tlul_data_integ_dec (
      .data_intg_i({tl_i.d_user.data_intg, DataMaxWidth'(tl_i.d_data)}),
      .data_err_o(rsp_data_err)
    );
  end else begin : gen_no_rsp_data_intg_check
    assign rsp_data_err = 1'b0;
  end

  // error is not permanently latched as rsp_intg_chk is typically
  // used near the host.
  // if the error is permanent, it would imply the host could forever
  // receive bus errors and lose all ability to debug.
  // It should be up to the host to determine the permanence of this error.
  assign err_o = tl_i.d_valid & (|rsp_err | rsp_data_err);

  logic unused_tl;
  assign unused_tl = |tl_i;

  `ASSERT_INIT(PayLoadWidthCheck, $bits(tl_d2h_rsp_intg_t) <= D2HRspMaxWidth)

endmodule // tlul_rsp_intg_chk


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package edn_reg_pkg;

  // Param list
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 7;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } edn_cmd_req_done;
    struct packed {
      logic        q;
    } edn_fatal_err;
  } edn_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } edn_cmd_req_done;
    struct packed {
      logic        q;
    } edn_fatal_err;
  } edn_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } edn_cmd_req_done;
    struct packed {
      logic        q;
      logic        qe;
    } edn_fatal_err;
  } edn_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_alert;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_alert;
  } edn_reg2hw_alert_test_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } edn_enable;
    struct packed {
      logic [3:0]  q;
    } boot_req_mode;
    struct packed {
      logic [3:0]  q;
    } auto_req_mode;
    struct packed {
      logic [3:0]  q;
    } cmd_fifo_rst;
  } edn_reg2hw_ctrl_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } edn_reg2hw_boot_ins_cmd_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } edn_reg2hw_boot_gen_cmd_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } edn_reg2hw_sw_cmd_req_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } edn_reg2hw_reseed_cmd_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } edn_reg2hw_generate_cmd_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } edn_reg2hw_max_num_reqs_between_reseeds_reg_t;

  typedef struct packed {
    logic [4:0]  q;
    logic        qe;
  } edn_reg2hw_err_code_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } edn_cmd_req_done;
    struct packed {
      logic        d;
      logic        de;
    } edn_fatal_err;
  } edn_hw2reg_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } cmd_rdy;
    struct packed {
      logic        d;
      logic        de;
    } cmd_sts;
  } edn_hw2reg_sw_cmd_sts_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } edn_enable_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } boot_req_mode_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } auto_req_mode_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } cmd_fifo_rst_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } edn_bus_cmp_alert;
  } edn_hw2reg_recov_alert_sts_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } sfifo_rescmd_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_gencmd_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_output_err;
    struct packed {
      logic        d;
      logic        de;
    } edn_ack_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } edn_main_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } edn_cntr_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_write_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_read_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_state_err;
  } edn_hw2reg_err_code_reg_t;

  typedef struct packed {
    logic [8:0]  d;
    logic        de;
  } edn_hw2reg_main_sm_state_reg_t;

  // Register -> HW type
  typedef struct packed {
    edn_reg2hw_intr_state_reg_t intr_state; // [229:228]
    edn_reg2hw_intr_enable_reg_t intr_enable; // [227:226]
    edn_reg2hw_intr_test_reg_t intr_test; // [225:222]
    edn_reg2hw_alert_test_reg_t alert_test; // [221:218]
    edn_reg2hw_ctrl_reg_t ctrl; // [217:202]
    edn_reg2hw_boot_ins_cmd_reg_t boot_ins_cmd; // [201:170]
    edn_reg2hw_boot_gen_cmd_reg_t boot_gen_cmd; // [169:138]
    edn_reg2hw_sw_cmd_req_reg_t sw_cmd_req; // [137:105]
    edn_reg2hw_reseed_cmd_reg_t reseed_cmd; // [104:72]
    edn_reg2hw_generate_cmd_reg_t generate_cmd; // [71:39]
    edn_reg2hw_max_num_reqs_between_reseeds_reg_t max_num_reqs_between_reseeds; // [38:6]
    edn_reg2hw_err_code_test_reg_t err_code_test; // [5:0]
  } edn_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    edn_hw2reg_intr_state_reg_t intr_state; // [45:42]
    edn_hw2reg_sw_cmd_sts_reg_t sw_cmd_sts; // [41:38]
    edn_hw2reg_recov_alert_sts_reg_t recov_alert_sts; // [37:28]
    edn_hw2reg_err_code_reg_t err_code; // [27:10]
    edn_hw2reg_main_sm_state_reg_t main_sm_state; // [9:0]
  } edn_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] EDN_INTR_STATE_OFFSET = 7'h 0;
  parameter logic [BlockAw-1:0] EDN_INTR_ENABLE_OFFSET = 7'h 4;
  parameter logic [BlockAw-1:0] EDN_INTR_TEST_OFFSET = 7'h 8;
  parameter logic [BlockAw-1:0] EDN_ALERT_TEST_OFFSET = 7'h c;
  parameter logic [BlockAw-1:0] EDN_REGWEN_OFFSET = 7'h 10;
  parameter logic [BlockAw-1:0] EDN_CTRL_OFFSET = 7'h 14;
  parameter logic [BlockAw-1:0] EDN_BOOT_INS_CMD_OFFSET = 7'h 18;
  parameter logic [BlockAw-1:0] EDN_BOOT_GEN_CMD_OFFSET = 7'h 1c;
  parameter logic [BlockAw-1:0] EDN_SW_CMD_REQ_OFFSET = 7'h 20;
  parameter logic [BlockAw-1:0] EDN_SW_CMD_STS_OFFSET = 7'h 24;
  parameter logic [BlockAw-1:0] EDN_RESEED_CMD_OFFSET = 7'h 28;
  parameter logic [BlockAw-1:0] EDN_GENERATE_CMD_OFFSET = 7'h 2c;
  parameter logic [BlockAw-1:0] EDN_MAX_NUM_REQS_BETWEEN_RESEEDS_OFFSET = 7'h 30;
  parameter logic [BlockAw-1:0] EDN_RECOV_ALERT_STS_OFFSET = 7'h 34;
  parameter logic [BlockAw-1:0] EDN_ERR_CODE_OFFSET = 7'h 38;
  parameter logic [BlockAw-1:0] EDN_ERR_CODE_TEST_OFFSET = 7'h 3c;
  parameter logic [BlockAw-1:0] EDN_MAIN_SM_STATE_OFFSET = 7'h 40;

  // Reset values for hwext registers and their fields
  parameter logic [1:0] EDN_INTR_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] EDN_INTR_TEST_EDN_CMD_REQ_DONE_RESVAL = 1'h 0;
  parameter logic [0:0] EDN_INTR_TEST_EDN_FATAL_ERR_RESVAL = 1'h 0;
  parameter logic [1:0] EDN_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] EDN_ALERT_TEST_RECOV_ALERT_RESVAL = 1'h 0;
  parameter logic [0:0] EDN_ALERT_TEST_FATAL_ALERT_RESVAL = 1'h 0;
  parameter logic [31:0] EDN_SW_CMD_REQ_RESVAL = 32'h 0;
  parameter logic [31:0] EDN_RESEED_CMD_RESVAL = 32'h 0;
  parameter logic [31:0] EDN_GENERATE_CMD_RESVAL = 32'h 0;

  // Register index
  typedef enum int {
    EDN_INTR_STATE,
    EDN_INTR_ENABLE,
    EDN_INTR_TEST,
    EDN_ALERT_TEST,
    EDN_REGWEN,
    EDN_CTRL,
    EDN_BOOT_INS_CMD,
    EDN_BOOT_GEN_CMD,
    EDN_SW_CMD_REQ,
    EDN_SW_CMD_STS,
    EDN_RESEED_CMD,
    EDN_GENERATE_CMD,
    EDN_MAX_NUM_REQS_BETWEEN_RESEEDS,
    EDN_RECOV_ALERT_STS,
    EDN_ERR_CODE,
    EDN_ERR_CODE_TEST,
    EDN_MAIN_SM_STATE
  } edn_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] EDN_PERMIT [17] = '{
    4'b 0001, // index[ 0] EDN_INTR_STATE
    4'b 0001, // index[ 1] EDN_INTR_ENABLE
    4'b 0001, // index[ 2] EDN_INTR_TEST
    4'b 0001, // index[ 3] EDN_ALERT_TEST
    4'b 0001, // index[ 4] EDN_REGWEN
    4'b 0011, // index[ 5] EDN_CTRL
    4'b 1111, // index[ 6] EDN_BOOT_INS_CMD
    4'b 1111, // index[ 7] EDN_BOOT_GEN_CMD
    4'b 1111, // index[ 8] EDN_SW_CMD_REQ
    4'b 0001, // index[ 9] EDN_SW_CMD_STS
    4'b 1111, // index[10] EDN_RESEED_CMD
    4'b 1111, // index[11] EDN_GENERATE_CMD
    4'b 1111, // index[12] EDN_MAX_NUM_REQS_BETWEEN_RESEEDS
    4'b 0011, // index[13] EDN_RECOV_ALERT_STS
    4'b 1111, // index[14] EDN_ERR_CODE
    4'b 0001, // index[15] EDN_ERR_CODE_TEST
    4'b 0011  // index[16] EDN_MAIN_SM_STATE
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//


package edn_pkg;
  ///////////////////////////
  // Peripheral Interfaces //
  ///////////////////////////

  parameter int unsigned   ENDPOINT_BUS_WIDTH = 32;
  parameter int unsigned   FIPS_ENDPOINT_BUS_WIDTH = entropy_src_pkg::FIPS_BUS_WIDTH +
                           ENDPOINT_BUS_WIDTH;

  // EDN request interface
  typedef struct packed {
    logic                                 edn_req;
  } edn_req_t;
  typedef struct packed {
    logic                                 edn_ack;
    logic                                 edn_fips;
    logic [ENDPOINT_BUS_WIDTH-1:0]        edn_bus;
  } edn_rsp_t;

  parameter edn_req_t EDN_REQ_DEFAULT = '0;
  parameter edn_rsp_t EDN_RSP_DEFAULT = '0;

  typedef enum logic [8:0] {
    Idle              = 9'b110000101, // idle
    BootLoadIns       = 9'b110110111, // boot: load the instantiate command
    BootLoadGen       = 9'b000000011, // boot: load the generate command
    BootInsAckWait    = 9'b011010010, // boot: wait for instantiate command ack
    BootCaptGenCnt    = 9'b010111010, // boot: capture the gen fifo count
    BootSendGenCmd    = 9'b011100100, // boot: send the generate command
    BootGenAckWait    = 9'b101101100, // boot: wait for generate command ack
    BootPulse         = 9'b100001010, // boot: signal a done pulse
    BootDone          = 9'b011011111, // boot: stay in done state until reset
    AutoLoadIns       = 9'b001110000, // auto: load the instantiate command
    AutoFirstAckWait  = 9'b001001101, // auto: wait for first instantiate command ack
    AutoAckWait       = 9'b101100011, // auto: wait for instantiate command ack
    AutoDispatch      = 9'b110101110, // auto: determine next command to be sent
    AutoCaptGenCnt    = 9'b000110101, // auto: capture the gen fifo count
    AutoSendGenCmd    = 9'b111111000, // auto: send the generate command
    AutoCaptReseedCnt = 9'b000100110, // auto: capture the reseed fifo count
    AutoSendReseedCmd = 9'b101010110, // auto: send the reseed command
    SWPortMode        = 9'b100111001, // swport: no hw request mode
    Error             = 9'b010010001  // illegal state reached and hang
  } state_e;

endpackage : edn_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

package otbn_pkg;

  // Global Constants ==============================================================================

  // Data path width for BN (wide) instructions, in bits.
  parameter int WLEN = 256;

  // "Extended" WLEN: the size of the datapath with added integrity bits
  parameter int ExtWLEN = WLEN * 39 / 32;

  // Width of base (32b) data path with added integrity bits
  parameter int BaseIntgWidth = 39;

  // Number of 32-bit words per WLEN
  parameter int BaseWordsPerWLEN = WLEN / 32;

  // Number of flag groups
  parameter int NFlagGroups = 2;

  // Width of the GPR index/address
  parameter int GprAw = 5;

  // Number of General Purpose Registers (GPRs)
  parameter int NGpr = 2 ** GprAw;

  // Width of the WDR index/address
  parameter int WdrAw = 5;

  // Number of Wide Data Registers (WDRs)
  parameter int NWdr = 2 ** WdrAw;

  // Width of entropy input
  parameter int EdnDataWidth = 256;

  parameter int SideloadKeyWidth = 384;

  parameter int unsigned LoopStackDepth = 8;

  // Zero word in the implemented ECC scheme. If changing the ECC scheme, this has to be changed,
  // and vice-versa.
  localparam logic [BaseIntgWidth-1:0] EccZeroWord     = prim_secded_pkg::SecdedInv3932ZeroWord;
  localparam logic [ExtWLEN-1:0]       EccWideZeroWord = {BaseWordsPerWLEN{EccZeroWord}};

  // Size of DMEM scratch area. The total DMEM size is OTBN_DMEM_SIZE + DmemScratchSizeByte. Note
  // that some of the Python tooling depends on this parameter (it needs to know the full DMEM size,
  // but regtool only gives it OTBN_DMEM_SIZE). If changing this, you'll also need to edit
  // _DmemScratchSizeBytes in util/shared/mem_layout.py
  parameter int DmemScratchSizeByte = 1024;

  // Toplevel constants ============================================================================

  parameter int AlertFatal = 0;
  parameter int AlertRecov = 1;

  // Register file implementation selection enum.
  typedef enum integer {
    RegFileFF    = 0, // Generic flip-flop based implementation
    RegFileFPGA  = 1  // FPGA implmentation, does infer RAM primitives.
  } regfile_e;

  // Command to execute. See the CMD register description in otbn.hjson for details.
  typedef enum logic [7:0] {
    CmdExecute     = 8'hd8,
    CmdSecWipeDmem = 8'hc3,
    CmdSecWipeImem = 8'h1e
  } cmd_e;

  // Status register values. See the STATUS register description in otbn.hjson for details.
  typedef enum logic [7:0] {
    StatusIdle            = 8'h00,
    StatusBusyExecute     = 8'h01,
    StatusBusySecWipeDmem = 8'h02,
    StatusBusySecWipeImem = 8'h03,
    StatusBusySecWipeInt  = 8'h04,
    StatusLocked          = 8'hFF
  } status_e;

  function automatic logic is_busy_status(status_e status);
    return status inside {StatusBusyExecute,
                          StatusBusySecWipeDmem,
                          StatusBusySecWipeImem,
                          StatusBusySecWipeInt};
  endfunction

  // Error bits
  //
  // Note: These errors are duplicated in other places. If updating them here, update those too.
  typedef struct packed {
    logic fatal_software;
    logic lifecycle_escalation;
    logic illegal_bus_access;
    logic bad_internal_state;
    logic bus_intg_violation;
    logic reg_intg_violation;
    logic dmem_intg_violation;
    logic imem_intg_violation;
    logic rnd_fips_chk_fail;
    logic rnd_rep_chk_fail;
    logic key_invalid;
    logic loop;
    logic illegal_insn;
    logic call_stack;
    logic bad_insn_addr;
    logic bad_data_addr;
  } err_bits_t;

  // Wrappers for classifying bad internal states
  typedef struct packed {
    logic alu_bignum_err;
    logic mac_bignum_err;
    logic ispr_bignum_err;
    logic controller_err;
    logic rf_err;
    logic rd_err;
  } predec_err_t;

  typedef struct packed {
    logic spr_urnd_acks;
    logic spr_rnd_acks;
    logic spr_secwipe_reqs;
    logic mubi_rma_err;
    logic mubi_urnd_err;
    logic state_err;
  } start_stop_bad_int_t;

  typedef struct packed {
    logic loop_hw_cnt_err;
    logic loop_hw_stack_cnt_err;
    logic loop_hw_intg_err;
    logic rf_base_call_stack_err;
    logic spr_secwipe_acks;
    logic state_err;
    logic controller_mubi_err;
  } controller_bad_int_t;

  typedef struct packed {
    logic imem_gnt_missed_err;
    logic dmem_gnt_missed_err;
  } missed_gnt_t;

  typedef struct packed {
    logic rf_base_intg_err;
    logic rf_bignum_intg_err;
    logic mod_ispr_intg_err;
    logic acc_ispr_intg_err;
    logic loop_stack_addr_intg_err;
    logic insn_fetch_intg_err;
  } internal_intg_err_t;

  // All the error signals that can be generated directly from the controller. Note that this is
  // organised to include every software error (including 'call_stack', which actually gets fed in
  // from the base register file)
  typedef struct packed {
    logic fatal_software;
    logic bad_internal_state;
    logic reg_intg_violation;
    logic key_invalid;
    logic loop;
    logic illegal_insn;
    logic call_stack;
    logic bad_insn_addr;
    logic bad_data_addr;
  } controller_err_bits_t;

  // All the error signals that can be generated somewhere inside otbn_core
  typedef struct packed {
    logic fatal_software;
    logic bad_internal_state;
    logic reg_intg_violation;
    logic dmem_intg_violation;
    logic imem_intg_violation;
    logic rnd_fips_chk_fail;
    logic rnd_rep_chk_fail;
    logic key_invalid;
    logic loop;
    logic illegal_insn;
    logic call_stack;
    logic bad_insn_addr;
    logic bad_data_addr;
  } core_err_bits_t;

  // The error signals that are generated outside of otbn_core
  typedef struct packed {
    logic lifecycle_escalation;
    logic illegal_bus_access;
    logic bad_internal_state;
    logic bus_intg_violation;
  } non_core_err_bits_t;

  // Constants =====================================================================================

  typedef enum logic {
    InsnSubsetBase = 1'b0,  // Base (RV32/Narrow) Instruction Subset
    InsnSubsetBignum = 1'b1 // Big Number (BN/Wide) Instruction Subset
  } insn_subset_e;

  // Opcodes (field [6:0] in the instruction), matching the RISC-V specification for the base
  // instruction subset.
  typedef enum logic [6:0] {
    InsnOpcodeBaseLoad       = 7'h03,
    InsnOpcodeBaseMemMisc    = 7'h0f,
    InsnOpcodeBaseOpImm      = 7'h13,
    InsnOpcodeBaseStore      = 7'h23,
    InsnOpcodeBaseOp         = 7'h33,
    InsnOpcodeBaseLui        = 7'h37,
    InsnOpcodeBaseBranch     = 7'h63,
    InsnOpcodeBaseJalr       = 7'h67,
    InsnOpcodeBaseJal        = 7'h6f,
    InsnOpcodeBaseSystem     = 7'h73,
    InsnOpcodeBignumMisc     = 7'h0B,
    InsnOpcodeBignumArith    = 7'h2B,
    InsnOpcodeBignumMulqacc  = 7'h3B,
    InsnOpcodeBignumBaseMisc = 7'h7B
  } insn_opcode_e;

  typedef enum logic [3:0] {
    AluOpBaseAdd,
    AluOpBaseSub,

    AluOpBaseXor,
    AluOpBaseOr,
    AluOpBaseAnd,
    AluOpBaseNot,

    AluOpBaseSra,
    AluOpBaseSrl,
    AluOpBaseSll
  } alu_op_base_e;

  typedef enum logic [3:0] {
    AluOpBignumAdd,
    AluOpBignumAddc,
    AluOpBignumAddm,

    AluOpBignumSub,
    AluOpBignumSubb,
    AluOpBignumSubm,

    AluOpBignumRshi,

    AluOpBignumXor,
    AluOpBignumOr,
    AluOpBignumAnd,
    AluOpBignumNot,

    AluOpBignumNone
  } alu_op_bignum_e;

  typedef enum logic [1:0] {
    AluOpLogicXor = 2'h0,
    AluOpLogicOr  = 2'h1,
    AluOpLogicAnd = 2'h2,
    AluOpLogicNot = 2'h3
  } alu_op_logic_e;

  typedef enum logic {
    ComparisonOpBaseEq,
    ComparisonOpBaseNeq
  } comparison_op_base_e;

  // Operand a source selection
  typedef enum logic [1:0] {
    OpASelRegister  = 'd0,
    OpASelZero = 'd1,
    OpASelCurrPc = 'd2
  } op_a_sel_e;

  // Operand b source selection
  typedef enum logic {
    OpBSelRegister  = 'd0,
    OpBSelImmediate = 'd1
  } op_b_sel_e;

  // Immediate b selection for base ISA
  typedef enum logic [2:0] {
    ImmBaseBI,
    ImmBaseBS,
    ImmBaseBB,
    ImmBaseBU,
    ImmBaseBJ,
    ImmBaseBL,
    ImmBaseBX
  } imm_b_sel_base_e;

  // Shift amount select for bignum ISA
  typedef enum logic [1:0] {
    ShamtSelBignumA,
    ShamtSelBignumS,
    ShamtSelBignumZero
  } shamt_sel_bignum_e;

  // Regfile write data selection
  typedef enum logic [2:0] {
    RfWdSelEx,
    RfWdSelNextPc,
    RfWdSelLsu,
    RfWdSelIspr,
    RfWdSelIncr,
    RfWdSelMac,
    RfWdSelMovSel
  } rf_wd_sel_e;

  // Control and Status Registers (CSRs)
  parameter int CsrNumWidth = 12;
  typedef enum logic [CsrNumWidth-1:0] {
    // Address ranges follow the RISC-V Privileged Specification v1.11
    // 0x7C0-0x7FF Custom read/write
    CsrFg0         = 12'h7C0,
    CsrFg1         = 12'h7C1,
    CsrFlags       = 12'h7C8,
    CsrMod0        = 12'h7D0,
    CsrMod1        = 12'h7D1,
    CsrMod2        = 12'h7D2,
    CsrMod3        = 12'h7D3,
    CsrMod4        = 12'h7D4,
    CsrMod5        = 12'h7D5,
    CsrMod6        = 12'h7D6,
    CsrMod7        = 12'h7D7,
    CsrRndPrefetch = 12'h7D8,

    // 0xFC0-0xFFF Custom read-only
    CsrRnd         = 12'hFC0,
    CsrUrnd        = 12'hFC1
  } csr_e;

  // Wide Special Purpose Registers (WSRs)
  parameter int NWsr = 8; // Number of WSRs
  parameter int WsrNumWidth = $clog2(NWsr);
  typedef enum logic [WsrNumWidth-1:0] {
    WsrMod    = 'd0,
    WsrRnd    = 'd1,
    WsrUrnd   = 'd2,
    WsrAcc    = 'd3,
    WsrKeyS0L = 'd4,
    WsrKeyS0H = 'd5,
    WsrKeyS1L = 'd6,
    WsrKeyS1H = 'd7
  } wsr_e;

  // Internal Special Purpose Registers (ISPRs)
  // CSRs and WSRs have some overlap into what they map into. ISPRs are the actual registers in the
  // design which CSRs and WSRs are mapped on to.
  parameter int NIspr = 9;
  parameter int IsprNumWidth = $clog2(NIspr);
  typedef enum logic [IsprNumWidth-1:0] {
    IsprMod    = 'd0,
    IsprRnd    = 'd1,
    IsprAcc    = 'd2,
    IsprFlags  = 'd3,
    IsprUrnd   = 'd4,
    IsprKeyS0L = 'd5,
    IsprKeyS0H = 'd6,
    IsprKeyS1L = 'd7,
    IsprKeyS1H = 'd8
  } ispr_e;

  typedef logic [$clog2(NFlagGroups)-1:0] flag_group_t;

  typedef struct packed {
    logic Z;
    logic L;
    logic M;
    logic C;
  } flags_t;

  localparam int FlagsWidth = $bits(flags_t);

  typedef enum logic [$clog2(FlagsWidth)-1:0] {
    FlagC = 'd0,
    FlagM = 'd1,
    FlagL = 'd2,
    FlagZ = 'd3
  } flag_e;

  // Structures for decoded instructions, grouped into three:
  // - insn_dec_shared_t - Anything that applies to both bignum and base microarchitecture
  // - insn_dec_base_t - Anything that only applies to the base side microarchitecture
  // - insn_dec_bignum_t - Anything that only applies to bignum side microarchitecture

  typedef struct packed {
    insn_subset_e           subset;
    logic                   ecall_insn;
    logic                   ld_insn;
    logic                   st_insn;
    logic                   branch_insn;
    logic                   jump_insn;
    logic                   loop_insn;
    logic                   ispr_rd_insn;
    logic                   ispr_wr_insn;
    logic                   ispr_rs_insn;
    logic [NFlagGroups-1:0] ispr_flags_wr;
  } insn_dec_shared_t;

  typedef struct packed {
    logic [4:0]          d;             // Destination register
    logic [4:0]          a;             // First source register
    logic [4:0]          b;             // Second source register
    logic [31:0]         i;             // Immediate
    alu_op_base_e        alu_op;
    comparison_op_base_e comparison_op;
    op_a_sel_e           op_a_sel;
    op_b_sel_e           op_b_sel;
    logic                rf_ren_a;
    logic                rf_ren_b;
    logic                rf_we;
    rf_wd_sel_e          rf_wdata_sel;
    logic [11:0]         loop_bodysize;
    logic                loop_immediate;
  } insn_dec_base_t;

  typedef struct packed {
    logic [WdrAw-1:0]        d;           // Destination register
    logic [WdrAw-1:0]        a;           // First source register
    logic [WdrAw-1:0]        b;           // Second source register
    logic [WLEN-1:0]         i;           // Immediate

    logic                    rf_a_indirect; // Indirect lookup, bignum register index a comes from
                                            // base register a read
    logic                    rf_b_indirect; // Indirect lookup, bignum register index b comes from
                                            // base register b read
    logic                    rf_d_indirect; // Indirect lookup, bignum register index d comes from
                                            // base register b read using d in this struct

    logic                    d_inc;           // Increment destination register index in base
                                              // register file
    logic                    a_inc;           // Increment source register index a in base register
                                              // file
    logic                    a_wlen_word_inc; // Increment source register a in base register file
                                              // by WLEN word size
    logic                    b_inc;           // Increment source register index b in base register
                                              // file

    // Shifting only applies to a subset of ALU operations
    logic [$clog2(WLEN)-1:0] alu_shift_amt;   // Shift amount
    logic                    alu_shift_right; // Shift right if set otherwise left

    flag_group_t             alu_flag_group;
    flag_e                   alu_sel_flag;
    logic                    alu_flag_en;
    logic                    mac_flag_en;
    alu_op_bignum_e          alu_op;
    op_b_sel_e               alu_op_b_sel;

    logic [1:0]              mac_op_a_qw_sel;
    logic [1:0]              mac_op_b_qw_sel;
    logic                    mac_wr_hw_sel_upper;
    logic [1:0]              mac_pre_acc_shift;
    logic                    mac_zero_acc;
    logic                    mac_shift_out;
    logic                    mac_en;

    logic                    rf_we;
    rf_wd_sel_e              rf_wdata_sel;
    logic                    rf_ren_a;
    logic                    rf_ren_b;

    logic                    sel_insn;
  } insn_dec_bignum_t;

  typedef struct packed {
    logic [NWdr-1:0] rf_ren_a;
    logic [NWdr-1:0] rf_ren_b;
    logic [NWdr-1:0] rf_we;
  } rf_predec_bignum_t;

  typedef struct packed {
    logic                    adder_x_en;
    logic                    x_res_operand_a_sel;
    logic                    adder_y_op_a_en;
    logic                    shift_mod_sel;
    logic                    adder_y_op_shifter_en;
    logic                    shifter_a_en;
    logic                    shifter_b_en;
    logic                    shift_right;
    logic [$clog2(WLEN)-1:0] shift_amt;
    logic                    logic_a_en;
    logic                    logic_shifter_en;
    logic [3:0]              logic_res_sel;
    logic [NFlagGroups-1:0]  flag_group_sel;
    flags_t                  flag_sel;
    logic [NFlagGroups-1:0]  flags_keep;
    logic [NFlagGroups-1:0]  flags_adder_update;
    logic [NFlagGroups-1:0]  flags_logic_update;
    logic [NFlagGroups-1:0]  flags_mac_update;
    logic [NFlagGroups-1:0]  flags_ispr_wr;
  } alu_predec_bignum_t;

  typedef struct packed {
    logic [NIspr-1:0] ispr_rd_en;
    logic [NIspr-1:0] ispr_wr_en;
  } ispr_predec_bignum_t;

  typedef struct packed {
    logic op_en;
    logic acc_rd_en;
  } mac_predec_bignum_t;

  typedef struct packed {
    logic call_stack_pop;
    logic call_stack_push;
    logic branch_insn;
    logic jump_insn;
    logic loop_insn;
    logic sel_insn;
  } ctrl_flow_predec_t;

  typedef struct packed {
    alu_op_base_e     op;
    logic [31:0] operand_a;
    logic [31:0] operand_b;
  } alu_base_operation_t;

  typedef struct packed {
    comparison_op_base_e op;
    logic [31:0] operand_a;
    logic [31:0] operand_b;
  } alu_base_comparison_t;

  typedef struct packed {
    alu_op_bignum_e op;
    logic [WLEN-1:0]         operand_a;
    logic [WLEN-1:0]         operand_b;
    logic                    shift_right;
    logic [$clog2(WLEN)-1:0] shift_amt;
    flag_group_t             flag_group;
    flag_e                   sel_flag;
    logic                    alu_flag_en;
    logic                    mac_flag_en;
  } alu_bignum_operation_t;

  typedef struct packed {
    logic [WLEN-1:0] operand_a;
    logic [WLEN-1:0] operand_b;
    logic [1:0]      operand_a_qw_sel;
    logic [1:0]      operand_b_qw_sel;
    logic            wr_hw_sel_upper;
    logic [1:0]      pre_acc_shift_imm;
    logic            zero_acc;
    logic            shift_acc;
  } mac_bignum_operation_t;

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 5 \
  //      -s 5799399942 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (66.67%)
  //  4: |||||||||| (33.33%)
  //  5: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4

  localparam int StateControllerWidth = 5;
  typedef enum logic [StateControllerWidth-1:0] {
    OtbnStateHalt        = 5'b00100,
    OtbnStateRun         = 5'b01010,
    OtbnStateStall       = 5'b10011,
    OtbnStateLocked      = 5'b11101
  } otbn_state_e;

  // States for start_stop_controller
  // Encoding generated with:
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 9 -n 7 \
  //      -s 573771984 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (44.44%)
  //  4: |||||||||||||||||| (41.67%)
  //  5: | (2.78%)
  //  6: | (2.78%)
  //  7: ||| (8.33%)
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 7
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 6
  //
  localparam int StateStartStopWidth = 7;
  typedef enum logic [StateStartStopWidth-1:0] {
    OtbnStartStopStateInitial             = 7'b1010011,
    OtbnStartStopStateHalt                = 7'b1111001,
    OtbnStartStopStateUrndRefresh         = 7'b0000110,
    OtbnStartStopStateRunning             = 7'b1001000,
    OtbnStartStopSecureWipeWdrUrnd        = 7'b0101100,
    OtbnStartStopSecureWipeAccModBaseUrnd = 7'b0010000,
    OtbnStartStopSecureWipeAllZero        = 7'b0110101,
    OtbnStartStopSecureWipeComplete       = 7'b0001011,
    OtbnStartStopStateLocked              = 7'b1101111
  } otbn_start_stop_state_e;

// Encoding generated with:
// $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 5 \
//      -s 2298830978 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (66.67%)
//  4: |||||||||| (33.33%)
//  5: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 4
// Minimum Hamming weight: 1
// Maximum Hamming weight: 4
//
localparam int StateScrambleCtrlWidth = 5;
typedef enum logic [StateScrambleCtrlWidth-1:0] {
  ScrambleCtrlIdle    = 5'b10011,
  ScrambleCtrlDmemReq = 5'b11110,
  ScrambleCtrlImemReq = 5'b01000,
  ScrambleCtrlError   = 5'b00101
} scramble_ctrl_state_e;

  // URNG PRNG default seed.
  // These parameters have been generated with
  // $ ./util/design/gen-lfsr-seed.py --width 256 --seed 2840984437 --prefix "Urnd"
  parameter int UrndPrngWidth = 256;
  typedef logic [UrndPrngWidth-1:0] urnd_prng_seed_t;
  parameter urnd_prng_seed_t RndCnstUrndPrngSeedDefault =
      256'h84ddfadaf7e1134d70aa1c59de6197ff25a4fe335d095f1e2cba89acbe4a07e9;

  parameter otp_ctrl_pkg::otbn_key_t RndCnstOtbnKeyDefault =
      128'h14e8cecae3040d5e12286bb3cc113298;
  parameter otp_ctrl_pkg::otbn_nonce_t RndCnstOtbnNonceDefault =
      64'hf79780bc735f3843;

  typedef logic [63:0] otbn_dmem_nonce_t;
  typedef logic [63:0] otbn_imem_nonce_t;
endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Common Library: Clock Gating cell with synchronizer

module prim_clock_gating_sync (
  input        clk_i,
  input        rst_ni,
  input        test_en_i,
  input        async_en_i,
  output logic en_o,
  output logic clk_o
);


  prim_flop_2sync #(
    .Width(1)
  ) i_sync (
    .clk_i,
    .rst_ni,
    .d_i(async_en_i),
    .q_o(en_o)
  );

  prim_clock_gating i_cg (
    .clk_i,
    .en_i(en_o),
    .test_en_i,
    .clk_o
  );


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// N:1 SRAM arbiter
//
// Parameter
//  N:  Number of requst port
//  DW: Data width (SECDED is not included)
//  Aw: Address width
//  ArbiterImpl: can be either PPC or BINTREE.
`include "prim_assert.sv"

module prim_sram_arbiter #(
  parameter int unsigned N  = 4,
  parameter int unsigned SramDw = 32,
  parameter int unsigned SramAw = 12,
  parameter ArbiterImpl = "PPC",
  parameter bit EnMask = 1'b 0 // Disable wmask if 0
) (
  input clk_i,
  input rst_ni,

  input        [     N-1:0] req_i,
  input        [SramAw-1:0] req_addr_i [N],
  input        [     N-1:0] req_write_i,
  input        [SramDw-1:0] req_wdata_i[N],
  input        [SramDw-1:0] req_wmask_i[N],
  output logic [     N-1:0] gnt_o,

  output logic [     N-1:0] rsp_rvalid_o,      // Pulse
  output logic [SramDw-1:0] rsp_rdata_o[N],
  output logic [       1:0] rsp_error_o[N],

  // SRAM Interface
  output logic              sram_req_o,
  output logic [SramAw-1:0] sram_addr_o,
  output logic              sram_write_o,
  output logic [SramDw-1:0] sram_wdata_o,
  output logic [SramDw-1:0] sram_wmask_o,
  input                     sram_rvalid_i,
  input        [SramDw-1:0] sram_rdata_i,
  input        [1:0]        sram_rerror_i
);

  typedef struct packed {
    logic write;
    logic [SramAw-1:0] addr;
    logic [SramDw-1:0] wdata;
    logic [SramDw-1:0] wmask;
  } req_t;

  req_t req_packed [N];

  for (genvar i = 0 ; i < N ; i++) begin : gen_reqs
    assign req_packed[i] = {
      req_write_i[i],
      req_addr_i [i],
      req_wdata_i[i],
      (EnMask) ? req_wmask_i[i] : {SramDw{1'b1}}
    };
  end

  localparam int ARB_DW = $bits(req_t);

  req_t sram_packed;
  assign sram_write_o = sram_packed.write;
  assign sram_addr_o  = sram_packed.addr;
  assign sram_wdata_o = sram_packed.wdata;
  assign sram_wmask_o = (EnMask) ? sram_packed.wmask : {SramDw{1'b1}};

  if (EnMask == 1'b 0) begin : g_unused
    logic unused_wmask;

    always_comb begin
      unused_wmask = 1'b 1;
      for (int unsigned i = 0 ; i < N ; i++) begin
        unused_wmask ^= ^req_wmask_i[i];
      end
      unused_wmask ^= ^sram_packed.wmask;
    end
  end


  if (ArbiterImpl == "PPC") begin : gen_arb_ppc
    prim_arbiter_ppc #(
      .N (N),
      .DW(ARB_DW)
    ) u_reqarb (
      .clk_i,
      .rst_ni,
      .req_chk_i ( 1'b1        ),
      .req_i,
      .data_i    ( req_packed  ),
      .gnt_o,
      .idx_o     (             ),
      .valid_o   ( sram_req_o  ),
      .data_o    ( sram_packed ),
      .ready_i   ( 1'b1        )
    );
  end else if (ArbiterImpl == "BINTREE") begin : gen_tree_arb
    prim_arbiter_tree #(
      .N (N),
      .DW(ARB_DW)
    ) u_reqarb (
      .clk_i,
      .rst_ni,
      .req_chk_i ( 1'b1        ),
      .req_i,
      .data_i    ( req_packed  ),
      .gnt_o,
      .idx_o     (             ),
      .valid_o   ( sram_req_o  ),
      .data_o    ( sram_packed ),
      .ready_i   ( 1'b1        )
    );
  end else begin : gen_unknown
    `ASSERT_INIT(UnknownArbImpl_A, 0)
  end


  logic [N-1:0] steer;    // Steering sram_rvalid_i
  logic sram_ack;         // Ack for rvalid. |sram_rvalid_i

  assign sram_ack = sram_rvalid_i & (|steer);

  // Request FIFO
  prim_fifo_sync #(
    .Width    (N),
    .Pass     (1'b0),
    .Depth    (4)        // Assume at most 4 pipelined
  ) u_req_fifo (
    .clk_i,
    .rst_ni,
    .clr_i    (1'b0),
    .wvalid_i (sram_req_o & ~sram_write_o),  // Push only for read
    .wready_o (),     // TODO: Generate Error
    .wdata_i  (gnt_o),
    .rvalid_o (),     // TODO; Generate error if sram_rvalid_i but rvalid==0
    .rready_i (sram_ack),
    .rdata_o  (steer),
    .full_o   (),
    .depth_o  (),     // Not used
    .err_o    ()
  );

  assign rsp_rvalid_o = steer & {N{sram_rvalid_i}};

  for (genvar i = 0 ; i < N ; i++) begin : gen_rsp
    assign rsp_rdata_o[i] = sram_rdata_i;
    assign rsp_error_o[i] = sram_rerror_i; // No SECDED yet
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Slicer chops the incoming bitstring into OutW granularity.
// It supports fractional InW/OutW which fills 0 at the end of message.

`include "prim_assert.sv"

module prim_slicer #(
  parameter int InW = 64,
  parameter int OutW = 8,

  parameter int IndexW = 4
) (
  input        [IndexW-1:0] sel_i,
  input        [InW-1:0]    data_i,
  output logic [OutW-1:0]   data_o
);

  localparam int UnrollW = OutW*(2**IndexW);

  logic [UnrollW-1:0] unrolled_data;

  assign unrolled_data = UnrollW'(data_i);

  assign data_o = unrolled_data[sel_i*OutW+:OutW];

  `ASSERT_INIT(ValidWidth_A, InW <= OutW*(2**IndexW))

endmodule



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// REQ/ACK synchronizer
//
// This module synchronizes a REQ/ACK handshake across a clock domain crossing.
// Both domains will see a handshake with the duration of one clock cycle.
//
// Notes:
// - Once asserted, the source (SRC) domain is not allowed to de-assert REQ without ACK.
// - The destination (DST) domain is not allowed to send an ACK without a REQ.
// - When resetting one domain, also the other domain needs to be reset with both resets being
//   active at the same time.
// - This module works both when syncing from a faster to a slower clock domain and vice versa.
// - Internally, this module uses a non-return-to-zero (NRZ), two-phase handshake protocol by
//   default. Assuming the DST domain responds with an ACK immediately, the latency from asserting
//   the REQ in the SRC domain is:
//   - 1 source + 2 destination clock cycles until the handshake is performed in the DST domain,
//   - 1 source + 2 destination + 1 destination + 2 source clock cycles until the handshake is
//     performed in the SRC domain.
// - Optionally, the module can also use a return-to-zero (RZ), four-phase handshake protocol.
//   That one has lower throughput, but it is safe to partially reset either side, since the
//   two FSMs cannot get out of sync due to persisting EVEN/ODD states. The handshake latencies
//   are the same as for the NRZ protocol, but the throughput is half that of the NRZ protocol
//   since the signals neet to return to zero first, causing two round-trips through the
//   synchronizers instead of just one.
//
// For further information, see Section 8.2.4 in H. Kaeslin, "Top-Down Digital VLSI Design: From
// Architecture to Gate-Level Circuits and FPGAs", 2015.

`include "prim_assert.sv"

module prim_sync_reqack #(
  parameter bit EnRstChks = 1'b0,   // Enable reset-related assertion checks, disabled by default.
  parameter bit EnRzHs = 1'b0       // By Default, the faster NRZ handshake protocol
                                    // (EnRzHs = 0) is used. Enable the RZ handshake protocol
                                    // if the FSMs need to be partial-reset-safe.
) (
  input  clk_src_i,       // REQ side, SRC domain
  input  rst_src_ni,      // REQ side, SRC domain
  input  clk_dst_i,       // ACK side, DST domain
  input  rst_dst_ni,      // ACK side, DST domain

  input  logic req_chk_i, // Used for gating assertions. Drive to 1 during normal operation.

  input  logic src_req_i, // REQ side, SRC domain
  output logic src_ack_o, // REQ side, SRC domain
  output logic dst_req_o, // ACK side, DST domain
  input  logic dst_ack_i  // ACK side, DST domain
);

  // req_chk_i is used for gating assertions only.
  logic unused_req_chk;
  assign unused_req_chk = req_chk_i;

  if (EnRzHs) begin : gen_rz_hs_protocol
    //////////////////
    // RZ protocol //
    //////////////////

    // Types
    typedef enum logic {
      LoSt, HiSt
    } rz_fsm_e;

    // Signals
    rz_fsm_e src_fsm_d, src_fsm_q;
    rz_fsm_e dst_fsm_d, dst_fsm_q;
    logic src_ack, dst_ack;
    logic src_req, dst_req;

    // REQ-side FSM (SRC domain)
    always_comb begin : src_fsm
      src_fsm_d = src_fsm_q;
      src_ack_o = 1'b0;
      src_req = 1'b0;

      unique case (src_fsm_q)
        LoSt: begin
          // Wait for the ack to go back to zero before starting
          // a new transaction.
          if (!src_ack && src_req_i) begin
            src_fsm_d = HiSt;
          end
        end
        HiSt: begin
          src_req = 1'b1;
          // Forward the acknowledgement.
          src_ack_o = src_ack;
          // If request drops out, we go back to LoSt.
          // If DST side asserts ack, we also go back to LoSt.
          if (!src_req_i || src_ack) begin
            src_fsm_d = LoSt;
          end
        end
        //VCS coverage off
        // pragma coverage off
        default: ;
        //VCS coverage on
        // pragma coverage on
      endcase
    end

    // Move ACK over to SRC domain.
    prim_flop_2sync #(
      .Width(1)
    ) ack_sync (
      .clk_i  (clk_src_i),
      .rst_ni (rst_src_ni),
      .d_i    (dst_ack),
      .q_o    (src_ack)
    );

    // Registers
    always_ff @(posedge clk_src_i or negedge rst_src_ni) begin
      if (!rst_src_ni) begin
        src_fsm_q <= LoSt;
      end else begin
        src_fsm_q <= src_fsm_d;
      end
    end

    // ACK-side FSM (DST domain)
    always_comb begin : dst_fsm
      dst_fsm_d = dst_fsm_q;
      dst_req_o = 1'b0;
      dst_ack = 1'b0;

      unique case (dst_fsm_q)
        LoSt: begin
          if (dst_req) begin
            // Forward the request.
            dst_req_o = 1'b1;
            // Wait for the request and acknowledge to be asserted
            // before responding to the SRC side.
            if (dst_ack_i) begin
              dst_fsm_d = HiSt;
            end
          end
        end
        HiSt: begin
          dst_ack = 1'b1;
          // Wait for the request to drop back to zero.
          if (!dst_req) begin
            dst_fsm_d = LoSt;
          end
        end
        //VCS coverage off
        // pragma coverage off
        default: ;
        //VCS coverage on
        // pragma coverage on
      endcase
    end

    // Move REQ over to DST domain.
    prim_flop_2sync #(
      .Width(1)
    ) req_sync (
      .clk_i  (clk_dst_i),
      .rst_ni (rst_dst_ni),
      .d_i    (src_req),
      .q_o    (dst_req)
    );

    // Registers
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        dst_fsm_q <= LoSt;
      end else begin
        dst_fsm_q <= dst_fsm_d;
      end
    end

  end else begin : gen_nrz_hs_protocol
    //////////////////
    // NRZ protocol //
    //////////////////

    // Types
    typedef enum logic {
      EVEN, ODD
    } sync_reqack_fsm_e;

    // Signals
    sync_reqack_fsm_e src_fsm_ns, src_fsm_cs;
    sync_reqack_fsm_e dst_fsm_ns, dst_fsm_cs;

    logic src_req_d, src_req_q, src_ack;
    logic dst_ack_d, dst_ack_q, dst_req;
    logic src_handshake, dst_handshake;

    assign src_handshake = src_req_i & src_ack_o;
    assign dst_handshake = dst_req_o & dst_ack_i;

    // Move REQ over to DST domain.
    prim_flop_2sync #(
      .Width(1)
    ) req_sync (
      .clk_i  (clk_dst_i),
      .rst_ni (rst_dst_ni),
      .d_i    (src_req_q),
      .q_o    (dst_req)
    );

    // Move ACK over to SRC domain.
    prim_flop_2sync #(
      .Width(1)
    ) ack_sync (
      .clk_i  (clk_src_i),
      .rst_ni (rst_src_ni),
      .d_i    (dst_ack_q),
      .q_o    (src_ack)
    );

    // REQ-side FSM (SRC domain)
    always_comb begin : src_fsm
      src_fsm_ns = src_fsm_cs;

      // By default, we keep the internal REQ value and don't ACK.
      src_req_d = src_req_q;
      src_ack_o = 1'b0;

      unique case (src_fsm_cs)

        EVEN: begin
          // Simply forward REQ and ACK.
          src_req_d = src_req_i;
          src_ack_o = src_ack;

          // The handshake is done for exactly 1 clock cycle.
          if (src_handshake) begin
            src_fsm_ns = ODD;
          end
        end

        ODD: begin
          // Internal REQ and ACK have inverted meaning now. If src_req_i is high again, this
          // signals a new transaction.
          src_req_d = ~src_req_i;
          src_ack_o = ~src_ack;

          // The handshake is done for exactly 1 clock cycle.
          if (src_handshake) begin
            src_fsm_ns = EVEN;
          end
        end

        //VCS coverage off
        // pragma coverage off

        default: ;

        //VCS coverage on
        // pragma coverage on

      endcase
    end

    // ACK-side FSM (DST domain)
    always_comb begin : dst_fsm
      dst_fsm_ns = dst_fsm_cs;

      // By default, we don't REQ and keep the internal ACK.
      dst_req_o = 1'b0;
      dst_ack_d = dst_ack_q;

      unique case (dst_fsm_cs)

        EVEN: begin
          // Simply forward REQ and ACK.
          dst_req_o = dst_req;
          dst_ack_d = dst_ack_i;

          // The handshake is done for exactly 1 clock cycle.
          if (dst_handshake) begin
            dst_fsm_ns = ODD;
          end
        end

        ODD: begin
          // Internal REQ and ACK have inverted meaning now. If dst_req goes low, this signals a new
          // transaction.
          dst_req_o = ~dst_req;
          dst_ack_d = ~dst_ack_i;

          // The handshake is done for exactly 1 clock cycle.
          if (dst_handshake) begin
            dst_fsm_ns = EVEN;
          end
        end

        //VCS coverage off
        // pragma coverage off

        default: ;

        //VCS coverage on
        // pragma coverage on

      endcase
    end

    // Registers
    always_ff @(posedge clk_src_i or negedge rst_src_ni) begin
      if (!rst_src_ni) begin
        src_fsm_cs <= EVEN;
        src_req_q  <= 1'b0;
      end else begin
        src_fsm_cs <= src_fsm_ns;
        src_req_q  <= src_req_d;
      end
    end
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        dst_fsm_cs <= EVEN;
        dst_ack_q  <= 1'b0;
      end else begin
        dst_fsm_cs <= dst_fsm_ns;
        dst_ack_q  <= dst_ack_d;
      end
    end
  end

  ////////////////
  // Assertions //
  ////////////////

  `ifdef INC_ASSERT
    //VCS coverage off
    // pragma coverage off

    logic effective_rst_n;
    assign effective_rst_n = rst_src_ni && rst_dst_ni;

    logic chk_flag;
    always_ff @(posedge clk_src_i or negedge effective_rst_n) begin
      if (!effective_rst_n) begin
        chk_flag <= '0;
      end else if (src_req_i && !chk_flag) begin
        chk_flag <= 1'b1;
      end
    end
    //VCS coverage on
    // pragma coverage on

    // SRC domain can only de-assert REQ after receiving ACK.
    `ASSERT(SyncReqAckHoldReq, $fell(src_req_i) && req_chk_i && chk_flag |->
        $fell(src_ack_o), clk_src_i, !rst_src_ni || !rst_dst_ni || !req_chk_i || !chk_flag)
  `endif

  // DST domain cannot assert ACK without REQ.
  `ASSERT(SyncReqAckAckNeedsReq, dst_ack_i |->
      dst_req_o, clk_dst_i, !rst_src_ni || !rst_dst_ni)

  if (EnRstChks) begin : gen_assert_en_rst_chks
  `ifdef INC_ASSERT

    //VCS coverage off
    // pragma coverage off
    // This assertion is written very oddly because it is difficult to reliably catch
    // when rst drops.
    // The problem is that reset assertion in the design is often associated with clocks
    // stopping, this means things like rise / fell don't work correctly since there are
    // no clocks.
    // As a result of this, we end up detecting way past the interest point (whenever
    // clocks are restored) and falsely assert an error.
    // The code below instead tries to use asynchronous flags to determine when and if
    // the two domains are properly reset.
    logic src_reset_flag;
    always_ff @(posedge clk_src_i or negedge rst_src_ni) begin
      if (!rst_src_ni) begin
        src_reset_flag <= '0;
      end else if(src_req_i) begin
        src_reset_flag <= 1'b1;
      end
    end

    logic dst_reset_flag;
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        dst_reset_flag <= '0;
      end else if (dst_req_o) begin
        dst_reset_flag <= 1'b1;
      end
    end
    //VCS coverage on
    // pragma coverage on

    // Always reset both domains. Both resets need to be active at the same time.
    `ASSERT(SyncReqAckRstSrc, $fell(rst_src_ni) |->
        (!src_reset_flag throughout !dst_reset_flag[->1]),
        clk_src_i, 0)
    `ASSERT(SyncReqAckRstDst, $fell(rst_dst_ni) |->
        (!dst_reset_flag throughout !src_reset_flag[->1]),
        clk_dst_i, 0)

  `endif


  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// REQ/ACK synchronizer with associated data.
//
// This module synchronizes a REQ/ACK handshake with associated data across a clock domain
// crossing (CDC). Both domains will see a handshake with the duration of one clock cycle. By
// default, the data itself is not registered. The main purpose of feeding the data through this
// module to have an anchor point for waiving CDC violations. If the data is configured to flow
// from the destination (DST) to the source (SRC) domain, an additional register stage can be
// inserted for data buffering.
//
// Under the hood, this module uses a prim_sync_reqack primitive for synchronizing the
// REQ/ACK handshake. See prim_sync_reqack.sv for more details.

`include "prim_assert.sv"

module prim_sync_reqack_data #(
  parameter int unsigned Width       = 1,
  parameter bit          EnRstChks   = 1'b0, // Enable reset-related assertion checks, disabled by
                                             // default.
  parameter bit          DataSrc2Dst = 1'b1, // Direction of data flow: 1'b1 = SRC to DST,
                                             //                         1'b0 = DST to SRC
  parameter bit          DataReg     = 1'b0, // Enable optional register stage for data,
                                             // only usable with DataSrc2Dst == 1'b0.
  parameter bit          EnRzHs      = 1'b0  // By Default, we the faster NRZ handshake protocol
                                             // (EnRzHs = 0) is used. Enable the RZ handshake
                                             // protocol if the FSMs need to be partial-reset-safe.
) (
  input  clk_src_i,       // REQ side, SRC domain
  input  rst_src_ni,      // REQ side, SRC domain
  input  clk_dst_i,       // ACK side, DST domain
  input  rst_dst_ni,      // ACK side, DST domain

  input  logic req_chk_i, // Used for gating assertions. Drive to 1 during normal operation.

  input  logic src_req_i, // REQ side, SRC domain
  output logic src_ack_o, // REQ side, SRC domain
  output logic dst_req_o, // ACK side, DST domain
  input  logic dst_ack_i, // ACK side, DST domain

  input  logic [Width-1:0] data_i,
  output logic [Width-1:0] data_o
);

  ////////////////////////////////////
  // REQ/ACK synchronizer primitive //
  ////////////////////////////////////
  prim_sync_reqack #(
    .EnRstChks(EnRstChks),
    .EnRzHs(EnRzHs)
  ) u_prim_sync_reqack (
    .clk_src_i,
    .rst_src_ni,
    .clk_dst_i,
    .rst_dst_ni,

    .req_chk_i,

    .src_req_i,
    .src_ack_o,
    .dst_req_o,
    .dst_ack_i
  );

  /////////////////////////
  // Data register stage //
  /////////////////////////
  // Optional - Only relevant if the data flows from DST to SRC. In this case, it must be ensured
  // that the data remains stable until the ACK becomes visible in the SRC domain.
  //
  // Note that for larger data widths, it is recommended to adjust the data sender to hold the data
  // stable until the next REQ in order to save the cost of this register stage.
  if (DataSrc2Dst == 1'b0 && DataReg == 1'b1) begin : gen_data_reg
    logic             data_we;
    logic [Width-1:0] data_d, data_q;

    // Sample the data when seing the REQ/ACK handshake in the DST domain.
    assign data_we = dst_req_o & dst_ack_i;
    assign data_d  = data_i;
    always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
      if (!rst_dst_ni) begin
        data_q <= '0;
      end else if (data_we) begin
        data_q <= data_d;
      end
    end
    assign data_o = data_q;

  end else begin : gen_no_data_reg
    // Just feed through the data.
    assign data_o = data_i;
  end

  ////////////////
  // Assertions //
  ////////////////
  if (DataSrc2Dst == 1'b1) begin : gen_assert_data_src2dst
`ifdef INC_ASSERT
    //VCS coverage off
    // pragma coverage off
    logic effective_rst_n;
    assign effective_rst_n = rst_src_ni && rst_dst_ni;

    logic chk_flag_d, chk_flag_q;
    assign chk_flag_d = src_req_i && !chk_flag_q ? 1'b1 : chk_flag_q;

    always_ff @(posedge clk_src_i or negedge effective_rst_n) begin
      if (!effective_rst_n) begin
        chk_flag_q <= '0;
      end else begin
        chk_flag_q <= chk_flag_d;
      end
    end
    //VCS coverage on
    // pragma coverage on

    // SRC domain cannot change data while waiting for ACK.
    `ASSERT(SyncReqAckDataHoldSrc2Dst, !$stable(data_i) && chk_flag_q |->
        (!src_req_i || (src_req_i && src_ack_o)),
        clk_src_i, !rst_src_ni || !rst_dst_ni || !chk_flag_q)

    // Register stage cannot be used.
    `ASSERT_INIT(SyncReqAckDataReg, DataSrc2Dst && !DataReg)
`endif
  end else if (DataSrc2Dst == 1'b0 && DataReg == 1'b0) begin : gen_assert_data_dst2src
    // DST domain shall not change data while waiting for SRC domain to latch it (together with
    // receiving ACK). It takes 2 SRC cycles for ACK to cross over from DST to SRC, and 1 SRC cycle
    // for the next REQ to cross over from SRC to DST.
    //
    // Denote the src clock where REQ & ACK as time zero. The data flowing through the CDC could be
    // corrupted if data_o was not stable over the previous 2 clock cycles (so we want to check time
    // points -2, -1 and 0). Moreover, the DST domain cannot know that it is allowed to change value
    // until at least one more SRC cycle (the time taken for REQ to cross back from SRC to DST).
    //
    // To make this assertion, we will sample at each of 4 time points (-2, -1, 0 and +1), asserting
    // that data_o is equal at each of these times. Note this won't detect glitches at intermediate
    // timepoints.
    //
    // The SVAs below are designed not to consume time, which means that they can be disabled with
    // an $assertoff(..) and won't linger to fail later. This wouldn't work properly if we used
    // something like |=> instead of the $past(...) function. That means that we have to trigger at
    // the "end" of the window. To make sure we don't miss a situation where the value changed at
    // time -1 (causing corruption), but reset was asserted between time 0 and 1, we split the
    // assertion into two pieces. The first (SyncReqAckDataHoldDst2SrcA) checks that data doesn't
    // change in a way that could cause data corruption. The second (SyncReqAckDataHoldDst2SrcB)
    // checks that the DST side doesn't do anything that it shouldn't know is safe.
`ifdef INC_ASSERT
    //VCS coverage off
    // pragma coverage off
    logic effective_rst_n;
    assign effective_rst_n = rst_src_ni && rst_dst_ni;

    logic chk_flag_d, chk_flag_q;
    assign chk_flag_d = src_req_i && !chk_flag_q ? 1'b1 : chk_flag_q;

    always_ff @(posedge clk_src_i or negedge effective_rst_n) begin
      if (!effective_rst_n) begin
        chk_flag_q <= '0;
      end else begin
        chk_flag_q <= chk_flag_d;
      end
    end
    //VCS coverage on
    // pragma coverage on

    `ASSERT(SyncReqAckDataHoldDst2SrcA,
            chk_flag_q && src_req_i && src_ack_o |->
            $past(data_o, 2) == data_o && $past(data_o) == data_o,
            clk_src_i, !rst_src_ni || !rst_dst_ni || !chk_flag_q)
    `ASSERT(SyncReqAckDataHoldDst2SrcB,
            chk_flag_q && $past(src_req_i && src_ack_o) |-> $past(data_o) == data_o,
            clk_src_i, !rst_src_ni || !rst_dst_ni || !chk_flag_q)
`endif
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Slow to fast clock synchronizer
// This module is designed to be used for efficient sampling of signals from a slow clock to a much
// faster clock.
//
// The data is captured into flops on the negative edge of the slow clock (when the data should be
// stable). Because the slow clock passes through a two-flop synchronizer, the ratio of clock speeds
// needs to be high to guarantee that the data will be stable when sampled.
//
// A ratio of at-least 10:1 in clock speeds is recommended.

module prim_sync_slow_fast #(
  parameter int unsigned Width = 32
) (
  input  logic             clk_slow_i,
  input  logic             clk_fast_i,
  input  logic             rst_fast_ni,
  input  logic [Width-1:0] wdata_i,    // Slow domain
  output logic [Width-1:0] rdata_o     // Fast domain
);

  logic             sync_clk_slow, sync_clk_slow_q;
  logic             wdata_en;
  logic [Width-1:0] wdata_q;

  // Synchronize the slow clock to the fast domain
  prim_flop_2sync #(.Width(1)) sync_slow_clk (
    .clk_i    (clk_fast_i),
    .rst_ni   (rst_fast_ni),
    .d_i      (clk_slow_i),
    .q_o      (sync_clk_slow));

  // Register the synchronized clk
  always_ff @(posedge clk_fast_i or negedge rst_fast_ni) begin
    if (!rst_fast_ni) begin
      sync_clk_slow_q <= 1'b0;
    end else begin
      sync_clk_slow_q <= sync_clk_slow;
    end
  end

  // Find the negative edge of the synchronized slow clk
  assign wdata_en = sync_clk_slow_q & !sync_clk_slow;

  // Sample the slow data on the negative edge
  always_ff @(posedge clk_fast_i or negedge rst_fast_ni) begin
    if (!rst_fast_ni) begin
      wdata_q <= '0;
    end else if (wdata_en) begin
      wdata_q <= wdata_i;
    end
  end

  assign rdata_o = wdata_q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// prim_keccak is single round permutation module
`include "prim_assert.sv"
module prim_keccak #(
  parameter int Width = 1600, // b= {25, 50, 100, 200, 400, 800, 1600}

  // Derived
  localparam int W        = Width/25,
  localparam int L        = $clog2(W),
  localparam int MaxRound = 12 + 2*L, // Keccak-f only
  localparam int RndW     = $clog2(MaxRound+1) // Representing up to MaxRound
) (
  input        [RndW-1:0]  rnd_i,   // Current Round
  input        [Width-1:0] s_i,
  output logic [Width-1:0] s_o
);
  ///////////
  // Types //
  ///////////
  //             x    y    z
  typedef logic [4:0][4:0][W-1:0] box_t;   // (x,y,z) state
  typedef logic           [W-1:0] lane_t;  // (z)
  typedef logic [4:0]     [W-1:0] plane_t; // (x,z)
  typedef logic [4:0][4:0]        slice_t; // (x,y)
  typedef logic      [4:0][W-1:0] sheet_t; // (y,z) identical to plane_t
  typedef logic [4:0]             row_t;   // (x)
  typedef logic      [4:0]        col_t;   // (y) identical to row_t

  //////////////
  // Keccak_f //
  //////////////
  box_t state_in, keccak_f;
  box_t theta_data, rho_data, pi_data, chi_data, iota_data;
  assign state_in = bitarray_to_box(s_i);
  assign theta_data = theta(state_in);
  // Commented out rho function as vcs complains z-Offset%W isn't constant
  //assign rho_data   = rho(theta_data);
  assign pi_data    = pi(rho_data);
  assign chi_data   = chi(pi_data);
  assign iota_data  = iota(chi_data, rnd_i);
  assign keccak_f   = iota_data;
  assign s_o        = box_to_bitarray(keccak_f);

  // Rho ======================================================================
  // As RhoOffset[x][y] is considered as variable int in VCS,
  // it is replaced with generate statement.
  localparam int RhoOffset [5][5]  = '{
    //y  0    1    2    3    4     x
    '{   0,  36,   3, 105, 210},// 0
    '{   1, 300,  10,  45,  66},// 1
    '{ 190,   6, 171,  15, 253},// 2
    '{  28,  55, 153,  21, 120},// 3
    '{  91, 276, 231, 136,  78} // 4
  };
  for (genvar x = 0 ; x < 5 ; x++) begin : gen_rho_x
    for (genvar y = 0 ; y < 5 ; y++) begin : gen_rho_y
      localparam int Offset = RhoOffset[x][y]%W;
      localparam int ShiftAmt = W- Offset;
      if (Offset == 0) begin : gen_offset0
        assign rho_data[x][y][W-1:0] = theta_data[x][y][W-1:0];
      end else begin : gen_others
        assign rho_data[x][y][W-1:0] = {theta_data[x][y][0+:ShiftAmt],
                                        theta_data[x][y][ShiftAmt+:Offset]};
      end
    end
  end

  ////////////////
  // Assertions //
  ////////////////

  `ASSERT_INIT(ValidWidth_A, Width inside {25, 50, 100, 200, 400, 800, 1600})
  `ASSERT_INIT(ValidW_A, W inside {1, 2, 4, 8, 16, 32, 64})
  `ASSERT_INIT(ValidL_A, L inside {0, 1, 2, 3, 4, 5, 6})
  `ASSERT_INIT(ValidRound_A, MaxRound <= 24) // Keccak-f only

  ///////////////
  // Functions //
  ///////////////

  // Convert bitarray to 3D box
  // Please take a look at FIPS PUB 202
  // https://nvlpubs.nist.gov/nistpubs/FIPS/NIST.FIPS.202.pdf
  // > For all triples (x,y,z) such that 0<=x<5, 0<=y<5, and 0<=z<w,
  // >    A[x,y,z]=S[w(5y+x)+z]
  function automatic box_t bitarray_to_box(logic [Width-1:0] s_in);
    automatic box_t box;
    for (int y = 0 ; y < 5 ; y++) begin
      for (int x = 0 ; x < 5 ; x++) begin
        for (int z = 0 ; z < W ; z++) begin
          box[x][y][z] = s_in[W*(5*y+x) + z];
        end
      end
    end
    return box;
  endfunction : bitarray_to_box

  // Convert 3D cube to bitarray
  function automatic logic [Width-1:0] box_to_bitarray(box_t state);
    automatic logic [Width-1:0] bitarray;
    for (int y = 0 ; y < 5 ; y++) begin
      for (int x = 0 ; x < 5 ; x++) begin
        for (int z = 0 ; z < W ; z++) begin
          bitarray[W*(5*y+x)+z] = state[x][y][z];
        end
      end
    end
    return bitarray;
  endfunction : box_to_bitarray

  // Step Mapping =============================================================
  // theta
  // XOR each bit in the state with the parity of two columns
  // C[x,z] = A[x,0,z] ^ A[x,1,z] ^ A[x,2,z] ^ A[x,3,z] ^ A[x,4,z]
  // D[x,z] = C[x-1,z] ^ C[x+1,z-1]
  // theta = A[x,y,z] ^ D[x,z]
  function automatic box_t theta(box_t state);
    plane_t c;
    plane_t d;
    box_t result;
    for (int x = 0 ; x < 5 ; x++) begin
      for (int z = 0 ; z < W ; z++) begin
        c[x][z] = state[x][0][z] ^ state[x][1][z]
                ^ state[x][2][z] ^ state[x][3][z] ^ state[x][4][z];
      end
    end
    for (int x = 0 ; x < 5 ; x++) begin
      int index_x1, index_x2;
      index_x1 = (x == 0) ? 4 : x-1; // (x-1)%5
      index_x2 = (x == 4) ? 0 : x+1; // (x+1)%5
      for (int z = 0 ; z < W ; z++) begin
        int index_z;
        index_z = (z == 0) ? W-1 : z-1; // (z+1)%W
        d[x][z] = c[index_x1][z] ^ c[index_x2][index_z];
      end
    end
    for (int x = 0 ; x < 5 ; x++) begin
      for (int y = 0 ; y < 5 ; y++) begin
        for (int z = 0 ; z < W ; z++) begin
          result[x][y][z] = state[x][y][z] ^ d[x][z];
        end
      end
    end
    return result;
  endfunction : theta

  // rho

  // Commented out entire rho function due to VCS elaboration error.
  // (z-RhoOffset[x][y]%W) isn't considered as a constant in VCS.
  // Even changing it to W-RhoOffset[x][y]%W and assign to ShiftAmt
  // creates same error.

  // Offset : Look at Table 2 in FIPS PUB 202
  //localparam int RhoOffset [5][5]  = '{
  //  //y  0    1    2    3    4     x
  //  '{   0,  36,   3, 105, 210},// 0
  //  '{   1, 300,  10,  45,  66},// 1
  //  '{ 190,   6, 171,  15, 253},// 2
  //  '{  28,  55, 153,  21, 120},// 3
  //  '{  91, 276, 231, 136,  78} // 4
  //};

  // rotate bits of each lane by offset
  // 1. rho[0,0,z] = A[0,0,z]
  // 2. Offset swap
  //    a. (x,y) := (1,0)
  //    b. for t [0..23]
  //       i. rho[x,y,z] = A[x,y,z-(t+1)(t+2)/2]
  //       ii. (x,y) = (y, (2x+3y))
  //function automatic box_t rho(box_t state);
  //  box_t result;
  //  for (int x = 0 ; x < 5 ; x++) begin
  //    for (int y = 0 ; y < 5 ; y++) begin
  //      for (int z = 0 ; z < W ; z++) begin
  //        automatic int index_z;
  //        index_z = (z-RhoOffset[x][y])%W;
  //        result[x][y][z] = state[x][y][(z-RhoOffset[x][y])%W];
  //      end
  //    end
  //  end
  //  return result;
  //endfunction : rho

  // pi
  // rearrange the position of lanes
  // pi[x,y,z] = state[(x+3y),x,z]
  localparam int PiRotate [5][5] = '{
    //y  0    1    2    3    4     x
    '{   0,   3,   1,   4,   2},// 0
    '{   1,   4,   2,   0,   3},// 1
    '{   2,   0,   3,   1,   4},// 2
    '{   3,   1,   4,   2,   0},// 3
    '{   4,   2,   0,   3,   1} // 4
  };
  function automatic box_t pi(box_t state);
    box_t result;
    for (int x = 0 ; x < 5 ; x++) begin
      for (int y = 0 ; y < 5 ; y++) begin
        int index_x;
        result[x][y][W-1:0] = state[PiRotate[x][y]][x][W-1:0];
      end
    end
    return result;
  endfunction : pi

  // chi
  // chi[x,y,z] = state[x,y,z] ^ ((state[x+1,y,z] ^ 1) & state[x+2,y,z])
  function automatic box_t chi(box_t state);
    box_t result;
    for (int x = 0 ; x < 5 ; x++) begin
      int index_x1, index_x2;
      index_x1 = (x == 4) ? 0 : x+1;
      index_x2 = (x >= 3) ? x-3 : x+2;
      for (int y = 0 ; y < 5 ; y++) begin
        for (int z = 0 ; z < W ; z++) begin
          result[x][y][z] = state[x][y][z] ^
                                ((~state[index_x1][y][z])
                                 & state[index_x2][y][z]);
        end
      end
    end
    return result;
  endfunction : chi

  // iota
  // XOR (x,y) = (0,0) with round constant

  // RC parameter: Precomputed by util/keccak_rc.py. Only up-to 0..L-1 is used
  // RC = '0
  // RC[2**j-1] = rc(j+7*rnd)
  // rc(t) =
  //    1. t%255 == 0 -> 1
  //    2. R[0:7] = 'b10000000
  //    3. for i = [1..t%255]
  //      a. R = 0 || R
  //      b. R[0] = R[0] ^ R[8]
  //      c. R[4] = R[4] ^ R[8]
  //      d. R[5] = R[5] ^ R[8]
  //      e. R[6] = R[6] ^ R[8]
  //      f. R = R[0:7]
  //    4. return R[0]
  // RC has L = [0..6]
  // for lower L case, only chopping lower part of 64bit RC is sufficient.
  localparam logic [63:0] RC [24] = '{
     64'h 0000_0000_0000_0001, // Round 0
     64'h 0000_0000_0000_8082, // Round 1
     64'h 8000_0000_0000_808A, // Round 2
     64'h 8000_0000_8000_8000, // Round 3
     64'h 0000_0000_0000_808B, // Round 4
     64'h 0000_0000_8000_0001, // Round 5
     64'h 8000_0000_8000_8081, // Round 6
     64'h 8000_0000_0000_8009, // Round 7
     64'h 0000_0000_0000_008A, // Round 8
     64'h 0000_0000_0000_0088, // Round 9
     64'h 0000_0000_8000_8009, // Round 10
     64'h 0000_0000_8000_000A, // Round 11
     64'h 0000_0000_8000_808B, // Round 12
     64'h 8000_0000_0000_008B, // Round 13
     64'h 8000_0000_0000_8089, // Round 14
     64'h 8000_0000_0000_8003, // Round 15
     64'h 8000_0000_0000_8002, // Round 16
     64'h 8000_0000_0000_0080, // Round 17
     64'h 0000_0000_0000_800A, // Round 18
     64'h 8000_0000_8000_000A, // Round 19
     64'h 8000_0000_8000_8081, // Round 20
     64'h 8000_0000_0000_8080, // Round 21
     64'h 0000_0000_8000_0001, // Round 22
     64'h 8000_0000_8000_8008  // Round 23
  };

  // iota: XOR with RC for (x,y) = (0,0)
  function automatic box_t iota(box_t state, logic [RndW-1:0] rnd);
    box_t result;
    result = state;
    result[0][0][W-1:0] = state[0][0][W-1:0] ^ RC[rnd][W-1:0];

    return result;
  endfunction : iota

  // Round function : Rnd(A,i_r)
  // Not used due to rho function issue described above.

  //function automatic box_t keccak_rnd(box_t state, logic [RndW-1:0] rnd);
  //  box_t keccak_state;
  //  keccak_state = iota(chi(pi(rho(theta(state)))), rnd);
  //
  //  return keccak_state;
  //endfunction : keccak_rnd

endmodule



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Combine InW data and write to OutW data if packed to full word or stop signal

`include "prim_assert.sv"

// ICEBOX(#12958): Revise to send out the empty status.
module prim_packer #(
  parameter int unsigned InW  = 32,
  parameter int unsigned OutW = 32,

  // If 1, The input/output are byte granularity
  parameter int HintByteData = 0,

  // Turn on protect against FI for the pos variable
  parameter bit EnProtection = 1'b 0
) (
  input clk_i ,
  input rst_ni,

  input                   valid_i,
  input        [InW-1:0]  data_i,
  input        [InW-1:0]  mask_i,
  output                  ready_o,

  output logic            valid_o,
  output logic [OutW-1:0] data_o,
  output logic [OutW-1:0] mask_o,
  input                   ready_i,

  input                   flush_i,  // If 1, send out remnant and clear state
  output logic            flush_done_o,

  // When EnProtection is set, err_o raises an error case (position variable
  // mismatch)
  output logic            err_o
);

  localparam int unsigned Width    = InW + OutW;  // storage width
  localparam int unsigned ConcatW  = Width + InW; // Input concatenated width
  localparam int unsigned PtrW     = $clog2(ConcatW+1);
  localparam int unsigned IdxW     = prim_util_pkg::vbits(InW);
  localparam int unsigned OnesCntW = $clog2(InW+1);

  logic valid_next, ready_next;
  logic [Width-1:0]   stored_data, stored_mask;
  logic [ConcatW-1:0] concat_data, concat_mask;
  logic [ConcatW-1:0] shiftl_data, shiftl_mask;
  logic [InW-1:0]     shiftr_data, shiftr_mask;

  logic [PtrW-1:0]     pos_q;         // Current write position
  logic [IdxW-1:0]     lod_idx;       // result of Leading One Detector
  logic [OnesCntW-1:0] inmask_ones;   // Counting Ones for mask_i

  logic ack_in, ack_out;

  logic flush_valid; // flush data out request
  logic flush_done;

  // Computing next position ==================================================
  always_comb begin
    // counting mask_i ones
    inmask_ones = '0;
    for (int i = 0 ; i < InW ; i++) begin
      inmask_ones = inmask_ones + OnesCntW'(mask_i[i]);
    end
  end

  logic [PtrW-1:0] pos_with_input;
  assign pos_with_input = pos_q + PtrW'(inmask_ones);

  if (EnProtection == 1'b 0) begin : g_pos_nodup
    logic [PtrW-1:0] pos_d;

    always_comb begin
      pos_d = pos_q;

      unique case ({ack_in, ack_out})
        2'b00: pos_d = pos_q;
        2'b01: pos_d = (int'(pos_q) <= OutW) ? '0 : pos_q - PtrW'(OutW);
        2'b10: pos_d = pos_with_input;
        2'b11: pos_d = (int'(pos_with_input) <= OutW) ? '0 : pos_with_input - PtrW'(OutW);
        default: pos_d = pos_q;
      endcase
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        pos_q <= '0;
      end else if (flush_done) begin
        pos_q <= '0;
      end else begin
        pos_q <= pos_d;
      end
    end

    assign err_o = 1'b 0; // No checker logic

  end else begin : g_pos_dupcnt // EnProtection == 1'b 1
    // incr_en: Increase the pos by cnt_step. ack_in && !ack_out
    // decr_en: Decrease the pos by cnt_step. !ack_in && ack_out
    // set_en:  Set to specific value in case of ack_in && ack_out.
    //          This case, the value could be increased or descreased based on
    //          the input size (inmask_ones)
    logic            cnt_incr_en, cnt_decr_en, cnt_set_en;
    logic [PtrW-1:0] cnt_step, cnt_set;

    assign cnt_incr_en =  ack_in && !ack_out;
    assign cnt_decr_en = !ack_in &&  ack_out;
    assign cnt_set_en  =  ack_in &&  ack_out;

    // counter has underflow protection.
    assign cnt_step = (cnt_incr_en) ? PtrW'(inmask_ones) : PtrW'(OutW);

    always_comb begin : cnt_set_logic

      // default, consuming all data
      cnt_set = '0;

      if (pos_with_input > PtrW'(OutW)) begin
        // pos_q + inmask_ones is bigger than Output width. Still data remained.
        cnt_set = pos_with_input - PtrW'(OutW);
      end
    end : cnt_set_logic


    prim_count #(
      .Width      (PtrW),
      .ResetValue ('0  )
    ) u_pos (
      .clk_i,
      .rst_ni,

      .clr_i      (flush_done),

      .set_i      (cnt_set_en),
      .set_cnt_i  (cnt_set   ),

      .incr_en_i  (cnt_incr_en),
      .decr_en_i  (cnt_decr_en),
      .step_i     (cnt_step   ),

      .cnt_o      (pos_q     ), // Current counter state
      .cnt_next_o (          ), // Next counter state

      .err_o
    );
  end // g_pos_dupcnt

  //---------------------------------------------------------------------------

  // Leading one detector for mask_i
  always_comb begin
    lod_idx = 0;
    for (int i = InW-1; i >= 0 ; i--) begin
      if (mask_i[i] == 1'b1) begin
        lod_idx = IdxW'(unsigned'(i));
      end
    end
  end

  assign ack_in  = valid_i & ready_o;
  assign ack_out = valid_o & ready_i;

  // Data process =============================================================
  //  shiftr : Input data shifted right to put the leading one at bit zero
  assign shiftr_data = (valid_i) ? data_i >> lod_idx : '0;
  assign shiftr_mask = (valid_i) ? mask_i >> lod_idx : '0;

  //  shiftl : Input data shifted into the current stored position
  assign shiftl_data = ConcatW'(shiftr_data) << pos_q;
  assign shiftl_mask = ConcatW'(shiftr_mask) << pos_q;

  // concat : Merging stored and shiftl
  assign concat_data = {{(InW){1'b0}}, stored_data & stored_mask} |
                       (shiftl_data & shiftl_mask);
  assign concat_mask = {{(InW){1'b0}}, stored_mask} | shiftl_mask;

  logic [Width-1:0] stored_data_next, stored_mask_next;

  always_comb begin
    unique case ({ack_in, ack_out})
      2'b 00: begin
        stored_data_next = stored_data;
        stored_mask_next = stored_mask;
      end
      2'b 01: begin
        // ack_out : shift the amount of OutW
        stored_data_next = {{OutW{1'b0}}, stored_data[Width-1:OutW]};
        stored_mask_next = {{OutW{1'b0}}, stored_mask[Width-1:OutW]};
      end
      2'b 10: begin
        // ack_in : Store concat data
        stored_data_next = concat_data[0+:Width];
        stored_mask_next = concat_mask[0+:Width];
      end
      2'b 11: begin
        // both : shift the concat_data
        stored_data_next = concat_data[ConcatW-1:OutW];
        stored_mask_next = concat_mask[ConcatW-1:OutW];
      end
      default: begin
        stored_data_next = stored_data;
        stored_mask_next = stored_mask;
      end
    endcase
  end

  // Store the data temporary if it doesn't exceed OutW
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      stored_data <= '0;
      stored_mask <= '0;
    end else if (flush_done) begin
      stored_data <= '0;
      stored_mask <= '0;
    end else begin
      stored_data <= stored_data_next;
      stored_mask <= stored_mask_next;
    end
  end
  //---------------------------------------------------------------------------

  // flush handling
  typedef enum logic {
    FlushIdle,
    FlushSend
  } flush_st_e;
  flush_st_e flush_st, flush_st_next;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      flush_st <= FlushIdle;
    end else begin
      flush_st <= flush_st_next;
    end
  end

  always_comb begin
    flush_st_next = FlushIdle;

    flush_valid = 1'b0;
    flush_done  = 1'b0;

    unique case (flush_st)
      FlushIdle: begin
        if (flush_i) begin
          flush_st_next = FlushSend;
        end else begin
          flush_st_next = FlushIdle;
        end
      end

      FlushSend: begin
        if (pos_q == '0) begin
          flush_st_next = FlushIdle;

          flush_valid = 1'b 0;
          flush_done  = 1'b 1;
        end else begin
          flush_st_next = FlushSend;

          flush_valid = 1'b 1;
          flush_done  = 1'b 0;
        end
      end
      default: begin
        flush_st_next = FlushIdle;

        flush_valid = 1'b 0;
        flush_done  = 1'b 0;
      end
    endcase
  end

  assign flush_done_o = flush_done;


  // Output signals ===========================================================
  assign valid_next = (int'(pos_q) >= OutW) ? 1'b 1 : flush_valid;

  // storage space is InW + OutW. So technically, ready_o can be asserted even
  // if `pos_q` is greater than OutW. But in order to do that, the logic should
  // use `inmask_ones` value whether pos_q+inmask_ones is less than (InW+OutW)
  // with `valid_i`. It creates a path from `valid_i` --> `ready_o`.
  // It may create a timing loop in some modules that use `ready_o` to
  // `valid_i` (which is not a good practice though)
  assign ready_next = int'(pos_q) <= OutW;

  // Output request
  assign valid_o = valid_next;
  assign data_o  = stored_data[OutW-1:0];
  assign mask_o  = stored_mask[OutW-1:0];

  // ready_o
  assign ready_o = ready_next;
  //---------------------------------------------------------------------------

  //////////////////////////////////////////////
  // Assertions, Assumptions, and Coverpoints //
  //////////////////////////////////////////////
  // Assumption: mask_i should be contiguous ones
  // e.g: 0011100 --> OK
  //      0100011 --> Not OK
  if (InW > 1) begin : gen_mask_assert
    `ASSUME(ContiguousOnesMask_M,
            valid_i |-> $countones(mask_i ^ {mask_i[InW-2:0],1'b0}) <= 2)
  end

  // Flush and Write Enable cannot be asserted same time
  `ASSUME(ExFlushValid_M, flush_i |-> !valid_i)

  // While in flush state, new request shouldn't come
  `ASSUME(ValidIDeassertedOnFlush_M,
          flush_st == FlushSend |-> $stable(valid_i))

  // If not acked, input port keeps asserting valid and data
  `ASSUME(DataIStable_M,
          ##1 valid_i && $past(valid_i) && !$past(ready_o)
          |-> $stable(data_i) && $stable(mask_i))

  `ASSERT(FlushFollowedByDone_A,
          ##1 $rose(flush_i) && !flush_done_o |-> !flush_done_o [*0:$] ##1 flush_done_o)

  // If not acked, valid_o should keep asserting
  `ASSERT(ValidOPairedWidthReadyI_A,
          valid_o && !ready_i |=> valid_o)

  // If stored data is greater than the output width, valid should be asserted
  `ASSERT(ValidOAssertedForStoredDataGTEOutW_A,
          ($countones(stored_mask) >= OutW) |-> valid_o)

  // If output port doesn't accept the data, the data should be stable
  `ASSERT(DataOStableWhenPending_A,
          ##1 valid_o && $past(valid_o)
          && !$past(ready_i) |-> $stable(data_o))

  // If input data & stored data are greater than OutW, remained should be stored
  `ASSERT(ExcessiveDataStored_A,
          ack_in && ack_out && (($countones(mask_i) + $countones(stored_mask)) > OutW)
          |=> (($past(data_i) &  $past(mask_i)) >>
               ($past(lod_idx)+OutW-$countones($past(stored_mask))))
               == stored_data)

  `ASSERT(ExcessiveMaskStored_A,
          ack_in && ack_out && (($countones(mask_i) + $countones(stored_mask)) > OutW)
          |=> ($past(mask_i) >>
               ($past(lod_idx)+OutW-$countones($past(stored_mask))))
              == stored_mask)

  // Assertions for byte hint enabled
  if (HintByteData != 0) begin : g_byte_assert
    `ASSERT_INIT(InputDividedBy8_A,  InW  % 8 == 0)
    `ASSERT_INIT(OutputDividedBy8_A, OutW % 8 == 0)

    // Masking[8*i+:8] should be all zero or all one
    for (genvar i = 0 ; i < InW/8 ; i++) begin : g_byte_input_masking
      `ASSERT(InputMaskContiguous_A,
              valid_i |-> (|mask_i[8*i+:8] == 1'b 0)
                       || (&mask_i[8*i+:8] == 1'b 1))
    end
    for (genvar i = 0 ; i < OutW/8 ; i++) begin : g_byte_output_masking
      `ASSERT(OutputMaskContiguous_A,
              valid_o |-> (|mask_o[8*i+:8] == 1'b 0)
                       || (&mask_o[8*i+:8] == 1'b 1))
    end
  end
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Supports packed and unpacked modes
// Uses FIFO timing on the control signals
// No masking or flush functions supported

// Timings - case where InW < OutW
// clk_i      __|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__
// wvalid_i   _____|~~~~|_____|~~~~|_____|~~~~|_____|~~~~|___________________
// wdata_i    Val N     |Val N+1   |Val N+2   |Val N+3   |-------------------
// wready_o   ~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~|__________|~~~~~~~~
// rvalid_o   ___________________________________________|~~~~~~~~~~|________
// rdata_o    -------------------------------------------|Val       |--------
// rready_i   _________________________________________________|~~~~|________
// depth_o    0000000000|1111111111|2222222222|3333333333|4444444444|00000000


// Timings - case where InW > OutW
// clk_i      __|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__
// wvalid_i   _____|~~~~|____________________________________________________
// wdata_i    -----|Val |----------------------------------------------------
// wready_o   ~~~~~~~~~~|___________________________________________|~~~~~~~~
// rvalid_o   __________|~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~|________
// rdata_o    ----------|Val N     |Val N+1   |Val N+2   |Val N+3   |--------
// rready_i   ________________|~~~~|_____|~~~~|_____|~~~~|_____|~~~~|________
// depth_o    0000000000|4444444444|3333333333|2222222222|1111111111|00000000


// Timings - case where InW = OutW
// clk_i      __|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__~~|__|~~|__
// wvalid_i   _____|~~~~|____________________________________________________
// wdata_i    -----|Val |----------------------------------------------------
// wready_o   ~~~~~~~~~~|__________|~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
// rvalid_o   __________|~~~~~~~~~~|_________________________________________
// rdata_o    ----------|Val       |-----------------------------------------
// rready_i   ________________|~~~~|_________________________________________
// depth_o    0000000000|1111111111|00000000000000000000000000000000000000000


`include "prim_assert.sv"

module prim_packer_fifo #(
  parameter int InW  = 32,
  parameter int OutW = 8,
  parameter bit ClearOnRead = 1'b1, // if == 1 always output 0 after read
  // derived parameters
  localparam int MaxW = (InW > OutW) ? InW : OutW,
  localparam int MinW = (InW < OutW) ? InW : OutW,
  localparam int DepthW = $clog2(MaxW/MinW)
) (
  input logic clk_i ,
  input logic rst_ni,

  input logic               clr_i,
  input logic               wvalid_i,
  input logic  [InW-1:0]    wdata_i,
  output logic              wready_o,

  output logic              rvalid_o,
  output logic [OutW-1:0]   rdata_o,
  input logic               rready_i,
  output logic [DepthW:0]   depth_o
);

  localparam int unsigned   WidthRatio = MaxW / MinW;
  localparam bit [DepthW:0] FullDepth = WidthRatio[DepthW:0];

  // signals
  logic  load_data;
  logic  clear_data;
  logic  clear_status;

  // flops
  logic [DepthW:0] depth_q, depth_d;
  logic [MaxW-1:0] data_q, data_d;
  logic            clr_q, clr_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      depth_q <= '0;
      data_q  <= '0;
      clr_q   <= 1'b1;
    end else begin
      depth_q <= depth_d;
      data_q  <= data_d;
      clr_q   <= clr_d;
    end
  end

  // flop for handling reset case for clr
  assign clr_d = clr_i;

  assign depth_o = depth_q;

  if (InW < OutW) begin : gen_pack_mode
    logic [MaxW-1:0] wdata_shifted;

    assign wdata_shifted = {{OutW - InW{1'b0}}, wdata_i} << (depth_q*InW);
    assign clear_status = (rready_i && rvalid_o) || clr_q;
    assign clear_data = (ClearOnRead && clear_status) || clr_q;
    assign load_data = wvalid_i && wready_o;

    assign depth_d =  clear_status ? '0 :
           load_data ? depth_q+1 :
           depth_q;

    assign data_d = clear_data ? '0 :
           load_data ? (wdata_shifted | (depth_q == 0 ? '0 : data_q)) :
           data_q;

    // set outputs
    assign wready_o = !(depth_q == FullDepth) && !clr_q;
    assign rdata_o =  data_q;
    assign rvalid_o = (depth_q == FullDepth) && !clr_q;

  end else begin : gen_unpack_mode
    logic [MaxW-1:0] rdata_shifted;
    logic            pull_data;
    logic [DepthW:0] ptr_q, ptr_d;
    logic [DepthW:0] lsb_is_one;
    logic [DepthW:0] max_value;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        ptr_q   <= '0;
      end else begin
        ptr_q   <= ptr_d;
      end
    end

    assign lsb_is_one = {{DepthW{1'b0}},1'b1};
    assign max_value = FullDepth;
    assign rdata_shifted = data_q >> ptr_q*OutW;
    assign clear_status = (rready_i && (depth_q == lsb_is_one)) || clr_q;
    assign clear_data = (ClearOnRead && clear_status) || clr_q;
    assign load_data = wvalid_i && wready_o;
    assign pull_data = rvalid_o && rready_i;

    assign depth_d =  clear_status ? '0 :
           load_data ? max_value :
           pull_data ? depth_q-1 :
           depth_q;

    assign ptr_d =  clear_status ? '0 :
           pull_data ? ptr_q+1 :
           ptr_q;

    assign data_d = clear_data ? '0 :
           load_data ? wdata_i :
           data_q;

    // set outputs
    assign wready_o = (depth_q == '0) && !clr_q;
    assign rdata_o =  rdata_shifted[OutW-1:0];
    assign rvalid_o = !(depth_q == '0) && !clr_q;

    // Avoid possible lint errors in case InW > OutW.
    if (InW > OutW) begin : gen_unused
      logic [MaxW-MinW-1:0] unused_rdata_shifted;
      assign unused_rdata_shifted = rdata_shifted[MaxW-1:MinW];
    end
  end


  //////////////////////////////////////////////
  // Assertions, Assumptions, and Coverpoints //
  //////////////////////////////////////////////

  // If not acked, valid_o should keep asserting
  `ASSERT(ValidOPairedWithReadyI_A,
          rvalid_o && !rready_i && !clr_i |=> rvalid_o)

  // If output port doesn't accept the data, the data should be stable
  `ASSERT(DataOStableWhenPending_A,
          ##1 rvalid_o && $past(rvalid_o)
          && !$past(rready_i) && !$past(clr_i) |-> $stable(rdata_o))

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Simple parameterizable gate generator. Used to fill up the netlist with gates that cannot be
// optimized away.
//
// The module leverages 4bit SBoxes from the PRINCE cipher, and interleaves them with registers,
// resulting in a split of around 50/50 between logic and sequential cells.
//
// This generator has been tested with 32bit wide data, and produces the following results:
//
// -------------+-----------+----------
// requested GE | actual GE | GE error
// -------------+-----------+----------
// 500          |  483      |  -17
// 1000         |  964      |  -36
// 1500         |  1447     |  -53
// 2500         |  2892     |  392
// 5000         |  5299     |  299
// 7500         |  8030     |  530
// 10000        |  10393    |  393
// 15000        |  15575    |  575
// 25000        |  26422    |  1422
// 50000        |  52859    |  2859
// 100000       |  105270   |  5270
//
// Note that the generator is not very accurate for smaller gate counts due to the generate loop
// granularity. Hence, do not use for fever than 500 GE.
//
// If valid_i constantly set to 1'b1, the gate generator produces around 2.5% smaller designs for
// the configurations listed in the table above.

`include "prim_assert.sv"
module prim_gate_gen #(
  parameter int DataWidth = 32,
  parameter int NumGates = 1000
) (
  input                        clk_i,
  input                        rst_ni,

  input                        valid_i,
  input        [DataWidth-1:0] data_i,
  output logic [DataWidth-1:0] data_o,
  output                       valid_o
);

  /////////////////////////////////////
  // Local parameters and assertions //
  /////////////////////////////////////

  // technology specific tuning, do not modify.
  // an inner round is comprised of a 2bit rotation, followed by a 4bit SBox Layer.
  localparam int NumInnerRounds = 2;
  localparam int GatesPerRound  = DataWidth * 14;
  // an outer round consists of NumInnerRounds, followed by a register.
  localparam int NumOuterRounds = (NumGates + GatesPerRound / 2) / GatesPerRound;

  // do not use for fewer than 500 GE
  `ASSERT(MinimumNumGates_A, NumGates >= 500)
  `ASSERT(DataMustBeMultipleOfFour_A, DataWidth % 4 == 0)

  /////////////////////
  // Generator Loops //
  /////////////////////

  logic [NumOuterRounds-1:0][DataWidth-1:0] regs_d, regs_q;
  logic [NumOuterRounds-1:0] valid_d, valid_q;

  for (genvar k = 0; k < NumOuterRounds; k++) begin : gen_outer_round

    logic [NumInnerRounds:0][DataWidth-1:0] inner_data;

    if (k==0) begin : gen_first
      assign inner_data[0] = data_i;
      assign valid_d[0]    = valid_i;
    end else begin : gen_others
      assign inner_data[0] = regs_q[k-1];
      assign valid_d[k]    = valid_q[k-1];
    end

    for (genvar l = 0; l < NumInnerRounds; l++) begin : gen_inner
      // 2bit rotation + sbox layer
      assign inner_data[l+1] = prim_cipher_pkg::sbox4_32bit({inner_data[l][1:0],
                                                             inner_data[l][DataWidth-1:2]},
                                                             prim_cipher_pkg::PRINCE_SBOX4);
    end

    assign regs_d[k] = inner_data[NumInnerRounds];
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : p_regs
    if (!rst_ni) begin
      regs_q <= '0;
      valid_q <= '0;
    end else begin
      valid_q <= valid_d;
      for (int k = 0; k < NumOuterRounds; k++) begin
        if (valid_d[k]) begin
          regs_q[k] <= regs_d[k];
        end
      end
    end
  end

  assign data_o = regs_q[NumOuterRounds-1];
  assign valid_o = valid_q[NumOuterRounds-1];

endmodule : prim_gate_gen


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Pulse synchronizer: synchronizes a pulse from source clock domain (clk_src)
// to destination clock domain (clk_dst). Each pulse has the length of one clock
// cycle of its respective clock domain. Consecutive pulses need to be spaced
// appropriately apart from each other depending on the clock frequency ratio
// of the two clock domains.

module prim_pulse_sync (
  // source clock domain
  input  logic clk_src_i,
  input  logic rst_src_ni,
  input  logic src_pulse_i,
  // destination clock domain
  input  logic clk_dst_i,
  input  logic rst_dst_ni,
  output logic dst_pulse_o
);

  ////////////////////////////////////////////////////////////////////////////////
  // convert src_pulse to a level signal so we can use double-flop synchronizer //
  ////////////////////////////////////////////////////////////////////////////////
  logic src_level;

  always_ff @(posedge clk_src_i or negedge rst_src_ni) begin
    if (!rst_src_ni) begin
      src_level <= 1'b0;
    end else begin
      src_level <= src_level ^ src_pulse_i;
    end
  end


  // source active must come far enough such that the destination domain has time
  // to create a valid pulse.
`ifdef INC_ASSERT
  //VCS coverage off
  // pragma coverage off

  // source active flag tracks whether there is an ongoing "toggle" event.
  // Until this toggle event is accepted by the destination domain (negative edge of
  // of the pulse output), the source side cannot toggle again.
  logic effective_rst_n;
  assign effective_rst_n = rst_src_ni && dst_pulse_o;

  logic src_active_flag_d, src_active_flag_q;
  assign src_active_flag_d = src_pulse_i || src_active_flag_q;

  always_ff @(posedge clk_src_i or negedge effective_rst_n) begin
    if (!effective_rst_n) begin
      src_active_flag_q <= '0;
    end else begin
      src_active_flag_q <= src_active_flag_d;
    end
  end

  //VCS coverage on
  // pragma coverage on

  `ASSERT(SrcPulseCheck_M, src_pulse_i |-> !src_active_flag_q, clk_src_i, !rst_src_ni)
`endif

  //////////////////////////////////////////////////////////
  // synchronize level signal to destination clock domain //
  //////////////////////////////////////////////////////////
  logic dst_level;

  prim_flop_2sync #(.Width(1)) prim_flop_2sync (
    // source clock domain
    .d_i    (src_level),
    // destination clock domain
    .clk_i  (clk_dst_i),
    .rst_ni (rst_dst_ni),
    .q_o    (dst_level)
  );

  ////////////////////////////////////////
  // convert level signal back to pulse //
  ////////////////////////////////////////
  logic dst_level_q;

  // delay dst_level by 1 cycle
  always_ff @(posedge clk_dst_i or negedge rst_dst_ni) begin
    if (!rst_dst_ni) begin
      dst_level_q <= 1'b0;
    end else begin
      dst_level_q <= dst_level;
    end
  end

  // edge detection
  assign dst_pulse_o = dst_level_q ^ dst_level;

  `ASSERT(DstPulseCheck_A, dst_pulse_o |=> !dst_pulse_o, clk_dst_i, !rst_dst_ni)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Primitive input filter, with enable.  Configurable number of cycles.
//
// when in reset, stored vector is zero
// when enable is false, output is input
// when enable is true, output is stored value,
//   new input must be opposite value from stored value for
//   #Cycles before switching to new value.

module prim_filter #(
  // If this parameter is set, an additional 2-stage synchronizer will be
  // added at the input.
  parameter bit AsyncOn = 0,
  parameter int unsigned Cycles = 4
) (
  input        clk_i,
  input        rst_ni,
  input        enable_i,
  input        filter_i,
  output logic filter_o
);

  logic [Cycles-1:0] stored_vector_q, stored_vector_d;
  logic stored_value_q, update_stored_value;
  logic unused_stored_vector_q_msb;

  logic filter_synced;

  if (AsyncOn) begin : gen_async
    // Run this through a 2 stage synchronizer to
    // prevent metastability.
    prim_flop_2sync #(
      .Width(1)
    ) prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(filter_i),
      .q_o(filter_synced)
    );
  end else begin : gen_sync
    assign filter_synced = filter_i;
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      stored_value_q <= 1'b0;
    end else if (update_stored_value) begin
      stored_value_q <= filter_synced;
    end
  end

  assign stored_vector_d = {stored_vector_q[Cycles-2:0],filter_synced};
  assign unused_stored_vector_q_msb = stored_vector_q[Cycles-1];

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      stored_vector_q <= '0;
    end else begin
      stored_vector_q <= stored_vector_d;
    end
  end

  assign update_stored_value =
             (stored_vector_d == {Cycles{1'b0}}) |
             (stored_vector_d == {Cycles{1'b1}});

  assign filter_o = enable_i ? stored_value_q : filter_synced;

endmodule



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Primitive counter-based input filter, with enable.
// Configurable number of cycles. Cheaper version of filter for
// large values of #Cycles
//
// when in reset, stored value is zero
// when enable is false, output is input
// when enable is true, output is stored value,
//   new input must be opposite value from stored value for
//   #Cycles before switching to new value.

module prim_filter_ctr #(
  // If this parameter is set, an additional 2-stage synchronizer will be
  // added at the input.
  parameter bit AsyncOn = 0,
  parameter int unsigned CntWidth = 2
) (
  input                clk_i,
  input                rst_ni,
  input                enable_i,
  input                filter_i,
  input [CntWidth-1:0] thresh_i,
  output logic         filter_o
);

  logic [CntWidth-1:0] diff_ctr_q, diff_ctr_d;
  logic filter_q, stored_value_q, update_stored_value;

  logic filter_synced;

  if (AsyncOn) begin : gen_async
    // Run this through a 2 stage synchronizer to
    // prevent metastability.
    prim_flop_2sync #(
      .Width(1)
    ) prim_flop_2sync (
      .clk_i,
      .rst_ni,
      .d_i(filter_i),
      .q_o(filter_synced)
    );
  end else begin : gen_sync
    assign filter_synced = filter_i;
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      filter_q <= 1'b0;
    end else begin
      filter_q <= filter_synced;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      stored_value_q <= 1'b0;
    end else if (update_stored_value) begin
      stored_value_q <= filter_synced;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      diff_ctr_q <= '0;
    end else begin
      diff_ctr_q <= diff_ctr_d;
    end
  end

  // always look for differences, even if not filter enabled
  assign update_stored_value = (diff_ctr_d == thresh_i);
  assign diff_ctr_d = (filter_synced != filter_q) ? '0       :           // restart
                      (diff_ctr_q >= thresh_i)    ? thresh_i :           // saturate
                                                    (diff_ctr_q + 1'b1); // count up

  assign filter_o = enable_i ? stored_value_q : filter_synced;

endmodule



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Primitive interrupt handler. This assumes the existence of three
// controller registers: INTR_ENABLE, INTR_STATE, INTR_TEST.
// This module can be instantiated once per interrupt field, or
// "bussified" with all fields of the interrupt vector.

module prim_intr_hw # (
  parameter int unsigned Width = 1,
  parameter bit FlopOutput = 1,

  // IntrT parameter is to hint the logic for the interrupt type. Module
  // supports two interrupt types, *Status* and *Event*.
  //
  // The differences between those two types are:
  // - Status is persistent. Until the root cause is alleviated, the interrupt
  //   keeps asserting.
  // - Event remains high for a relatively short period time without SW
  //   intervention. One distinct example is an error (error could be status
  //   though). If a certain error condition is captured, HW logic may create a
  //   pulse. In this case the interrupt is assumed as an Event interrupt.
  parameter IntrT = "Event" // Event or Status
) (
  // event
  input  clk_i,
  input  rst_ni,
  input  [Width-1:0]  event_intr_i,

  // register interface
  input  [Width-1:0]  reg2hw_intr_enable_q_i,
  input  [Width-1:0]  reg2hw_intr_test_q_i,
  input               reg2hw_intr_test_qe_i,
  input  [Width-1:0]  reg2hw_intr_state_q_i,
  output              hw2reg_intr_state_de_o,
  output [Width-1:0]  hw2reg_intr_state_d_o,

  // outgoing interrupt
  output logic [Width-1:0]  intr_o
);

  logic [Width-1:0] status; // incl. test

  if (IntrT == "Event") begin : g_intr_event
    logic  [Width-1:0]    new_event;
    assign new_event =
               (({Width{reg2hw_intr_test_qe_i}} & reg2hw_intr_test_q_i) | event_intr_i);
    assign hw2reg_intr_state_de_o = |new_event;
    // for scalar interrupts, this resolves to '1' with new event
    // for vector interrupts, new events are OR'd in to existing interrupt state
    assign hw2reg_intr_state_d_o  =  new_event | reg2hw_intr_state_q_i;

    assign status = reg2hw_intr_state_q_i ;
  end : g_intr_event
  else if (IntrT == "Status") begin : g_intr_status
    logic [Width-1:0] test_q; // Storing test. Cleared by SW

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) test_q <= '0;
      else if (reg2hw_intr_test_qe_i) test_q <= reg2hw_intr_test_q_i;
    end

    // TODO: In Status type, INTR_STATE is better to be external type and RO.
    assign hw2reg_intr_state_de_o = 1'b 1; // always represent the status
    assign hw2reg_intr_state_d_o  = event_intr_i | test_q;

    assign status = event_intr_i | test_q;

    // To make the timing same to event type, status signal does not use CSR.q,
    // rather the input of the CSR.
    logic unused_reg2hw;
    assign unused_reg2hw = ^reg2hw_intr_state_q_i;
  end : g_intr_status


  if (FlopOutput == 1) begin : gen_flop_intr_output
    // flop the interrupt output
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        intr_o <= '0;
      end else begin
        intr_o <= status & reg2hw_intr_enable_q_i;
      end
    end

  end else begin : gen_intr_passthrough_output
    logic unused_clk;
    logic unused_rst_n;
    assign unused_clk = clk_i;
    assign unused_rst_n = rst_ni;
    assign intr_o = reg2hw_intr_state_q_i & reg2hw_intr_enable_q_i;
  end

  `ASSERT_INIT(IntrTKind_A, IntrT inside {"Event", "Status"})

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// TL-UL fifo, used to add elasticity or an asynchronous clock crossing
// to an TL-UL bus.  This instantiates two FIFOs, one for the request side,
// and one for the response side.

module tlul_fifo_sync #(
  parameter bit          ReqPass = 1'b1,
  parameter bit          RspPass = 1'b1,
  parameter int unsigned ReqDepth = 2,
  parameter int unsigned RspDepth = 2,
  parameter int unsigned SpareReqW = 1,
  parameter int unsigned SpareRspW = 1
) (
  input                     clk_i,
  input                     rst_ni,
  input  tlul_pkg::tl_h2d_t tl_h_i,
  output tlul_pkg::tl_d2h_t tl_h_o,
  output tlul_pkg::tl_h2d_t tl_d_o,
  input  tlul_pkg::tl_d2h_t tl_d_i,
  input  [SpareReqW-1:0]    spare_req_i,
  output [SpareReqW-1:0]    spare_req_o,
  input  [SpareRspW-1:0]    spare_rsp_i,
  output [SpareRspW-1:0]    spare_rsp_o
);

  // Put everything on the request side into one FIFO
  localparam int unsigned REQFIFO_WIDTH = $bits(tlul_pkg::tl_h2d_t) -2 + SpareReqW;

  prim_fifo_sync #(.Width(REQFIFO_WIDTH), .Pass(ReqPass), .Depth(ReqDepth)) reqfifo (
    .clk_i,
    .rst_ni,
    .clr_i         (1'b0          ),
    .wvalid_i      (tl_h_i.a_valid),
    .wready_o      (tl_h_o.a_ready),
    .wdata_i       ({tl_h_i.a_opcode ,
                     tl_h_i.a_param  ,
                     tl_h_i.a_size   ,
                     tl_h_i.a_source ,
                     tl_h_i.a_address,
                     tl_h_i.a_mask   ,
                     tl_h_i.a_data   ,
                     tl_h_i.a_user   ,
                     spare_req_i}),
    .rvalid_o      (tl_d_o.a_valid),
    .rready_i      (tl_d_i.a_ready),
    .rdata_o       ({tl_d_o.a_opcode ,
                     tl_d_o.a_param  ,
                     tl_d_o.a_size   ,
                     tl_d_o.a_source ,
                     tl_d_o.a_address,
                     tl_d_o.a_mask   ,
                     tl_d_o.a_data   ,
                     tl_d_o.a_user   ,
                     spare_req_o}),
    .full_o        (),
    .depth_o       (),
    .err_o         ());

  // Put everything on the response side into the other FIFO

  localparam int unsigned RSPFIFO_WIDTH = $bits(tlul_pkg::tl_d2h_t) -2 + SpareRspW;

  prim_fifo_sync #(.Width(RSPFIFO_WIDTH), .Pass(RspPass), .Depth(RspDepth)) rspfifo (
    .clk_i,
    .rst_ni,
    .clr_i         (1'b0          ),
    .wvalid_i      (tl_d_i.d_valid),
    .wready_o      (tl_d_o.d_ready),
    .wdata_i       ({tl_d_i.d_opcode,
                     tl_d_i.d_param ,
                     tl_d_i.d_size  ,
                     tl_d_i.d_source,
                     tl_d_i.d_sink  ,
                     (tl_d_i.d_opcode == tlul_pkg::AccessAckData) ? tl_d_i.d_data :
                                                                    {top_pkg::TL_DW{1'b0}} ,
                     tl_d_i.d_user  ,
                     tl_d_i.d_error ,
                     spare_rsp_i}),
    .rvalid_o      (tl_h_o.d_valid),
    .rready_i      (tl_h_i.d_ready),
    .rdata_o       ({tl_h_o.d_opcode,
                     tl_h_o.d_param ,
                     tl_h_o.d_size  ,
                     tl_h_o.d_source,
                     tl_h_o.d_sink  ,
                     tl_h_o.d_data  ,
                     tl_h_o.d_user  ,
                     tl_h_o.d_error ,
                     spare_rsp_o}),
    .full_o        (),
    .depth_o       (),
    .err_o         ());

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// TL-UL fifo, used to add elasticity or an asynchronous clock crossing
// to an TL-UL bus.  This instantiates two FIFOs, one for the request side,
// and one for the response side.

`include "prim_assert.sv"

module tlul_fifo_async #(
  parameter int unsigned ReqDepth = 3,
  parameter int unsigned RspDepth = 3
) (
  input                      clk_h_i,
  input                      rst_h_ni,
  input                      clk_d_i,
  input                      rst_d_ni,
  input  tlul_pkg::tl_h2d_t  tl_h_i,
  output tlul_pkg::tl_d2h_t  tl_h_o,
  output tlul_pkg::tl_h2d_t  tl_d_o,
  input  tlul_pkg::tl_d2h_t  tl_d_i
);

  // Put everything on the request side into one FIFO
  localparam int unsigned REQFIFO_WIDTH = $bits(tlul_pkg::tl_h2d_t)-2;

  prim_fifo_async #(
    .Width(REQFIFO_WIDTH),
    .Depth(ReqDepth),
    .OutputZeroIfInvalid(1)
  ) reqfifo (
    .clk_wr_i      (clk_h_i),
    .rst_wr_ni     (rst_h_ni),
    .clk_rd_i      (clk_d_i),
    .rst_rd_ni     (rst_d_ni),
    .wvalid_i      (tl_h_i.a_valid),
    .wready_o      (tl_h_o.a_ready),
    .wdata_i       ({tl_h_i.a_opcode ,
                     tl_h_i.a_param  ,
                     tl_h_i.a_size   ,
                     tl_h_i.a_source ,
                     tl_h_i.a_address,
                     tl_h_i.a_mask   ,
                     tl_h_i.a_data   ,
                     tl_h_i.a_user   }),
    .rvalid_o      (tl_d_o.a_valid),
    .rready_i      (tl_d_i.a_ready),
    .rdata_o       ({tl_d_o.a_opcode ,
                     tl_d_o.a_param  ,
                     tl_d_o.a_size   ,
                     tl_d_o.a_source ,
                     tl_d_o.a_address,
                     tl_d_o.a_mask   ,
                     tl_d_o.a_data   ,
                     tl_d_o.a_user   }),
    .wdepth_o      (),
    .rdepth_o      ()
  );

  // Put everything on the response side into the other FIFO

  localparam int unsigned RSPFIFO_WIDTH = $bits(tlul_pkg::tl_d2h_t) -2;

  prim_fifo_async #(
    .Width(RSPFIFO_WIDTH),
    .Depth(RspDepth),
    .OutputZeroIfInvalid(1)
  ) rspfifo (
    .clk_wr_i      (clk_d_i),
    .rst_wr_ni     (rst_d_ni),
    .clk_rd_i      (clk_h_i),
    .rst_rd_ni     (rst_h_ni),
    .wvalid_i      (tl_d_i.d_valid),
    .wready_o      (tl_d_o.d_ready),
    .wdata_i       ({tl_d_i.d_opcode,
                     tl_d_i.d_param ,
                     tl_d_i.d_size  ,
                     tl_d_i.d_source,
                     tl_d_i.d_sink  ,
                     tl_d_i.d_data  ,
                     tl_d_i.d_user  ,
                     tl_d_i.d_error }),
    .rvalid_o      (tl_h_o.d_valid),
    .rready_i      (tl_h_i.d_ready),
    .rdata_o       ({tl_h_o.d_opcode,
                     tl_h_o.d_param ,
                     tl_h_o.d_size  ,
                     tl_h_o.d_source,
                     tl_h_o.d_sink  ,
                     tl_h_o.d_data  ,
                     tl_h_o.d_user  ,
                     tl_h_o.d_error }),
    .wdepth_o      (),
    .rdepth_o      ()
  );

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Protocol checker for TL-UL ports using assertions. Supports interface-widths
// up to 64bit.

`include "prim_assert.sv"

module tlul_assert #(
  parameter EndpointType = "Device" // can be either "Host" or "Device"
) (
  input clk_i,
  input rst_ni,

  // tile link ports
  input tlul_pkg::tl_h2d_t h2d,
  input tlul_pkg::tl_d2h_t d2h
);

`ifndef VERILATOR
`ifndef SYNTHESIS

`ifdef UVM
  import uvm_pkg::*;
`endif
  import tlul_pkg::*;
  import top_pkg::*;

  //////////////////////////////////
  // check requests and responses //
  //////////////////////////////////

  // There are up to 2**TL_AIW possible source-IDs. Below array "pend_req" has one entry
  // for each source-ID. Each entry has the following fields:
  //  - pend   : is set to 1 to indicate up to 1 pending request for the source ID
  //  - opcode : "Get" requires "AccessAckData" response, "Put*" require "AccessAck"
  //  - size   : d_size of response must match a_size of request
  //  - mask   : is used to allow X for bytes whose mask bit is 0
  typedef struct packed {
    bit                         pend; // set to 1 to indicate a pending request
    tl_a_op_e                   opcode;
    logic [top_pkg::TL_SZW-1:0] size;
    logic [top_pkg::TL_DBW-1:0] mask;
  } pend_req_t;

  pend_req_t [2**TL_AIW-1:0] pend_req;

  // set `disable_sva` before testing TLUL error cases
  bit disable_sva;
  // d_error related SVA doesn't work for xbar, as it doesn't return d_error for protocol errors
  // set this to disable the check
  bit disable_d_error_sva;

  logic [7:0]  a_mask, d_mask;
  logic [63:0] a_data, d_data;
  assign a_mask = 8'(h2d.a_mask);
  assign a_data = 64'(h2d.a_data);
  assign d_mask = 8'(pend_req[d2h.d_source].mask);
  assign d_data = 64'(d2h.d_data);

  ////////////////////////////////////
  // keep track of pending requests //
  ////////////////////////////////////

  // use negedge clk to avoid possible race conditions
  always_ff @(negedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      pend_req <= '0;
    end else begin
      if (h2d.a_valid) begin
        // store each request in pend_req array (we use blocking statements below so
        // that we can handle the case where request and response for the same
        // source-ID happen in the same cycle)
        if (d2h.a_ready) begin
          pend_req[h2d.a_source].pend    <= 1;
          pend_req[h2d.a_source].opcode  <= h2d.a_opcode;
          pend_req[h2d.a_source].size    <= h2d.a_size;
          pend_req[h2d.a_source].mask    <= h2d.a_mask;
        end
      end // h2d.a_valid

      if (d2h.d_valid) begin
        // update pend_req array
        if (h2d.d_ready) begin
          pend_req[d2h.d_source].pend <= 0;
        end
      end //d2h.d_valid
    end
  end

  /////////////////////////////////////////
  // define sequences for request checks //
  /////////////////////////////////////////

  sequence h2d_pre_S;
    h2d.a_valid;
  endsequence

  // a_opcode: only 3 opcodes are legal for requests
  sequence legalAOpcode_S;
    (h2d.a_opcode === PutFullData) ||
    (h2d.a_opcode === Get) ||
    (h2d.a_opcode === PutPartialData);
  endsequence

  // a_param is reserved
  sequence legalAParam_S;
    h2d.a_param === '0;
  endsequence

  // a_size: Size shouldn't be greater than the bus width in TL-UL (not in TL-UH)
  //         This assertion can be covered by below
  //         (a_size must less than or equal to ones of a_mask)

  // a_size: 2**a_size must greater than or equal to $countones(a_mask) for PutPartial and Get
  sequence sizeGTEMask_S;
    (h2d.a_opcode == PutFullData) || ((1 << h2d.a_size) >= $countones(h2d.a_mask));
  endsequence

  // a_size: 2**a_size must equal to $countones(a_mask) for PutFull
  sequence sizeMatchesMask_S;
    (h2d.a_opcode inside {PutPartialData, Get}) ||
    ((1 << h2d.a_size) === $countones(h2d.a_mask));
  endsequence

  // a_source: there should be no more than one pending request per each source ID
  sequence pendingReqPerSrc_S;
    pend_req[h2d.a_source].pend == 0;
  endsequence

  // a_address must be aligned to a_size: a_address & ((1 << a_size) - 1) == 0
  sequence addrSizeAligned_S;
    (h2d.a_address & ((1 << h2d.a_size)-1)) == '0;
  endsequence

  // a_mask must be contiguous for Get and PutFullData requests
  //    the spec talks about "naturally aligned". Does this mean that bit [0] of
  //    mask is always 1? If that's true, then below code could be much simpler.
  //    However, the spec shows a timing diagram where bit 0 of mask is 0.
  sequence contigMask_pre_S;
    h2d.a_opcode != PutPartialData;
  endsequence

  sequence contigMask_S;
    $countones(h2d.a_mask ^ {h2d.a_mask[$bits(h2d.a_mask)-2:0], 1'b0}) <= 2;
  endsequence

  // a_data must be known for opcode == Put*(depending on mask bits)
  sequence aDataKnown_pre_S;
    (h2d.a_opcode != Get);
  endsequence

  sequence aDataKnown_S;
    // no check if this lane mask is inactive
    ((!a_mask[0]) || (a_mask[0] && !$isunknown(a_data[8*0 +: 8]))) &&
    ((!a_mask[1]) || (a_mask[1] && !$isunknown(a_data[8*1 +: 8]))) &&
    ((!a_mask[2]) || (a_mask[2] && !$isunknown(a_data[8*2 +: 8]))) &&
    ((!a_mask[3]) || (a_mask[3] && !$isunknown(a_data[8*3 +: 8]))) &&
    ((!a_mask[4]) || (a_mask[4] && !$isunknown(a_data[8*4 +: 8]))) &&
    ((!a_mask[5]) || (a_mask[5] && !$isunknown(a_data[8*5 +: 8]))) &&
    ((!a_mask[6]) || (a_mask[6] && !$isunknown(a_data[8*6 +: 8]))) &&
    ((!a_mask[7]) || (a_mask[7] && !$isunknown(a_data[8*7 +: 8])));
  endsequence

  /////////////////////////////////////////
  // define sequences for request checks //
  /////////////////////////////////////////

  sequence d2h_pre_S;
    d2h.d_valid;
  endsequence

  // d_opcode: if request was Get, then response must be AccessAckData
  sequence respOpcode_S;
    d2h.d_opcode === ((pend_req[d2h.d_source].opcode == Get) ? AccessAckData : AccessAck);
  endsequence

  // d_param is reserved
  sequence legalDParam_S;
    d2h.d_param === '0;
  endsequence

  // d_size must equal the a_size of the corresponding request
  sequence respSzEqReqSz_S;
    d2h.d_size === pend_req[d2h.d_source].size;
  endsequence

  // d_source: each response should have a pending request using same source ID
  sequence respMustHaveReq_S;
    pend_req[d2h.d_source].pend;
  endsequence

// d_data must be known for AccessAckData (depending on mask bits)
  sequence dDataKnown_pre_S;
    d2h.d_opcode == AccessAckData;
  endsequence

  sequence dDataKnown_S;
    // no check if this lane mask is inactive
    ((!d_mask[0]) || (d_mask[0] && !$isunknown(d_data[8*0 +: 8]))) &&
    ((!d_mask[1]) || (d_mask[1] && !$isunknown(d_data[8*1 +: 8]))) &&
    ((!d_mask[2]) || (d_mask[2] && !$isunknown(d_data[8*2 +: 8]))) &&
    ((!d_mask[3]) || (d_mask[3] && !$isunknown(d_data[8*3 +: 8]))) &&
    ((!d_mask[4]) || (d_mask[4] && !$isunknown(d_data[8*4 +: 8]))) &&
    ((!d_mask[5]) || (d_mask[5] && !$isunknown(d_data[8*5 +: 8]))) &&
    ((!d_mask[6]) || (d_mask[6] && !$isunknown(d_data[8*6 +: 8]))) &&
    ((!d_mask[7]) || (d_mask[7] && !$isunknown(d_data[8*7 +: 8])));
  endsequence

  /////////////////////////////////////////
  // define sequences for d_error checks //
  /////////////////////////////////////////

  sequence d_error_pre_S;
    h2d.a_valid && d2h.a_ready;
  endsequence

  sequence legalAOpcodeErr_S;
    !(h2d.a_opcode inside {PutFullData, Get, PutPartialData});
  endsequence

  sequence sizeGTEMaskErr_S;
    (1 << h2d.a_size) < $countones(h2d.a_mask);
  endsequence

  sequence sizeMatchesMaskErr_S;
    (h2d.a_opcode == PutFullData) && ((1 << h2d.a_size) != $countones(h2d.a_mask));
  endsequence

  sequence addrSizeAlignedErr_S;
    (h2d.a_address & ((1 << h2d.a_size)-1)) != '0;
  endsequence

  ///////////////////////////////////
  // assemble properties and check //
  ///////////////////////////////////

  // note: use negedge clk to avoid possible race conditions
  // in this case all signals coming from the device side have an assumed property
  if (EndpointType == "Host") begin : gen_host
    // h2d
    `ASSERT(legalAOpcode_A,     h2d_pre_S |-> legalAOpcode_S,     !clk_i, !rst_ni || disable_sva)
    `ASSERT(legalAParam_A,      h2d_pre_S |-> legalAParam_S,      !clk_i, !rst_ni)
    `ASSERT(sizeGTEMask_A,      h2d_pre_S |-> sizeGTEMask_S,      !clk_i, !rst_ni || disable_sva)
    `ASSERT(sizeMatchesMask_A,  h2d_pre_S |-> sizeMatchesMask_S,  !clk_i, !rst_ni || disable_sva)
    `ASSERT(pendingReqPerSrc_A, h2d_pre_S |-> pendingReqPerSrc_S, !clk_i, !rst_ni)
    `ASSERT(addrSizeAligned_A,  h2d_pre_S |-> addrSizeAligned_S,  !clk_i, !rst_ni || disable_sva)
    `ASSERT(contigMask_A,       h2d_pre_S and contigMask_pre_S |-> contigMask_S,
          !clk_i, !rst_ni || disable_sva)
    `ASSERT(aDataKnown_A,       h2d_pre_S and aDataKnown_pre_S |-> aDataKnown_S, !clk_i, !rst_ni)
    // d2h
    `ASSUME(respOpcode_M,       d2h_pre_S |-> respOpcode_S,       !clk_i, !rst_ni)
    `ASSUME(legalDParam_M,      d2h_pre_S |-> legalDParam_S,      !clk_i, !rst_ni)
    `ASSUME(respSzEqReqSz_M,    d2h_pre_S |-> respSzEqReqSz_S,    !clk_i, !rst_ni)
    `ASSUME(respMustHaveReq_M,  d2h_pre_S |-> respMustHaveReq_S,  !clk_i, !rst_ni)
    `ASSUME(dDataKnown_M,       d2h_pre_S and dDataKnown_pre_S |-> dDataKnown_S,
          !clk_i, !rst_ni || disable_sva)
  // in this case all signals coming from the host side have an assumed property
  end else if (EndpointType == "Device") begin : gen_device
    // h2d
    `ASSUME(legalAParam_M,       h2d_pre_S |-> legalAParam_S,      !clk_i, !rst_ni)
    `ASSUME(pendingReqPerSrc_M,  h2d_pre_S |-> pendingReqPerSrc_S, !clk_i, !rst_ni)
    `ASSUME(aDataKnown_M,        h2d_pre_S and aDataKnown_pre_S |-> aDataKnown_S, !clk_i, !rst_ni)
    `ASSUME(contigMask_M,        h2d_pre_S and contigMask_pre_S |-> contigMask_S,
            !clk_i, !rst_ni || disable_sva)
    // d2h
    `ASSERT(respOpcode_A,        d2h_pre_S |-> respOpcode_S,       !clk_i, !rst_ni)
    `ASSERT(legalDParam_A,       d2h_pre_S |-> legalDParam_S,      !clk_i, !rst_ni)
    `ASSERT(respSzEqReqSz_A,     d2h_pre_S |-> respSzEqReqSz_S,    !clk_i, !rst_ni)
    `ASSERT(respMustHaveReq_A,   d2h_pre_S |-> respMustHaveReq_S,  !clk_i, !rst_ni)
    `ASSERT(dDataKnown_A,        d2h_pre_S and dDataKnown_pre_S |-> dDataKnown_S,
          !clk_i, !rst_ni || disable_sva)
    // d2h error cases
    `ASSERT(legalAOpcodeErr_A, d_error_pre_S and legalAOpcodeErr_S |=>
            s_eventually (d2h.d_valid && d2h.d_error), , !rst_ni || disable_d_error_sva)
    `ASSERT(sizeGTEMaskErr_A, d_error_pre_S and sizeGTEMaskErr_S |=>
            s_eventually (d2h.d_valid && d2h.d_error), , !rst_ni || disable_d_error_sva)
    `ASSERT(sizeMatchesMaskErr_A, d_error_pre_S and sizeMatchesMaskErr_S |=>
            s_eventually (d2h.d_valid && d2h.d_error), , !rst_ni || disable_d_error_sva)
    `ASSERT(addrSizeAlignedErr_A, d_error_pre_S and addrSizeAlignedErr_S |=>
            s_eventually (d2h.d_valid && d2h.d_error), , !rst_ni || disable_d_error_sva)
  end else begin : gen_unknown
    initial begin : p_unknonw
      `ASSERT_I(unknownConfig_A, 0 == 1)
    end
  end

  initial begin : p_dbw
    // widths up to 64bit / 8 Byte are supported
    `ASSERT_I(TlDbw_A, TL_DBW <= 8)
  end

  // make sure all "pending" bits are 0 at the end of the sim
  for (genvar ii = 0; ii < 2**TL_AIW; ii++) begin : gen_assert_final
    `ASSERT_FINAL(noOutstandingReqsAtEndOfSim_A, (pend_req[ii].pend == 0))
  end

  ////////////////////////////////////
  // additional checks for X values //
  ////////////////////////////////////

  // a_* should be known when a_valid == 1 (a_opcode and a_param are already covered above)
  // This also covers ASSERT_KNOWN of a_valid
  `ASSERT_KNOWN_IF(aKnown_A, {h2d.a_size, h2d.a_source, h2d.a_address, h2d.a_mask, h2d.a_user},
    h2d.a_valid)

  // d_* should be known when d_valid == 1 (d_opcode, d_param, d_size already covered above)
  // This also covers ASSERT_KNOWN of d_valid
  `ASSERT_KNOWN_IF(dKnown_A, {d2h.d_source, d2h.d_sink, d2h.d_error, d2h.d_user}, d2h.d_valid)

  //  make sure ready is not X after reset
  `ASSERT_KNOWN(aReadyKnown_A, d2h.a_ready)
  `ASSERT_KNOWN(dReadyKnown_A, h2d.d_ready)

  ////////////////////////////////////
  // SVA coverage //
  ////////////////////////////////////
  `define TLUL_COVER(SEQ) `COVER(``SEQ``_C, ``SEQ``_S, !clk_i, !rst_ni || disable_sva)

  // host sends back2back requests
  sequence b2bReq_S;
    h2d.a_valid && d2h.a_ready ##1 h2d.a_valid;
  endsequence

  // device sends back2back responses
  sequence b2bRsp_S;
    d2h.d_valid && h2d.d_ready ##1 d2h.d_valid;
  endsequence

  // host sends back2back requests with same address
  // UVM RAL can't issue this scenario, add this cover to make sure it's tested in some other seq
  sequence b2bReqWithSameAddr_S;
    bit [top_pkg::TL_AW-1:0] pre_addr;
    (h2d.a_valid && d2h.a_ready, pre_addr = h2d.a_address)
        ##1 h2d.a_valid && pre_addr == h2d.a_address;
  endsequence

  // a_valid is dropped without a_ready
  sequence aValidNotAccepted_S;
    h2d.a_valid && !d2h.a_ready ##1 !h2d.a_valid;
  endsequence

  // d_valid is dropped without a_ready
  sequence dValidNotAccepted_S;
    d2h.d_valid && !h2d.d_ready ##1 !d2h.d_valid;
  endsequence

  // host uses same source for back2back items
  sequence b2bSameSource_S;
    bit [top_pkg::TL_AIW-1:0] pre_source;
    (h2d.a_valid && d2h.a_ready, pre_source = h2d.a_source) ##1 h2d.a_valid[->1]
        ##0 pre_source == h2d.a_source;
  endsequence

  // a channal content is changed without being accepted
  `define TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(NAME) \
    sequence a_``NAME``ChangedNotAccepted_S; \
      int pre; \
      (h2d.a_valid && !d2h.a_ready, pre = h2d.a_``NAME``) ##1 h2d.a_valid[->1] \
          ##0 pre != h2d.a_``NAME``; \
    endsequence \
    `TLUL_COVER(a_``NAME``ChangedNotAccepted)

  // d channal content is changed without being accepted
  `define TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(NAME) \
    sequence d_``NAME``ChangedNotAccepted_S; \
      int pre; \
      (d2h.d_valid && !h2d.d_ready, pre = d2h.d_``NAME``) ##1 d2h.d_valid[->1] \
          ##0 pre != d2h.d_``NAME``; \
    endsequence \
    `TLUL_COVER(d_``NAME``ChangedNotAccepted)

  if (EndpointType == "Host") begin : gen_host_cov // DUT is host
    `TLUL_COVER(b2bRsp)
    `TLUL_COVER(dValidNotAccepted)
    `TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(data)
    `TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(opcode)
    `TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(size)
    `TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(source)
    `TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(sink)
    `TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED(error)
  end else if (EndpointType == "Device") begin : gen_device_cov // DUT is device
    `TLUL_COVER(b2bReq)
    `TLUL_COVER(b2bReqWithSameAddr)
    `TLUL_COVER(aValidNotAccepted)
    `TLUL_COVER(b2bSameSource)
    `TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(address)
    `TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(data)
    `TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(opcode)
    `TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(size)
    `TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(source)
    `TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED(mask)
  end else begin : gen_unknown_cov
    initial begin : p_unknonw_cov
      `ASSERT_I(unknownConfig_A, 0 == 1)
    end
  end

  `ifdef UVM
    initial forever begin
      bit tlul_assert_en;
      uvm_config_db#(bit)::wait_modified(null, "%m", "tlul_assert_en");
      if (!uvm_config_db#(bit)::get(null, "%m", "tlul_assert_en", tlul_assert_en)) begin
        `uvm_fatal("tlul_assert", "Can't find tlul_assert_en")
      end
      disable_sva = !tlul_assert_en;
    end
    initial forever begin
      bit tlul_assert_en;
      uvm_config_db#(bit)::wait_modified(null, "%m", "tlul_d_error_assert_en");
      if (!uvm_config_db#(bit)::get(null, "%m", "tlul_d_error_assert_en", tlul_assert_en)) begin
        `uvm_fatal("tlul_assert", "Can't find tlul_d_error_assert_en")
      end
      disable_d_error_sva = !tlul_assert_en;
    end
  `endif

  `undef TLUL_COVER
  `undef TLUL_A_CHAN_CONTENT_CHANGED_WO_ACCEPTED
  `undef TLUL_D_CHAN_CONTENT_CHANGED_WO_ACCEPTED
`endif
`endif
endmodule : tlul_assert


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0


`include "prim_assert.sv"

module tlul_err import tlul_pkg::*; (
  input clk_i,
  input rst_ni,

  input tl_h2d_t tl_i,

  output logic err_o
);

  localparam int IW  = $bits(tl_i.a_source);
  localparam int SZW = $bits(tl_i.a_size);
  localparam int DW  = $bits(tl_i.a_data);
  localparam int MW  = $bits(tl_i.a_mask);
  localparam int SubAW = $clog2(DW/8);

  logic opcode_allowed, a_config_allowed;

  logic op_full, op_partial, op_get;
  assign op_full    = (tl_i.a_opcode == PutFullData);
  assign op_partial = (tl_i.a_opcode == PutPartialData);
  assign op_get     = (tl_i.a_opcode == Get);

  // An instruction type transaction cannot be write
  logic instr_wr_err;
  assign instr_wr_err = prim_mubi_pkg::mubi4_test_true_strict(tl_i.a_user.instr_type) &
                        (op_full | op_partial);

  logic instr_type_err;
  assign instr_type_err = prim_mubi_pkg::mubi4_test_invalid(tl_i.a_user.instr_type);

  // Anything that doesn't fall into the permitted category, it raises an error
  assign err_o = ~(opcode_allowed & a_config_allowed) | instr_wr_err | instr_type_err;

  // opcode check
  assign opcode_allowed = (tl_i.a_opcode == PutFullData)
                        | (tl_i.a_opcode == PutPartialData)
                        | (tl_i.a_opcode == Get);

  // a channel configuration check
  logic addr_sz_chk;    // address and size alignment check
  logic mask_chk;       // inactive lane a_mask check
  logic fulldata_chk;   // PutFullData should have size match to mask

  logic [MW-1:0] mask;

  assign mask = (1 << tl_i.a_address[SubAW-1:0]);

  always_comb begin
    addr_sz_chk  = 1'b0;
    mask_chk     = 1'b0;
    fulldata_chk = 1'b0; // Only valid when opcode is PutFullData

    if (tl_i.a_valid) begin
      unique case (tl_i.a_size)
        'h0: begin // 1 Byte
          addr_sz_chk  = 1'b1;
          mask_chk     = ~|(tl_i.a_mask & ~mask);
          fulldata_chk = |(tl_i.a_mask & mask);
        end

        'h1: begin // 2 Byte
          addr_sz_chk  = ~tl_i.a_address[0];
          // check inactive lanes if lower 2B, check a_mask[3:2], if uppwer 2B, a_mask[1:0]
          mask_chk     = (tl_i.a_address[1]) ? ~|(tl_i.a_mask & 4'b0011)
                       : ~|(tl_i.a_mask & 4'b1100);
          fulldata_chk = (tl_i.a_address[1]) ? &tl_i.a_mask[3:2] : &tl_i.a_mask[1:0] ;
        end

        'h2: begin // 4 Byte
          addr_sz_chk  = ~|tl_i.a_address[SubAW-1:0];
          mask_chk     = 1'b1;
          fulldata_chk = &tl_i.a_mask[3:0];
        end

        default: begin // else
          addr_sz_chk  = 1'b0;
          mask_chk     = 1'b0;
          fulldata_chk = 1'b0;
        end
      endcase
    end else begin
      addr_sz_chk  = 1'b0;
      mask_chk     = 1'b0;
      fulldata_chk = 1'b0;
    end
  end

  assign a_config_allowed = addr_sz_chk
                          & mask_chk
                          & (op_get | op_partial | fulldata_chk) ;

  // Only 32 bit data width for current tlul_err
  `ASSERT_INIT(dataWidthOnly32_A, DW == 32)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0


`include "prim_assert.sv"

module tlul_err64 import tlul_pkg::*; (
  input clk_i,
  input rst_ni,

  input tl_h2d_t64 tl_i,

  output logic err_o
);

  localparam int IW  = $bits(tl_i.a_source);
  localparam int SZW = $bits(tl_i.a_size);
  localparam int DW  = $bits(tl_i.a_data);
  localparam int MW  = $bits(tl_i.a_mask);
  localparam int SubAW = $clog2(DW/8);

  logic opcode_allowed, a_config_allowed;

  logic op_full, op_partial, op_get;
  assign op_full    = (tl_i.a_opcode == PutFullData);
  assign op_partial = (tl_i.a_opcode == PutPartialData);
  assign op_get     = (tl_i.a_opcode == Get);

  // An instruction type transaction cannot be write
  logic instr_wr_err;
  assign instr_wr_err = prim_mubi_pkg::mubi4_test_true_strict(tl_i.a_user.instr_type) &
                        (op_full | op_partial);

  logic instr_type_err;
  assign instr_type_err = prim_mubi_pkg::mubi4_test_invalid(tl_i.a_user.instr_type);

  // Anything that doesn't fall into the permitted category, it raises an error
  assign err_o = ~(opcode_allowed & a_config_allowed) | instr_wr_err | instr_type_err;

  // opcode check
  assign opcode_allowed = (tl_i.a_opcode == PutFullData)
                        | (tl_i.a_opcode == PutPartialData)
                        | (tl_i.a_opcode == Get);

  // a channel configuration check
  logic addr_sz_chk;    // address and size alignment check
  logic mask_chk;       // inactive lane a_mask check
  logic fulldata_chk;   // PutFullData should have size match to mask

  logic [MW-1:0] mask;

  assign mask = (1 << tl_i.a_address[SubAW-1:0]);

  always_comb begin
    addr_sz_chk  = 1'b0;
    mask_chk     = 1'b0;
    fulldata_chk = 1'b0; // Only valid when opcode is PutFullData

    if (tl_i.a_valid) begin
      unique case (tl_i.a_size)
        'h0: begin // 1 Byte
          addr_sz_chk  = 1'b1;
          mask_chk     = ~|(tl_i.a_mask & ~mask);
          fulldata_chk = |(tl_i.a_mask & mask);
        end

        'h1: begin // 2 Byte
          addr_sz_chk  = ~tl_i.a_address[0];
          // check inactive lanes if lower 2B, check a_mask[3:2], if uppwer 2B, a_mask[1:0]
          mask_chk     = (tl_i.a_address[1]) ? ~|(tl_i.a_mask & 4'b0011)
                       : ~|(tl_i.a_mask & 4'b1100);
          fulldata_chk = (tl_i.a_address[1]) ? &tl_i.a_mask[3:2] : &tl_i.a_mask[1:0] ;
        end

        'h2: begin // 4 Byte
          addr_sz_chk  = ~|tl_i.a_address[SubAW-1:0];
          mask_chk     = 1'b1;
          fulldata_chk = &tl_i.a_mask[3:0];
        end

        default: begin // else
          addr_sz_chk  = 1'b0;
          mask_chk     = 1'b0;
          fulldata_chk = 1'b0;
        end
      endcase
    end else begin
      addr_sz_chk  = 1'b0;
      mask_chk     = 1'b0;
      fulldata_chk = 1'b0;
    end
  end

  assign a_config_allowed = addr_sz_chk
                          & mask_chk
                          & (op_get | op_partial | fulldata_chk) ;

  // Only 32 bit data width for current tlul_err
  `ASSERT_INIT(dataWidthOnly32_A, DW == 32)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

// Protocol checker for multiple TL-UL ports

module tlul_assert_multiple #(
  parameter int unsigned N = 2,
  parameter EndpointType = "Device" // can be "Device" or "Host"
) (
  input clk_i,
  input rst_ni,

  // tile link ports
  input tlul_pkg::tl_h2d_t h2d [N],
  input tlul_pkg::tl_d2h_t d2h [N]
);

  // instantiate N tlul_assert modules
  for (genvar ii = 0; ii < N; ii++) begin : gen_assert
    tlul_assert #(
      .EndpointType(EndpointType)
    ) tlul_assert (
      .clk_i,
      .rst_ni,
      // TL-UL ports
      .h2d (h2d[ii]),
      .d2h (d2h[ii])
    );
  end
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Flash Controller module.
//

package flash_ctrl_pkg;

  // design parameters that can be altered through topgen
  parameter int unsigned NumBanks        = flash_ctrl_reg_pkg::RegNumBanks;
  parameter int unsigned PagesPerBank    = flash_ctrl_reg_pkg::RegPagesPerBank;
  parameter int unsigned BusPgmResBytes  = flash_ctrl_reg_pkg::RegBusPgmResBytes;
  // How many types of info per bank
  parameter int InfoTypes                = flash_ctrl_reg_pkg::NumInfoTypes;

  // fixed parameters of flash derived from topgen parameters
  parameter int DataWidth       = 64;
  parameter int MetaDataWidth   = 12;

// The following hard-wired values are there to work-around verilator.
// For some reason if the values are assigned through parameters verilator thinks
// they are not constant
  parameter int InfoTypeSize [InfoTypes] = '{
    10,
    1,
    2
  };
  parameter int InfosPerBank    = max_info_pages('{
    10,
    1,
    2
  });
  parameter int WordsPerPage    = 256; // Number of flash words per page
  parameter int BusWidth        = top_pkg::TL_DW;
  parameter int BusIntgWidth    = tlul_pkg::DataIntgWidth;
  parameter int BusFullWidth    = BusWidth + BusIntgWidth;
  parameter int MpRegions       = 8;  // flash controller protection regions
  //parameter int FifoDepth       = 16; // rd / prog fifos
  parameter int InfoTypesWidth  = prim_util_pkg::vbits(InfoTypes);

  // flash phy parameters
  parameter int DataByteWidth   = prim_util_pkg::vbits(DataWidth / 8);
  parameter int BankW           = prim_util_pkg::vbits(NumBanks);
  parameter int InfoPageW       = prim_util_pkg::vbits(InfosPerBank);
  parameter int PageW           = prim_util_pkg::vbits(PagesPerBank);
  parameter int WordW           = prim_util_pkg::vbits(WordsPerPage);
  parameter int AddrW           = BankW + PageW + WordW; // all flash range
  parameter int BankAddrW       = PageW + WordW;         // 1 bank of flash range
  parameter int AllPagesW       = BankW + PageW;

  // flash ctrl / bus parameters
  // flash / bus width may be different from actual flash word width
  parameter int BusBytes        = BusWidth / 8;
  parameter int BusByteWidth    = prim_util_pkg::vbits(BusBytes);
  parameter int WidthMultiple   = DataWidth / BusWidth;
  // Number of bus words that can be programmed at once
  parameter int BusPgmRes       = BusPgmResBytes / BusBytes;
  parameter int BusPgmResWidth  = prim_util_pkg::vbits(BusPgmRes);
  parameter int BusWordsPerPage = WordsPerPage * WidthMultiple;
  parameter int BusWordW        = prim_util_pkg::vbits(BusWordsPerPage);
  parameter int BusAddrW        = BankW + PageW + BusWordW;
  parameter int BusAddrByteW    = BusAddrW + BusByteWidth;
  parameter int BusBankAddrW    = PageW + BusWordW;
  parameter int PhyAddrStart    = BusWordW - WordW;

  // fifo parameters
  //parameter int FifoDepthW      = prim_util_pkg::vbits(FifoDepth+1);

  // The end address in bus words for each kind of partition in each bank
  parameter logic [PageW-1:0] DataPartitionEndAddr = PageW'(PagesPerBank - 1);
  //parameter logic [PageW-1:0] InfoPartitionEndAddr [InfoTypes] = '{
  //  9,
  //  0,
  //  1
  //};
  parameter logic [PageW-1:0] InfoPartitionEndAddr [InfoTypes] = '{
    PageW'(InfoTypeSize[0] - 1),
    PageW'(InfoTypeSize[1] - 1),
    PageW'(InfoTypeSize[2] - 1)
  };

  // Flash Disable usage
  typedef enum logic [3:0] {
    PhyDisableIdx,
    ArbFsmDisableIdx,
    LcMgrDisableIdx,
    MpDisableIdx,
    HostDisableIdx,
    IFetchDisableIdx,
    RdFifoIdx,
    ProgFifoIdx,
    FlashDisableLast
  } flash_disable_pos_e;

  ////////////////////////////
  // All memory protection, seed related parameters
  // Those related for seed pages should be template candidates
  ////////////////////////////

  // parameters for connected components
  parameter int SeedWidth = 256;
  parameter int KeyWidth  = 128;
  parameter int EdnWidth  = edn_pkg::ENDPOINT_BUS_WIDTH;
  typedef logic [KeyWidth-1:0] flash_key_t;

  // Default Lfsr configurations
  // These LFSR parameters have been generated with
  // $ util/design/gen-lfsr-seed.py --width 32 --seed 1274809145 --prefix ""
  parameter int LfsrWidth = 32;
  typedef logic [LfsrWidth-1:0] lfsr_seed_t;
  typedef logic [LfsrWidth-1:0][$clog2(LfsrWidth)-1:0] lfsr_perm_t;
  parameter lfsr_seed_t RndCnstLfsrSeedDefault = 32'ha8cee782;
  parameter lfsr_perm_t RndCnstLfsrPermDefault = {
    160'hd60bc7d86445da9347e0ccdd05b281df95238bb5
  };

  // These LFSR parameters have been generated with
  // $ util/design/gen-lfsr-seed.py --width 64 --seed 691876113 --prefix ""


  // lcmgr phase enum
  typedef enum logic [1:0] {
    PhaseSeed,
    PhaseRma,
    PhaseNone,
    PhaseInvalid
  } flash_lcmgr_phase_e;

  import flash_ctrl_reg_pkg::flash_ctrl_reg2hw_mp_bank_cfg_shadowed_mreg_t;
  import flash_ctrl_reg_pkg::flash_ctrl_reg2hw_mp_region_mreg_t;
  import flash_ctrl_reg_pkg::flash_ctrl_reg2hw_mp_region_cfg_mreg_t;
  import flash_ctrl_reg_pkg::flash_ctrl_reg2hw_bank0_info0_page_cfg_mreg_t;
  import flash_ctrl_reg_pkg::flash_ctrl_reg2hw_default_region_reg_t;

  typedef flash_ctrl_reg2hw_mp_bank_cfg_shadowed_mreg_t sw_bank_cfg_t;
  typedef flash_ctrl_reg2hw_mp_region_mreg_t sw_region_t;
  typedef flash_ctrl_reg2hw_mp_region_cfg_mreg_t sw_region_cfg_t;
  typedef flash_ctrl_reg2hw_default_region_reg_t sw_default_cfg_t;
  typedef flash_ctrl_reg2hw_bank0_info0_page_cfg_mreg_t sw_info_cfg_t;

  // alias for super long reg_pkg typedef
  typedef struct packed {
    logic        q;
  } bank_cfg_t;

  import prim_mubi_pkg::mubi4_t;
  import prim_mubi_pkg::MuBi4True;
  import prim_mubi_pkg::MuBi4False;

  // This is identical to the reg structures but do not have err_updates / storage
  typedef struct packed {
    mubi4_t en;
    mubi4_t rd_en;
    mubi4_t prog_en;
    mubi4_t erase_en;
    mubi4_t scramble_en;
    mubi4_t ecc_en;
    mubi4_t he_en;
  } info_page_cfg_t;

  // This is identical to the reg structures but do not have err_updates / storage
  typedef struct packed {
    mubi4_t en;
    mubi4_t rd_en;
    mubi4_t prog_en;
    mubi4_t erase_en;
    mubi4_t scramble_en;
    mubi4_t ecc_en;
    mubi4_t he_en;
    logic [8:0] base;
    logic [9:0] size;
  } mp_region_cfg_t;

  // memory protection specific structs
  typedef struct packed {
    logic [InfoTypesWidth-1:0] sel;
    logic [AllPagesW-1:0] addr;
  } page_addr_t;

  typedef struct packed {
    page_addr_t           page;
    flash_lcmgr_phase_e   phase;
    info_page_cfg_t       cfg;
  } info_page_attr_t;

  typedef struct packed {
    flash_lcmgr_phase_e   phase;
    mp_region_cfg_t cfg;
  } data_region_attr_t;

  // flash life cycle / key manager management constants
  // One page for creator seeds
  // One page for owner seeds
  // One page for isolated flash page
  parameter int NumSeeds = 2;
  parameter bit [BankW-1:0] SeedBank = 0;
  parameter bit [InfoTypesWidth-1:0] SeedInfoSel = 0;
  parameter bit [0:0] CreatorSeedIdx = 0;
  parameter bit [0:0] OwnerSeedIdx = 1;
  parameter bit [PageW-1:0] CreatorInfoPage = 1;
  parameter bit [PageW-1:0] OwnerInfoPage = 2;
  parameter bit [PageW-1:0] IsolatedInfoPage = 3;

  parameter int TotalSeedWidth = SeedWidth * NumSeeds;
  typedef logic [TotalSeedWidth-1:0] all_seeds_t;

  // which page of which info type of which bank for seed selection
  parameter page_addr_t SeedInfoPageSel [NumSeeds] = '{
    '{
      sel:  SeedInfoSel,
      addr: {SeedBank, CreatorInfoPage}
     },

    '{
      sel:  SeedInfoSel,
      addr: {SeedBank, OwnerInfoPage}
     }
  };

  // which page of which info type of which bank for isolated partition
  parameter page_addr_t IsolatedPageSel = '{
    sel:  SeedInfoSel,
    addr: {SeedBank, IsolatedInfoPage}
  };

  // hardware interface memory protection rules
  parameter int HwInfoRules = 5;
  parameter int HwDataRules = 1;

  parameter info_page_cfg_t CfgAllowRead = '{
    en:          MuBi4True,
    rd_en:       MuBi4True,
    prog_en:     MuBi4False,
    erase_en:    MuBi4False,
    scramble_en: MuBi4True,
    ecc_en:      MuBi4True,
    he_en:       MuBi4True
  };

  parameter info_page_cfg_t CfgAllowReadProgErase = '{
    en:          MuBi4True,
    rd_en:       MuBi4True,
    prog_en:     MuBi4True,
    erase_en:    MuBi4True,
    scramble_en: MuBi4True,
    ecc_en:      MuBi4True,
    he_en:       MuBi4True   // HW assumes high endurance
  };

  parameter info_page_cfg_t CfgInfoDisable = '{
    en:          MuBi4False,
    rd_en:       MuBi4False,
    prog_en:     MuBi4False,
    erase_en:    MuBi4False,
    scramble_en: MuBi4False,
    ecc_en:      MuBi4False,
    he_en:       MuBi4False
  };

  parameter info_page_attr_t HwInfoPageAttr[HwInfoRules] = '{
    '{
       page:  SeedInfoPageSel[CreatorSeedIdx],
       phase: PhaseSeed,
       cfg:   CfgAllowRead
     },

    '{
       page:  SeedInfoPageSel[OwnerSeedIdx],
       phase: PhaseSeed,
       cfg:   CfgAllowRead
     },

    '{
       page:  SeedInfoPageSel[CreatorSeedIdx],
       phase: PhaseRma,
       cfg:   CfgAllowReadProgErase
     },

    '{
       page:  SeedInfoPageSel[OwnerSeedIdx],
       phase: PhaseRma,
       cfg:   CfgAllowReadProgErase
     },

    '{
       page:  IsolatedPageSel,
       phase: PhaseRma,
       cfg:   CfgAllowReadProgErase
     }
  };

  parameter data_region_attr_t HwDataAttr[HwDataRules] = '{
    '{
       phase: PhaseRma,
       cfg:   '{
                 en:          MuBi4True,
                 rd_en:       MuBi4True,
                 prog_en:     MuBi4True,
                 erase_en:    MuBi4True,
                 scramble_en: MuBi4True,
                 ecc_en:      MuBi4True,
                 he_en:       MuBi4True, // HW assumes high endurance
                 base:        '0,
                 size:        NumBanks * PagesPerBank
                }
     }
  };


  ////////////////////////////
  // Design time constants
  ////////////////////////////
  parameter flash_key_t RndCnstAddrKeyDefault =
    128'h5d707f8a2d01d400928fa691c6a6e0a4;
  parameter flash_key_t RndCnstDataKeyDefault =
    128'h39953618f2ca6f674af39f64975ea1f5;
  parameter all_seeds_t RndCnstAllSeedsDefault = {
    256'h3528874c0d9e481ead4d240eb6238a2c6218896f5315edb5ccefe029a6d04091,
    256'h9cde77e25a313a76984ab0ebf990983432b03b48186dcd556565fe721b447477
  };


  ////////////////////////////
  // Flash operation related enums
  ////////////////////////////

  // Flash Operations Supported
  typedef enum logic [1:0] {
    FlashOpRead     = 2'h0,
    FlashOpProgram  = 2'h1,
    FlashOpErase    = 2'h2,
    FlashOpInvalid  = 2'h3
  } flash_op_e;

  // Flash Program Operations Supported
  typedef enum logic {
    FlashProgNormal = 0,
    FlashProgRepair = 1
  } flash_prog_e;
  parameter int ProgTypes = 2;

  // Flash Erase Operations Supported
  typedef enum logic  {
    FlashErasePage  = 0,
    FlashEraseBank  = 1
  } flash_erase_e;

  // Flash function select
  typedef enum logic [1:0] {
    NoneSel,
    SwSel,
    HwSel
  } flash_sel_e;

  // Flash tlul to fifo direction
  typedef enum logic  {
    WriteDir     = 1'b0,
    ReadDir      = 1'b1
  } flash_flfo_dir_e;

  // Flash partition type
  typedef enum logic {
    FlashPartData = 1'b0,
    FlashPartInfo = 1'b1
  } flash_part_e;

  // Flash controller to memory
  typedef struct packed {
    logic                 req;
    logic                 scramble_en;
    logic                 ecc_en;
    logic                 he_en;
    logic                 rd_buf_en;
    logic                 rd;
    logic                 prog;
    logic                 pg_erase;
    logic                 bk_erase;
    logic                 erase_suspend;
    flash_part_e          part;
    logic [InfoTypesWidth-1:0] info_sel;
    logic [BusAddrW-1:0]  addr;
    logic [BusFullWidth-1:0] prog_data;
    logic                 prog_last;
    flash_prog_e          prog_type;
    mp_region_cfg_t [MpRegions:0] region_cfgs;
    logic [KeyWidth-1:0]  addr_key;
    logic [KeyWidth-1:0]  data_key;
    logic [KeyWidth-1:0]  rand_addr_key;
    logic [KeyWidth-1:0]  rand_data_key;
    logic                 alert_trig;
    logic                 alert_ack;
    jtag_pkg::jtag_req_t  jtag_req;
    prim_mubi_pkg::mubi4_t flash_disable;
  } flash_req_t;

  // default value of flash_req_t (for dangling ports)
  parameter flash_req_t FLASH_REQ_DEFAULT = '{
    req:           '0,
    scramble_en:   '0,
    ecc_en:        '0,
    he_en:         '0,
    rd_buf_en:     1'b0,
    rd:            '0,
    prog:          '0,
    pg_erase:      '0,
    bk_erase:      '0,
    erase_suspend: '0,
    part:          FlashPartData,
    info_sel:      '0,
    addr:          '0,
    prog_data:     '0,
    prog_last:     '0,
    prog_type:     FlashProgNormal,
    region_cfgs:   '0,
    addr_key:      RndCnstAddrKeyDefault,
    data_key:      RndCnstDataKeyDefault,
    rand_addr_key: '0,
    rand_data_key: '0,
    alert_trig:    1'b0,
    alert_ack:     1'b0,
    jtag_req:      '0,
    flash_disable: prim_mubi_pkg::MuBi4False
  };

  // memory to flash controller
  typedef struct packed {
    logic [ProgTypes-1:0]    prog_type_avail;
    logic                    rd_done;
    logic                    prog_done;
    logic                    erase_done;
    logic                    rd_err;
    logic [BusFullWidth-1:0] rd_data;
    logic                    init_busy;
    logic                    macro_err;
    logic [NumBanks-1:0]     ecc_single_err;
    logic [NumBanks-1:0][BusAddrW-1:0] ecc_addr;
    jtag_pkg::jtag_rsp_t     jtag_rsp;
    logic                    prog_intg_err;
    logic                    storage_relbl_err;
    logic                    storage_intg_err;
    logic                    fsm_err;
    logic                    spurious_ack;
    logic                    arb_err;
    logic                    host_gnt_err;
    logic                    fifo_err;
  } flash_rsp_t;

  // default value of flash_rsp_t (for dangling ports)
  parameter flash_rsp_t FLASH_RSP_DEFAULT = '{
    prog_type_avail:    {ProgTypes{1'b1}},
    rd_done:            1'b0,
    prog_done:          1'b0,
    erase_done:         1'b0,
    rd_err:             '0,
    rd_data:            '0,
    init_busy:          1'b0,
    macro_err:          1'b0,
    ecc_single_err:     '0,
    ecc_addr:           '0,
    jtag_rsp:           '0,
    prog_intg_err:      '0,
    storage_relbl_err:  '0,
    storage_intg_err:   '0,
    fsm_err:            '0,
    spurious_ack:       '0,
    arb_err:            '0,
    host_gnt_err:       '0,
    fifo_err:           '0
  };

  // RMA entries
  typedef struct packed {
    logic [BankW-1:0] bank;
    flash_part_e part;
    logic [InfoTypesWidth-1:0] info_sel;
    logic [PageW:0] start_page;
    logic [PageW:0] num_pages;
  } rma_wipe_entry_t;

  // entries to be wiped
  parameter int WipeEntries = 5;
  parameter rma_wipe_entry_t RmaWipeEntries[WipeEntries] = '{
    '{
       bank: SeedBank,
       part: FlashPartInfo,
       info_sel: SeedInfoSel,
       start_page: {1'b0, CreatorInfoPage},
       num_pages: 1
     },

    '{
       bank: SeedBank,
       part: FlashPartInfo,
       info_sel: SeedInfoSel,
       start_page: {1'b0, OwnerInfoPage},
       num_pages: 1
     },

    '{
       bank: SeedBank,
       part: FlashPartInfo,
       info_sel: SeedInfoSel,
       start_page: {1'b0, IsolatedInfoPage},
       num_pages: 1
     },

    '{
       bank: 0,
       part: FlashPartData,
       info_sel: 0,
       start_page: 0,
       num_pages: (PageW + 1)'(PagesPerBank)
     },

    '{
       bank: 1,
       part: FlashPartData,
       info_sel: 0,
       start_page: 0,
       num_pages: (PageW + 1)'(PagesPerBank)
     }
  };


  // flash_ctrl to keymgr
  typedef struct packed {
    logic [NumSeeds-1:0][SeedWidth-1:0] seeds;
  } keymgr_flash_t;

  parameter keymgr_flash_t KEYMGR_FLASH_DEFAULT = '{
    seeds: '{
     256'h9152e32c9380a4bcc3e0ab263581e6b0e8825186e1e445631646e8bef8c45d47,
     256'hfa365df52da48cd752fb3a026a8e608f0098cfe5fa9810494829d0cd9479eb78
    }
  };

  // dft_en jtag selection
  typedef enum logic [2:0] {
    FlashLcTckSel,
    FlashLcTdiSel,
    FlashLcTmsSel,
    FlashLcTdoSel,
    FlashBistSel,
    FlashLcDftLast
  } flash_lc_jtag_e;

  // Error bit positioning
  typedef struct packed {
    logic invalid_op_err;
    logic oob_err;
    logic mp_err;
    logic rd_err;
    logic prog_err;
    logic prog_win_err;
    logic prog_type_err;
  } flash_ctrl_err_t;

  // interrupt bit positioning
  typedef enum logic[2:0] {
    ProgEmpty,
    ProgLvl,
    RdFull,
    RdLvl,
    OpDone,
    CorrErr,
    LastIntrIdx
  } flash_ctrl_intr_e;

  // find the max number pages among info types
  function automatic integer max_info_pages(int infos[InfoTypes]);
    int current_max = 0;
    for (int i = 0; i < InfoTypes; i++) begin
      if (infos[i] > current_max) begin
        current_max = infos[i];
      end
    end
    return current_max;
  endfunction // max_info_banks

  // RMA control FSM encoding
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 7 -n 10   //      -s 3319803877 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||||||| (47.62%)
  //  6: |||||||||||||||| (38.10%)
  //  7: |||| (9.52%)
  //  8: || (4.76%)
  //  9: --
  // 10: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 8
  // Minimum Hamming weight: 3
  // Maximum Hamming weight: 6
  //
  localparam int RmaStateWidth = 11;
  typedef enum logic [RmaStateWidth-1:0] {
    StRmaIdle        = 11'b11110001010,
    StRmaPageSel     = 11'b10111100111,
    StRmaErase       = 11'b11000010111,
    StRmaEraseWait   = 11'b01010100110,
    StRmaWordSel     = 11'b00010011001,
    StRmaProgram     = 11'b11011111101,
    StRmaProgramWait = 11'b00111110000,
    StRmaRdVerify    = 11'b00101001100,
    StRmaDisabled    = 11'b01001011010,
    StRmaInvalid     = 11'b10100111011
  } rma_state_e;


  // find the max number pages among info types
  function automatic info_page_cfg_t info_cfg_qual(info_page_cfg_t in_cfg,
                                                   info_page_cfg_t qual_cfg);

    info_page_cfg_t out_cfg;
    out_cfg = '{
      en:          prim_mubi_pkg::mubi4_and_hi(in_cfg.en,          qual_cfg.en),
      rd_en:       prim_mubi_pkg::mubi4_and_hi(in_cfg.rd_en,       qual_cfg.rd_en),
      prog_en:     prim_mubi_pkg::mubi4_and_hi(in_cfg.prog_en,     qual_cfg.prog_en),
      erase_en:    prim_mubi_pkg::mubi4_and_hi(in_cfg.erase_en,    qual_cfg.erase_en),
      scramble_en: prim_mubi_pkg::mubi4_and_hi(in_cfg.scramble_en, qual_cfg.scramble_en),
      ecc_en:      prim_mubi_pkg::mubi4_and_hi(in_cfg.ecc_en,      qual_cfg.ecc_en),
      he_en :      prim_mubi_pkg::mubi4_and_hi(in_cfg.he_en,       qual_cfg.he_en)
    };

    return out_cfg;
  endfunction // max_info_banks

endpackage : flash_ctrl_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package keymgr_reg_pkg;

  // Param list
  parameter int NumSaltReg = 8;
  parameter int NumSwBindingReg = 8;
  parameter int NumOutReg = 8;
  parameter int NumKeyVersion = 1;
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 8;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    logic        q;
  } keymgr_reg2hw_intr_state_reg_t;

  typedef struct packed {
    logic        q;
  } keymgr_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    logic        q;
    logic        qe;
  } keymgr_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_operation_err;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_fault_err;
  } keymgr_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic        q;
  } keymgr_reg2hw_start_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  q;
    } operation;
    struct packed {
      logic        q;
    } cdi_sel;
    struct packed {
      logic [1:0]  q;
    } dest_sel;
  } keymgr_reg2hw_control_shadowed_reg_t;

  typedef struct packed {
    logic [2:0]  q;
  } keymgr_reg2hw_sideload_clear_reg_t;

  typedef struct packed {
    logic [15:0] q;
  } keymgr_reg2hw_reseed_interval_shadowed_reg_t;

  typedef struct packed {
    logic        q;
    logic        qe;
  } keymgr_reg2hw_sw_binding_regwen_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_sealing_sw_binding_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_attest_sw_binding_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_salt_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_key_version_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_max_creator_key_ver_shadowed_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_max_owner_int_key_ver_shadowed_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } keymgr_reg2hw_max_owner_key_ver_shadowed_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } cmd;
    struct packed {
      logic        q;
    } kmac_fsm;
    struct packed {
      logic        q;
    } kmac_done;
    struct packed {
      logic        q;
    } kmac_op;
    struct packed {
      logic        q;
    } kmac_out;
    struct packed {
      logic        q;
    } regfile_intg;
    struct packed {
      logic        q;
    } shadow;
    struct packed {
      logic        q;
    } ctrl_fsm_intg;
    struct packed {
      logic        q;
    } ctrl_fsm_chk;
    struct packed {
      logic        q;
    } ctrl_fsm_cnt;
    struct packed {
      logic        q;
    } reseed_cnt;
    struct packed {
      logic        q;
    } side_ctrl_fsm;
    struct packed {
      logic        q;
    } side_ctrl_sel;
    struct packed {
      logic        q;
    } key_ecc;
  } keymgr_reg2hw_fault_status_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } keymgr_hw2reg_intr_state_reg_t;

  typedef struct packed {
    logic        d;
  } keymgr_hw2reg_cfg_regwen_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } keymgr_hw2reg_start_reg_t;

  typedef struct packed {
    logic        d;
  } keymgr_hw2reg_sw_binding_regwen_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } keymgr_hw2reg_sw_share0_output_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } keymgr_hw2reg_sw_share1_output_mreg_t;

  typedef struct packed {
    logic [2:0]  d;
    logic        de;
  } keymgr_hw2reg_working_state_reg_t;

  typedef struct packed {
    logic [1:0]  d;
    logic        de;
  } keymgr_hw2reg_op_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } invalid_op;
    struct packed {
      logic        d;
      logic        de;
    } invalid_kmac_input;
    struct packed {
      logic        d;
      logic        de;
    } invalid_shadow_update;
  } keymgr_hw2reg_err_code_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } cmd;
    struct packed {
      logic        d;
      logic        de;
    } kmac_fsm;
    struct packed {
      logic        d;
      logic        de;
    } kmac_done;
    struct packed {
      logic        d;
      logic        de;
    } kmac_op;
    struct packed {
      logic        d;
      logic        de;
    } kmac_out;
    struct packed {
      logic        d;
      logic        de;
    } regfile_intg;
    struct packed {
      logic        d;
      logic        de;
    } shadow;
    struct packed {
      logic        d;
      logic        de;
    } ctrl_fsm_intg;
    struct packed {
      logic        d;
      logic        de;
    } ctrl_fsm_chk;
    struct packed {
      logic        d;
      logic        de;
    } ctrl_fsm_cnt;
    struct packed {
      logic        d;
      logic        de;
    } reseed_cnt;
    struct packed {
      logic        d;
      logic        de;
    } side_ctrl_fsm;
    struct packed {
      logic        d;
      logic        de;
    } side_ctrl_sel;
    struct packed {
      logic        d;
      logic        de;
    } key_ecc;
  } keymgr_hw2reg_fault_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } invalid_creator_seed;
    struct packed {
      logic        d;
      logic        de;
    } invalid_owner_seed;
    struct packed {
      logic        d;
      logic        de;
    } invalid_dev_id;
    struct packed {
      logic        d;
      logic        de;
    } invalid_health_state;
    struct packed {
      logic        d;
      logic        de;
    } invalid_key_version;
    struct packed {
      logic        d;
      logic        de;
    } invalid_key;
    struct packed {
      logic        d;
      logic        de;
    } invalid_digest;
  } keymgr_hw2reg_debug_reg_t;

  // Register -> HW type
  typedef struct packed {
    keymgr_reg2hw_intr_state_reg_t intr_state; // [945:945]
    keymgr_reg2hw_intr_enable_reg_t intr_enable; // [944:944]
    keymgr_reg2hw_intr_test_reg_t intr_test; // [943:942]
    keymgr_reg2hw_alert_test_reg_t alert_test; // [941:938]
    keymgr_reg2hw_start_reg_t start; // [937:937]
    keymgr_reg2hw_control_shadowed_reg_t control_shadowed; // [936:931]
    keymgr_reg2hw_sideload_clear_reg_t sideload_clear; // [930:928]
    keymgr_reg2hw_reseed_interval_shadowed_reg_t reseed_interval_shadowed; // [927:912]
    keymgr_reg2hw_sw_binding_regwen_reg_t sw_binding_regwen; // [911:910]
    keymgr_reg2hw_sealing_sw_binding_mreg_t [7:0] sealing_sw_binding; // [909:654]
    keymgr_reg2hw_attest_sw_binding_mreg_t [7:0] attest_sw_binding; // [653:398]
    keymgr_reg2hw_salt_mreg_t [7:0] salt; // [397:142]
    keymgr_reg2hw_key_version_mreg_t [0:0] key_version; // [141:110]
    keymgr_reg2hw_max_creator_key_ver_shadowed_reg_t max_creator_key_ver_shadowed; // [109:78]
    keymgr_reg2hw_max_owner_int_key_ver_shadowed_reg_t max_owner_int_key_ver_shadowed; // [77:46]
    keymgr_reg2hw_max_owner_key_ver_shadowed_reg_t max_owner_key_ver_shadowed; // [45:14]
    keymgr_reg2hw_fault_status_reg_t fault_status; // [13:0]
  } keymgr_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    keymgr_hw2reg_intr_state_reg_t intr_state; // [588:587]
    keymgr_hw2reg_cfg_regwen_reg_t cfg_regwen; // [586:586]
    keymgr_hw2reg_start_reg_t start; // [585:584]
    keymgr_hw2reg_sw_binding_regwen_reg_t sw_binding_regwen; // [583:583]
    keymgr_hw2reg_sw_share0_output_mreg_t [7:0] sw_share0_output; // [582:319]
    keymgr_hw2reg_sw_share1_output_mreg_t [7:0] sw_share1_output; // [318:55]
    keymgr_hw2reg_working_state_reg_t working_state; // [54:51]
    keymgr_hw2reg_op_status_reg_t op_status; // [50:48]
    keymgr_hw2reg_err_code_reg_t err_code; // [47:42]
    keymgr_hw2reg_fault_status_reg_t fault_status; // [41:14]
    keymgr_hw2reg_debug_reg_t debug; // [13:0]
  } keymgr_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] KEYMGR_INTR_STATE_OFFSET = 8'h 0;
  parameter logic [BlockAw-1:0] KEYMGR_INTR_ENABLE_OFFSET = 8'h 4;
  parameter logic [BlockAw-1:0] KEYMGR_INTR_TEST_OFFSET = 8'h 8;
  parameter logic [BlockAw-1:0] KEYMGR_ALERT_TEST_OFFSET = 8'h c;
  parameter logic [BlockAw-1:0] KEYMGR_CFG_REGWEN_OFFSET = 8'h 10;
  parameter logic [BlockAw-1:0] KEYMGR_START_OFFSET = 8'h 14;
  parameter logic [BlockAw-1:0] KEYMGR_CONTROL_SHADOWED_OFFSET = 8'h 18;
  parameter logic [BlockAw-1:0] KEYMGR_SIDELOAD_CLEAR_OFFSET = 8'h 1c;
  parameter logic [BlockAw-1:0] KEYMGR_RESEED_INTERVAL_REGWEN_OFFSET = 8'h 20;
  parameter logic [BlockAw-1:0] KEYMGR_RESEED_INTERVAL_SHADOWED_OFFSET = 8'h 24;
  parameter logic [BlockAw-1:0] KEYMGR_SW_BINDING_REGWEN_OFFSET = 8'h 28;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_0_OFFSET = 8'h 2c;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_1_OFFSET = 8'h 30;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_2_OFFSET = 8'h 34;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_3_OFFSET = 8'h 38;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_4_OFFSET = 8'h 3c;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_5_OFFSET = 8'h 40;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_6_OFFSET = 8'h 44;
  parameter logic [BlockAw-1:0] KEYMGR_SEALING_SW_BINDING_7_OFFSET = 8'h 48;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_0_OFFSET = 8'h 4c;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_1_OFFSET = 8'h 50;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_2_OFFSET = 8'h 54;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_3_OFFSET = 8'h 58;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_4_OFFSET = 8'h 5c;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_5_OFFSET = 8'h 60;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_6_OFFSET = 8'h 64;
  parameter logic [BlockAw-1:0] KEYMGR_ATTEST_SW_BINDING_7_OFFSET = 8'h 68;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_0_OFFSET = 8'h 6c;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_1_OFFSET = 8'h 70;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_2_OFFSET = 8'h 74;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_3_OFFSET = 8'h 78;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_4_OFFSET = 8'h 7c;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_5_OFFSET = 8'h 80;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_6_OFFSET = 8'h 84;
  parameter logic [BlockAw-1:0] KEYMGR_SALT_7_OFFSET = 8'h 88;
  parameter logic [BlockAw-1:0] KEYMGR_KEY_VERSION_OFFSET = 8'h 8c;
  parameter logic [BlockAw-1:0] KEYMGR_MAX_CREATOR_KEY_VER_REGWEN_OFFSET = 8'h 90;
  parameter logic [BlockAw-1:0] KEYMGR_MAX_CREATOR_KEY_VER_SHADOWED_OFFSET = 8'h 94;
  parameter logic [BlockAw-1:0] KEYMGR_MAX_OWNER_INT_KEY_VER_REGWEN_OFFSET = 8'h 98;
  parameter logic [BlockAw-1:0] KEYMGR_MAX_OWNER_INT_KEY_VER_SHADOWED_OFFSET = 8'h 9c;
  parameter logic [BlockAw-1:0] KEYMGR_MAX_OWNER_KEY_VER_REGWEN_OFFSET = 8'h a0;
  parameter logic [BlockAw-1:0] KEYMGR_MAX_OWNER_KEY_VER_SHADOWED_OFFSET = 8'h a4;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_0_OFFSET = 8'h a8;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_1_OFFSET = 8'h ac;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_2_OFFSET = 8'h b0;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_3_OFFSET = 8'h b4;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_4_OFFSET = 8'h b8;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_5_OFFSET = 8'h bc;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_6_OFFSET = 8'h c0;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE0_OUTPUT_7_OFFSET = 8'h c4;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_0_OFFSET = 8'h c8;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_1_OFFSET = 8'h cc;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_2_OFFSET = 8'h d0;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_3_OFFSET = 8'h d4;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_4_OFFSET = 8'h d8;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_5_OFFSET = 8'h dc;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_6_OFFSET = 8'h e0;
  parameter logic [BlockAw-1:0] KEYMGR_SW_SHARE1_OUTPUT_7_OFFSET = 8'h e4;
  parameter logic [BlockAw-1:0] KEYMGR_WORKING_STATE_OFFSET = 8'h e8;
  parameter logic [BlockAw-1:0] KEYMGR_OP_STATUS_OFFSET = 8'h ec;
  parameter logic [BlockAw-1:0] KEYMGR_ERR_CODE_OFFSET = 8'h f0;
  parameter logic [BlockAw-1:0] KEYMGR_FAULT_STATUS_OFFSET = 8'h f4;
  parameter logic [BlockAw-1:0] KEYMGR_DEBUG_OFFSET = 8'h f8;

  // Reset values for hwext registers and their fields
  parameter logic [0:0] KEYMGR_INTR_TEST_RESVAL = 1'h 0;
  parameter logic [0:0] KEYMGR_INTR_TEST_OP_DONE_RESVAL = 1'h 0;
  parameter logic [1:0] KEYMGR_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] KEYMGR_ALERT_TEST_RECOV_OPERATION_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] KEYMGR_ALERT_TEST_FATAL_FAULT_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] KEYMGR_CFG_REGWEN_RESVAL = 1'h 1;
  parameter logic [0:0] KEYMGR_CFG_REGWEN_EN_RESVAL = 1'h 1;
  parameter logic [0:0] KEYMGR_SW_BINDING_REGWEN_RESVAL = 1'h 1;
  parameter logic [0:0] KEYMGR_SW_BINDING_REGWEN_EN_RESVAL = 1'h 1;

  // Register index
  typedef enum int {
    KEYMGR_INTR_STATE,
    KEYMGR_INTR_ENABLE,
    KEYMGR_INTR_TEST,
    KEYMGR_ALERT_TEST,
    KEYMGR_CFG_REGWEN,
    KEYMGR_START,
    KEYMGR_CONTROL_SHADOWED,
    KEYMGR_SIDELOAD_CLEAR,
    KEYMGR_RESEED_INTERVAL_REGWEN,
    KEYMGR_RESEED_INTERVAL_SHADOWED,
    KEYMGR_SW_BINDING_REGWEN,
    KEYMGR_SEALING_SW_BINDING_0,
    KEYMGR_SEALING_SW_BINDING_1,
    KEYMGR_SEALING_SW_BINDING_2,
    KEYMGR_SEALING_SW_BINDING_3,
    KEYMGR_SEALING_SW_BINDING_4,
    KEYMGR_SEALING_SW_BINDING_5,
    KEYMGR_SEALING_SW_BINDING_6,
    KEYMGR_SEALING_SW_BINDING_7,
    KEYMGR_ATTEST_SW_BINDING_0,
    KEYMGR_ATTEST_SW_BINDING_1,
    KEYMGR_ATTEST_SW_BINDING_2,
    KEYMGR_ATTEST_SW_BINDING_3,
    KEYMGR_ATTEST_SW_BINDING_4,
    KEYMGR_ATTEST_SW_BINDING_5,
    KEYMGR_ATTEST_SW_BINDING_6,
    KEYMGR_ATTEST_SW_BINDING_7,
    KEYMGR_SALT_0,
    KEYMGR_SALT_1,
    KEYMGR_SALT_2,
    KEYMGR_SALT_3,
    KEYMGR_SALT_4,
    KEYMGR_SALT_5,
    KEYMGR_SALT_6,
    KEYMGR_SALT_7,
    KEYMGR_KEY_VERSION,
    KEYMGR_MAX_CREATOR_KEY_VER_REGWEN,
    KEYMGR_MAX_CREATOR_KEY_VER_SHADOWED,
    KEYMGR_MAX_OWNER_INT_KEY_VER_REGWEN,
    KEYMGR_MAX_OWNER_INT_KEY_VER_SHADOWED,
    KEYMGR_MAX_OWNER_KEY_VER_REGWEN,
    KEYMGR_MAX_OWNER_KEY_VER_SHADOWED,
    KEYMGR_SW_SHARE0_OUTPUT_0,
    KEYMGR_SW_SHARE0_OUTPUT_1,
    KEYMGR_SW_SHARE0_OUTPUT_2,
    KEYMGR_SW_SHARE0_OUTPUT_3,
    KEYMGR_SW_SHARE0_OUTPUT_4,
    KEYMGR_SW_SHARE0_OUTPUT_5,
    KEYMGR_SW_SHARE0_OUTPUT_6,
    KEYMGR_SW_SHARE0_OUTPUT_7,
    KEYMGR_SW_SHARE1_OUTPUT_0,
    KEYMGR_SW_SHARE1_OUTPUT_1,
    KEYMGR_SW_SHARE1_OUTPUT_2,
    KEYMGR_SW_SHARE1_OUTPUT_3,
    KEYMGR_SW_SHARE1_OUTPUT_4,
    KEYMGR_SW_SHARE1_OUTPUT_5,
    KEYMGR_SW_SHARE1_OUTPUT_6,
    KEYMGR_SW_SHARE1_OUTPUT_7,
    KEYMGR_WORKING_STATE,
    KEYMGR_OP_STATUS,
    KEYMGR_ERR_CODE,
    KEYMGR_FAULT_STATUS,
    KEYMGR_DEBUG
  } keymgr_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] KEYMGR_PERMIT [63] = '{
    4'b 0001, // index[ 0] KEYMGR_INTR_STATE
    4'b 0001, // index[ 1] KEYMGR_INTR_ENABLE
    4'b 0001, // index[ 2] KEYMGR_INTR_TEST
    4'b 0001, // index[ 3] KEYMGR_ALERT_TEST
    4'b 0001, // index[ 4] KEYMGR_CFG_REGWEN
    4'b 0001, // index[ 5] KEYMGR_START
    4'b 0011, // index[ 6] KEYMGR_CONTROL_SHADOWED
    4'b 0001, // index[ 7] KEYMGR_SIDELOAD_CLEAR
    4'b 0001, // index[ 8] KEYMGR_RESEED_INTERVAL_REGWEN
    4'b 0011, // index[ 9] KEYMGR_RESEED_INTERVAL_SHADOWED
    4'b 0001, // index[10] KEYMGR_SW_BINDING_REGWEN
    4'b 1111, // index[11] KEYMGR_SEALING_SW_BINDING_0
    4'b 1111, // index[12] KEYMGR_SEALING_SW_BINDING_1
    4'b 1111, // index[13] KEYMGR_SEALING_SW_BINDING_2
    4'b 1111, // index[14] KEYMGR_SEALING_SW_BINDING_3
    4'b 1111, // index[15] KEYMGR_SEALING_SW_BINDING_4
    4'b 1111, // index[16] KEYMGR_SEALING_SW_BINDING_5
    4'b 1111, // index[17] KEYMGR_SEALING_SW_BINDING_6
    4'b 1111, // index[18] KEYMGR_SEALING_SW_BINDING_7
    4'b 1111, // index[19] KEYMGR_ATTEST_SW_BINDING_0
    4'b 1111, // index[20] KEYMGR_ATTEST_SW_BINDING_1
    4'b 1111, // index[21] KEYMGR_ATTEST_SW_BINDING_2
    4'b 1111, // index[22] KEYMGR_ATTEST_SW_BINDING_3
    4'b 1111, // index[23] KEYMGR_ATTEST_SW_BINDING_4
    4'b 1111, // index[24] KEYMGR_ATTEST_SW_BINDING_5
    4'b 1111, // index[25] KEYMGR_ATTEST_SW_BINDING_6
    4'b 1111, // index[26] KEYMGR_ATTEST_SW_BINDING_7
    4'b 1111, // index[27] KEYMGR_SALT_0
    4'b 1111, // index[28] KEYMGR_SALT_1
    4'b 1111, // index[29] KEYMGR_SALT_2
    4'b 1111, // index[30] KEYMGR_SALT_3
    4'b 1111, // index[31] KEYMGR_SALT_4
    4'b 1111, // index[32] KEYMGR_SALT_5
    4'b 1111, // index[33] KEYMGR_SALT_6
    4'b 1111, // index[34] KEYMGR_SALT_7
    4'b 1111, // index[35] KEYMGR_KEY_VERSION
    4'b 0001, // index[36] KEYMGR_MAX_CREATOR_KEY_VER_REGWEN
    4'b 1111, // index[37] KEYMGR_MAX_CREATOR_KEY_VER_SHADOWED
    4'b 0001, // index[38] KEYMGR_MAX_OWNER_INT_KEY_VER_REGWEN
    4'b 1111, // index[39] KEYMGR_MAX_OWNER_INT_KEY_VER_SHADOWED
    4'b 0001, // index[40] KEYMGR_MAX_OWNER_KEY_VER_REGWEN
    4'b 1111, // index[41] KEYMGR_MAX_OWNER_KEY_VER_SHADOWED
    4'b 1111, // index[42] KEYMGR_SW_SHARE0_OUTPUT_0
    4'b 1111, // index[43] KEYMGR_SW_SHARE0_OUTPUT_1
    4'b 1111, // index[44] KEYMGR_SW_SHARE0_OUTPUT_2
    4'b 1111, // index[45] KEYMGR_SW_SHARE0_OUTPUT_3
    4'b 1111, // index[46] KEYMGR_SW_SHARE0_OUTPUT_4
    4'b 1111, // index[47] KEYMGR_SW_SHARE0_OUTPUT_5
    4'b 1111, // index[48] KEYMGR_SW_SHARE0_OUTPUT_6
    4'b 1111, // index[49] KEYMGR_SW_SHARE0_OUTPUT_7
    4'b 1111, // index[50] KEYMGR_SW_SHARE1_OUTPUT_0
    4'b 1111, // index[51] KEYMGR_SW_SHARE1_OUTPUT_1
    4'b 1111, // index[52] KEYMGR_SW_SHARE1_OUTPUT_2
    4'b 1111, // index[53] KEYMGR_SW_SHARE1_OUTPUT_3
    4'b 1111, // index[54] KEYMGR_SW_SHARE1_OUTPUT_4
    4'b 1111, // index[55] KEYMGR_SW_SHARE1_OUTPUT_5
    4'b 1111, // index[56] KEYMGR_SW_SHARE1_OUTPUT_6
    4'b 1111, // index[57] KEYMGR_SW_SHARE1_OUTPUT_7
    4'b 0001, // index[58] KEYMGR_WORKING_STATE
    4'b 0001, // index[59] KEYMGR_OP_STATUS
    4'b 0001, // index[60] KEYMGR_ERR_CODE
    4'b 0011, // index[61] KEYMGR_FAULT_STATUS
    4'b 0001  // index[62] KEYMGR_DEBUG
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// key manager package
//

package keymgr_pkg;

  parameter int KeyWidth = 256;
  parameter int CDIs = 2; // 2 different CDIs, sealing / attestation
  parameter int CdiWidth = prim_util_pkg::vbits(CDIs);
  parameter int OtbnKeyWidth = 384;
  parameter int DigestWidth = 128;     // uses truncated hash
  parameter int KmacDataIfWidth = 64;  // KMAC interface data width
  parameter int KeyMgrStages = 3; // Number of key manager stages (creator, ownerInt, owner)
  parameter int SwBindingWidth = 32 * keymgr_reg_pkg::NumSwBindingReg;
  parameter int SaltWidth = 32 * keymgr_reg_pkg::NumSaltReg;
  parameter int Shares = 2; // number of key shares
  parameter int EdnWidth = edn_pkg::ENDPOINT_BUS_WIDTH;

  // These should be defined in another module's package
  parameter int HealthStateWidth = 128;
  parameter int DevIdWidth = 256;
  parameter int MaxWidth = 256;

  // Default seeds
  // These are generated using random.org byte dumper
  typedef logic [KeyWidth-1:0] seed_t;
  parameter seed_t RndCnstRevisionSeedDefault =
    256'h3a0a6d73cd50897de4d744bd65ebdb3837ea77087d878651c517c18a5742b2f9;
  parameter seed_t RndCnstCreatorIdentitySeedDefault =
    256'h6d234651d535ebb0dce4d82f503096614355fc7b84595e4f67a866177d421df6;
  parameter seed_t RndCnstOwnerIntIdentitySeedDefault =
    256'hdba98db4fb1413b32fd5a4deac3ce546966a4bc2761235643358c8e76083d382;
  parameter seed_t RndCnstOwnerIdentitySeedDefault =
    256'h8c0a27ef53e0e0bf5f5f5e26a30a0d0db10761ed802c6d2fd22873209976021e;
  parameter seed_t RndCnstSoftOutputSeedDefault =
    256'h99cadb2c2d9b438591d943a89bc64dbb3bc2abc842eeea5faf74d27f7a7c99b6;
  parameter seed_t RndCnstHardOutputSeedDefault =
    256'hd551b351decbb6f687c7f5c845363f12d6411fae812e16b23bc8ae59885a56b1;

  // Target based deriviation seeds
  // These are used during the generation stages for sideload
  parameter seed_t RndCnstNoneSeedDefault =
    256'h6EECBF9FC3C64230421DA1EAEC48F871070A3582E71AD4059D5D550784E9B9DE;
  parameter seed_t RndCnstAesSeedDefault =
    256'hC1104CD94EBA084FA6438188038006489F3DF38771214AE0BBA65CEB9BC2366F;
  parameter seed_t RndCnstKmacSeedDefault =
    256'h0A5CCCD9627BF6169B3A765D3D6D0CD89DBDCB7B6DF8D3C03746D60A0145D3ED;
  parameter seed_t RndCnstOtbnSeedDefault =
    256'h17B0AF865F8ACDDFC7580C2B7BC3FB33FC9BB5A4B292216C123ACF99A7861F96;
  parameter seed_t RndCnstCdiDefault =
    256'hC69C544D153A692AEEC4A0887BD5255F5C588C63A8BD94479BCFF7432DC55E3B;

  // Default Lfsr configurations
  // These LFSR parameters have been generated with
  // $ util/design/gen-lfsr-seed.py --width 64 --seed 691876113 --prefix ""
  parameter int LfsrWidth = 64;
  typedef logic [LfsrWidth-1:0] lfsr_seed_t;
  typedef logic [LfsrWidth-1:0][$clog2(LfsrWidth)-1:0] lfsr_perm_t;
  parameter lfsr_seed_t RndCnstLfsrSeedDefault = 64'h22d326255bd24320;
  parameter lfsr_perm_t RndCnstLfsrPermDefault = {
    128'h16108c9f9008aa37e5118d1ec1df64a7,
    256'h24f3f1b73537f42d38383ee8f897286df81d49ab54b6bbbb666cbd1a16c41252
  };

  // Random permutation
  parameter int RandWidth = LfsrWidth / 2;
  typedef logic [RandWidth-1:0][$clog2(RandWidth)-1:0] rand_perm_t;
  parameter rand_perm_t RndCnstRandPermDefault = {
    160'h62089181d2a6be2ce145e2e27099ededbd7dceb0
  };

  // Width calculations
  // These are the largest calculations in use across all stages
  parameter int AdvDataWidth = SwBindingWidth + 3*KeyWidth + DevIdWidth + HealthStateWidth;
  parameter int IdDataWidth = KeyWidth;
  // key version + salt + key ID + constant
  parameter int GenDataWidth = 32 + SaltWidth + KeyWidth*2;
  parameter int StageWidth = $clog2(KeyMgrStages);
  // Max Payload Width to derivation function
  // see security strength description https://keccak.team/keccak.html
  // The max width here is chosen arbitrarily to ensure we do not get out of hand.
  // Since KMAC is a MAC operation, the data can be as long as we need.
  parameter int KDFMaxWidth = 1600;

  // Enumeration for operations
  typedef enum logic [1:0] {
    Creator,
    OwnerInt,
    Owner,
    Disable
  } keymgr_stage_e;

  // Enumeration for sideload sel
  typedef enum logic [1:0] {
    None,
    Aes,
    Kmac,
    Otbn
  } keymgr_key_dest_e;

  // Enumeration for actual key slot idx
  typedef enum logic [1:0] {
    AesIdx,
    KmacIdx,
    OtbnIdx,
    LastIdx
  } keymgr_sideload_slot_idx_e;

  // Enumeration for key select
  typedef enum logic {
    HwKey = 0,
    SwKey = 1
  } keymgr_gen_out_e;

  // Enumeration for operation
  typedef enum logic [2:0] {
    OpAdvance = 0,
    OpGenId = 1,
    OpGenSwOut = 2,
    OpGenHwOut = 3,
    OpDisable = 4
  } keymgr_ops_e;

  // Enumeration for working state exposed to software
  typedef enum logic [2:0] {
    StReset,
    StInit,
    StCreatorRootKey,
    StOwnerIntKey,
    StOwnerKey,
    StDisabled,
    StInvalid
  } keymgr_working_state_e;

  // Enumeration for operation status
  typedef enum logic [1:0] {
    OpIdle = 0,
    OpWip = 1,
    OpDoneSuccess = 2,
    OpDoneFail = 3
  } keymgr_op_status_e;

  // keymgr has 4 categories of errors
  // sync errors  - recoverable errors that happen during keymgr operation
  // async errors - recoverable errors that happen asynchronously
  // sync faults  - fatal errors that happen during keymgr operation
  // async faults - fatal errors that happen asynchronously

  typedef enum logic [1:0] {
    SyncErrInvalidOp,
    SyncErrInvalidIn,
    SyncErrLastIdx
  } keymgr_sync_error_e;

  typedef enum logic [1:0] {
    AsyncErrShadowUpdate,
    AsyncErrLastIdx
  } keymgr_async_error_e;

  typedef enum logic [1:0] {
    SyncFaultKmacOp,
    SyncFaultKmacOut,
    SyncFaultSideSel,
    SyncFaultLastIdx
  } keymgr_sync_fault_e;

  typedef enum logic [3:0] {
    AsyncFaultKmacCmd,
    AsyncFaultKmacFsm,
    AsyncFaultKmacDone,
    AsyncFaultRegIntg,
    AsyncFaultShadow,
    AsyncFaultFsmIntg,
    AsyncFaultFsmChk,
    AsyncFaultCntErr,
    AsyncFaultRCntErr,
    AsyncFaultSideErr,
    AsyncFaultKeyEcc,
    AsyncFaultLastIdx
  } keymgr_async_fault_e;


  // Bit position of error code
  // Error is encoded as 1 error per bit
  typedef enum logic [2:0] {
    ErrInvalidOp,
    ErrInvalidIn,
    ErrShadowUpdate,
    ErrLastPos
  } keymgr_err_pos_e;

  // Bit position of fault status
  typedef enum logic [3:0] {
    FaultKmacCmd,
    FaultKmacFsm,
    FaultKmacDone,
    FaultKmacOp,
    FaultKmacOut,
    FaultRegIntg,
    FaultShadow,
    FaultCtrlFsm,
    FaultCtrlFsmChk,
    FaultCtrlCnt,
    FaultReseedCnt,
    FaultSideFsm,
    FaultSideSel,
    FaultKeyEcc,
    FaultLastPos
  } keymgr_fault_pos_e;

  typedef enum logic [2:0] {
    KeyUpdateIdle,
    KeyUpdateRandom,
    KeyUpdateRoot,
    KeyUpdateKmac,
    KeyUpdateWipe
  } keymgr_key_update_e;

  typedef enum logic [2:0] {
    SideLoadClrIdle,
    SideLoadClrAes,
    SideLoadClrKmac,
    SideLoadClrOtbn
  } keymgr_sideload_clr_e;

  // Key connection to various symmetric modules
  typedef struct packed {
    logic valid;
    logic [Shares-1:0][KeyWidth-1:0] key;
  } hw_key_req_t;

  // Key connection to otbn
  typedef struct packed {
    logic valid;
    logic [Shares-1:0][OtbnKeyWidth-1:0] key;
  } otbn_key_req_t;

  parameter hw_key_req_t HW_KEY_REQ_DEFAULT = '{
    valid: 1'b0,
    key: {Shares{KeyWidth'(32'hDEADBEEF)}}
  };

  parameter otbn_key_req_t OTBN_KEY_REQ_DEFAULT = '{
    valid: 1'b0,
    key: {Shares{OtbnKeyWidth'(32'hDEADBEEF)}}
  };

  // The following structs should be sourced from other modules
  // defined here temporarily

  // lc keymgr enable usage
  typedef enum logic [1:0] {
    KeyMgrEnCtrl,
    KeyMgrEnCfgEn,
    KeyMgrEnSwBindingEn,
    KeyMgrEnLast
  } keymgr_lc_en_usage_e;

  // perm_data
  function automatic logic[RandWidth-1:0] perm_data (logic [RandWidth-1:0] data,
    rand_perm_t perm_sel);

    for (int k = 0; k < 32; k++) begin : gen_data_loop
      perm_data[k] = data[perm_sel[k]];
    end

  endfunction

endpackage : keymgr_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module can be used as a "gadget" to adapt the native 32bit width of the EDN network
// locally to the width needed by the consuming logic. For example, if the local consumer
// needs 128bit, this module would request four 32 bit words from EDN and stack them accordingly.
//
// The module also uses a req/ack synchronizer to synchronize the EDN data over to the local
// clock domain. Note that this assumes that the EDN data bus remains stable between subsequent
// requests.
//

`include "prim_assert.sv"

module prim_edn_req
  import prim_alert_pkg::*;
#(
  parameter int OutWidth = 32,
  // Repetition check for incoming edn data
  parameter bit RepCheck = 0,
  // Disable reset-related assertion checks inside prim_sync_reqack primitives.
  parameter bit EnRstChks = 0,

  // EDN Request latency checker
  //
  //  Each consumer IP may have the maximum expected latency. MaxLatency
  //  parameter describes the expected latency in terms of the consumer clock
  //  cycles. If the edn request comes later than that, the assertion will be
  //  fired.
  //
  //  The default value is 0, which disables the assertion.
  parameter int unsigned MaxLatency = 0
) (
  // Design side
  input                       clk_i,
  input                       rst_ni,
  input                       req_chk_i, // Used for gating assertions. Drive to 1 during normal
                                         // operation.
  input                       req_i,
  output logic                ack_o,
  output logic [OutWidth-1:0] data_o,
  output logic                fips_o,
  output logic                err_o,  // current data_o failed repetition check
  // EDN side
  input                       clk_edn_i,
  input                       rst_edn_ni,
  output edn_pkg::edn_req_t   edn_o,
  input  edn_pkg::edn_rsp_t   edn_i
);

  // Stop requesting words from EDN once desired amount of data is available.
  logic word_req, word_ack;
  assign word_req = req_i & ~ack_o;

  logic [edn_pkg::ENDPOINT_BUS_WIDTH-1:0] word_data;
  logic word_fips;
  localparam int SyncWidth = $bits({edn_i.edn_fips, edn_i.edn_bus});
  prim_sync_reqack_data #(
    .Width(SyncWidth),
    .EnRstChks(EnRstChks),
    .DataSrc2Dst(1'b0),
    .DataReg(1'b0)
  ) u_prim_sync_reqack_data (
    .clk_src_i  ( clk_i                           ),
    .rst_src_ni ( rst_ni                          ),
    .clk_dst_i  ( clk_edn_i                       ),
    .rst_dst_ni ( rst_edn_ni                      ),
    .req_chk_i  ( req_chk_i                       ),
    .src_req_i  ( word_req                        ),
    .src_ack_o  ( word_ack                        ),
    .dst_req_o  ( edn_o.edn_req                   ),
    .dst_ack_i  ( edn_i.edn_ack                   ),
    .data_i     ( {edn_i.edn_fips, edn_i.edn_bus} ),
    .data_o     ( {word_fips,      word_data}     )
  );

  if (RepCheck) begin : gen_rep_chk
    logic [edn_pkg::ENDPOINT_BUS_WIDTH-1:0] word_data_q;
    always_ff @(posedge clk_i) begin
      if (word_ack) begin
        word_data_q <= word_data;
      end
    end

    // do not check until we have received at least the first entry
    logic chk_rep;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        chk_rep <= '0;
      end else if (word_ack) begin
        chk_rep <= 1'b1;
      end
    end

    // Need to track if any of the packed words has failed the repetition check, i.e., is identical
    // to the last packed word.
    logic err_d, err_q;
    assign err_d = (req_i && ack_o)                                  ? 1'b0 : // clear
                   (chk_rep && word_ack && word_data == word_data_q) ? 1'b1 : // set
                                                                       err_q; // keep
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        err_q <= 1'b0;
      end else begin
        err_q <= err_d;
      end
    end
    assign err_o = err_q;

  end else begin : gen_no_rep_chk // block: gen_rep_chk
    assign err_o = '0;
  end

  prim_packer_fifo #(
    .InW(edn_pkg::ENDPOINT_BUS_WIDTH),
    .OutW(OutWidth),
    .ClearOnRead(1'b0)
  ) u_prim_packer_fifo (
    .clk_i,
    .rst_ni,
    .clr_i    ( 1'b0          ), // not needed
    .wvalid_i ( word_ack      ),
    .wdata_i  ( word_data     ),
    // no need for backpressure since we're always ready to
    // sink data at this point.
    .wready_o (               ),
    .rvalid_o ( ack_o         ),
    .rdata_o  ( data_o        ),
    // we're always ready to receive the packed output word
    // at this point.
    .rready_i ( 1'b1          ),
    .depth_o  (               )
  );

  // Need to track if any of the packed words has been generated with a pre-FIPS seed, i.e., has
  // fips == 1'b0.
  logic fips_d, fips_q;
  assign fips_d = (req_i && ack_o) ? 1'b1               : // clear
                  (word_ack)       ? fips_q & word_fips : // accumulate
                                     fips_q;              // keep
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      fips_q <= 1'b1;
    end else begin
      fips_q <= fips_d;
    end
  end
  assign fips_o = fips_q;

  ////////////////
  // Assertions //
  ////////////////

  // Check EDN data is valid: Not all zeros, all ones, or not the same as previous data.
`ifdef INC_ASSERT
  //VCS coverage off
  // pragma coverage off

  logic [OutWidth-1:0] data_prev, data_curr;

  always_ff @(posedge ack_o or negedge rst_ni) begin
    if (!rst_ni) begin
      data_prev <= '0;
      data_curr <= '0;
    end else if (ack_o) begin
      data_curr <= data_o;
      data_prev <= data_curr;
    end
  end
  //VCS coverage on
  // pragma coverage on

  `ASSERT(DataOutputValid_A, ack_o |-> (data_o != 0) && (data_o != '1))
  `ASSERT(DataOutputDiffFromPrev_A, data_prev != 0 |-> data_prev != data_o)
`endif

  // EDN Max Latency Checker
`ifndef SYNTHESIS
  if (MaxLatency != 0) begin: g_maxlatency_assertion
    //VCS coverage off
    // pragma coverage off
    localparam int unsigned LatencyW = $clog2(MaxLatency+1);
    logic [LatencyW-1:0] latency_counter;
    logic reset_counter;
    logic enable_counter;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) latency_counter <= '0;
      else if (reset_counter) latency_counter <= '0;
      else if (enable_counter) latency_counter <= latency_counter + 1'b1;
    end

    assign reset_counter  = ack_o;
    assign enable_counter = req_i;
    //VCS coverage on
    // pragma coverage on

    `ASSERT(MaxLatency_A, latency_counter <= MaxLatency)

    // TODO: Is it worth to check req & ack pair?
    //         _________________________________
    // req  __/                                 \______
    //                                           ____
    // ack  ____________________________________/    \_
    //
    //                                          | error

  end // g_maxlatency_assertion
`else // SYNTHESIS
  logic unused_param_maxlatency;
  assign unused_param_maxlatency = ^MaxLatency;
`endif // SYNTHESIS

endmodule : prim_edn_req


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL adapter for Register interface
 *
 * ICEBOX(#15822): Note that due to some modules with special needs (like
 * the vendored-in RV_DM), this module has been extended so that it
 * supports use cases outside of the generated reg_top module. This makes
 * this adapter and its parameterization options a bit heavy.
 *
 * We should in the future come back to this and refactor / align the
 * module and its parameterization needs.
 */

module tlul_adapter_reg
  import tlul_pkg::*;
  import prim_mubi_pkg::mubi4_t;
#(
  parameter  bit CmdIntgCheck      = 0,  // 1: Enable command integrity check
  parameter  bit EnableRspIntgGen  = 0,  // 1: Generate response integrity
  parameter  bit EnableDataIntgGen = 0,  // 1: Generate response data integrity
  parameter  int RegAw             = 8,  // Width of register address
  parameter  int RegDw             = 32, // Shall be matched with TL_DW
  parameter  int AccessLatency     = 0,  // 0: same cycle, 1: next cycle
  localparam int RegBw             = RegDw/8
) (
  input clk_i,
  input rst_ni,

  // TL-UL interface
  input  tl_h2d_t tl_i,
  output tl_d2h_t tl_o,

  // control interface
  input  mubi4_t  en_ifetch_i,
  output logic    intg_error_o,

  // Register interface
  output logic             re_o,
  output logic             we_o,
  output logic [RegAw-1:0] addr_o,
  output logic [RegDw-1:0] wdata_o,
  output logic [RegBw-1:0] be_o,
  input                    busy_i,
  // The following two signals are expected
  // to be returned in AccessLatency cycles.
  input        [RegDw-1:0] rdata_i,
  // This can be a write or read error.
  input                    error_i
);

  `ASSERT_INIT(AllowedLatency_A, AccessLatency inside {0, 1})

  localparam int IW  = $bits(tl_i.a_source);
  localparam int SZW = $bits(tl_i.a_size);

  logic outstanding_q;    // Indicates current request is pending
  logic a_ack, d_ack;

  logic [RegDw-1:0] rdata, rdata_q;
  logic             error_q, error, err_internal, instr_error, intg_error;

  logic addr_align_err;     // Size and alignment
  logic malformed_meta_err; // User signal format error or unsupported
  logic tl_err;             // Common TL-UL error checker

  logic [IW-1:0]  reqid_q;
  logic [SZW-1:0] reqsz_q;
  tl_d_op_e       rspop_q;

  logic rd_req, wr_req;

  assign a_ack   = tl_i.a_valid & tl_o.a_ready;
  assign d_ack   = tl_o.d_valid & tl_i.d_ready;
  // Request signal
  assign wr_req  = a_ack & ((tl_i.a_opcode == PutFullData) | (tl_i.a_opcode == PutPartialData));
  assign rd_req  = a_ack & (tl_i.a_opcode == Get);

  assign we_o    = wr_req & ~err_internal;
  assign re_o    = rd_req & ~err_internal;
  assign wdata_o = tl_i.a_data;
  assign be_o    = tl_i.a_mask;

  if (RegAw <= 2) begin : gen_only_one_reg
    assign addr_o  = '0;
  end else begin : gen_more_regs
    assign addr_o  = {tl_i.a_address[RegAw-1:2], 2'b00}; // generate always word-align
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)    outstanding_q <= 1'b0;
    else if (a_ack) outstanding_q <= 1'b1;
    else if (d_ack) outstanding_q <= 1'b0;
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      reqid_q <= '0;
      reqsz_q <= '0;
      rspop_q <= AccessAck;
    end else if (a_ack) begin
      reqid_q <= tl_i.a_source;
      reqsz_q <= tl_i.a_size;
      // Return AccessAckData regardless of error
      rspop_q <= (rd_req) ? AccessAckData : AccessAck ;
    end
  end

  if (AccessLatency == 1) begin : gen_access_latency1
    logic wr_req_q, rd_req_q;
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        rdata_q  <= '0;
        error_q  <= 1'b0;
        wr_req_q <= 1'b0;
        rd_req_q <= 1'b0;
      end else begin
        rd_req_q <= rd_req;
        wr_req_q <= wr_req;
        // Addressing phase
        if (a_ack) begin
          error_q <= err_internal;
        // Response phase
        end else begin
          error_q <= error;
          rdata_q <= rdata;
        end
      end
    end
    assign rdata = (error_i || error_q || wr_req_q) ? '1      :
                   (rd_req_q)                       ? rdata_i :
                                                      rdata_q; // backpressure case
    assign error = (rd_req_q || wr_req_q) ? (error_q || error_i) :
                                            error_q; // backpressure case
  end else begin : gen_access_latency0
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        rdata_q <= '0;
        error_q <= 1'b0;
      end else if (a_ack) begin
        rdata_q <= (error_i || err_internal || wr_req) ? '1 : rdata_i;
        error_q <= error_i || err_internal;
      end
    end
    assign rdata = rdata_q;
    assign error = error_q;
  end

  tlul_pkg::tl_d2h_t tl_o_pre;
  assign tl_o_pre = '{
    // busy is selected based on address
    // thus if there is no valid transaction, we should ignore busy
    a_ready:  ~(outstanding_q | tl_i.a_valid & busy_i),
    d_valid:  outstanding_q,
    d_opcode: rspop_q,
    d_param:  '0,
    d_size:   reqsz_q,
    d_source: reqid_q,
    d_sink:   '0,
    d_data:   rdata,
    d_user:   '0,
    d_error:  error
  };

  // outgoing integrity generation
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(EnableRspIntgGen),
    .EnableDataIntgGen(EnableDataIntgGen)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  if (CmdIntgCheck) begin : gen_cmd_intg_check
    logic intg_error_q;
    tlul_cmd_intg_chk u_cmd_intg_chk (
      .tl_i(tl_i),
      .err_o(intg_error)
    );
    // permanently latch integrity error until reset
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        intg_error_q <= 1'b0;
      end else if (intg_error) begin
        intg_error_q <= 1'b1;
      end
    end
    assign intg_error_o = intg_error_q;
  end else begin : gen_no_cmd_intg_check
    assign intg_error = 1'b0;
    assign intg_error_o = 1'b0;
  end

  ////////////////////
  // Error Handling //
  ////////////////////

  // An instruction type transaction is only valid if en_ifetch is enabled
  // If the instruction type is completely invalid, also considered an instruction error
  assign instr_error = prim_mubi_pkg::mubi4_test_invalid(tl_i.a_user.instr_type) |
                       (prim_mubi_pkg::mubi4_test_true_strict(tl_i.a_user.instr_type) &
                        prim_mubi_pkg::mubi4_test_false_loose(en_ifetch_i));

  assign err_internal = addr_align_err | malformed_meta_err | tl_err | instr_error | intg_error;

  // Don't allow unsupported values.
  assign malformed_meta_err = tl_a_user_chk(tl_i.a_user);

  // addr_align_err
  //    Raised if addr isn't aligned with the size
  //    Read size error is checked in tlul_assert.sv
  //    Here is it added due to the limitation of register interface.
  always_comb begin
    if (wr_req) begin
      // Only word-align is accepted based on comportability spec
      addr_align_err = |tl_i.a_address[1:0];
    end else begin
      // No request
      addr_align_err = 1'b0;
    end
  end

  // tl_err : separate checker
  tlul_err u_err (
    .clk_i,
    .rst_ni,
    .tl_i,
    .err_o (tl_err)
  );

  `ASSERT_INIT(MatchedWidthAssert, RegDw == top_pkg::TL_DW)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL adapter for SRAM-like devices
 *
 * This module handles byte writes for tlul integrity.
 * When a byte write is received, the downstream data is read first
 * to correctly create the integrity constant.
 *
 * A tlul transaction goes through this module.  If required, a
 * tlul read transaction is generated out first.  If not required, the
 * incoming tlul transaction is directly muxed out.
 */
module tlul_sram_byte import tlul_pkg::*; #(
  parameter bit EnableIntg  = 0,  // Enable integrity handling at byte level
  parameter int Outstanding = 1
) (
  input clk_i,
  input rst_ni,

  input tl_h2d_t tl_i,
  output tl_d2h_t tl_o,

  output tl_h2d_t tl_sram_o,
  input tl_d2h_t tl_sram_i,

  // if incoming transaction already has an error, do not
  // attempt to handle the byte-write access.  Instead treat as
  // feedthrough and allow the system to directly error back.
  // The error indication is also fed through
  input error_i,
  output logic error_o
);

  if (EnableIntg) begin : gen_integ_handling

    // state enumeration
    typedef enum logic [1:0] {
      StPassThru,
      StWaitRd,
      StWriteCmd
    } state_e;

    // state and selection
    logic stall_host;
    logic rd_phase;
    logic rd_wait;
    logic wr_phase;
    state_e state_d, state_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        state_q <= StPassThru;
      end else begin
        state_q <= state_d;
      end
    end

    // transaction qualifying signals
    logic a_ack;  // upstream a channel acknowledgement
    logic d_ack;  // upstream d channel acknowledgement
    logic sram_a_ack; // downstream a channel acknowledgement
    logic sram_d_ack; // downstream d channel acknowledgement
    logic wr_txn;
    logic byte_wr_txn;
    logic byte_req_ack;
    logic [prim_util_pkg::vbits(Outstanding+1)-1:0] pending_txn_cnt;

    assign a_ack = tl_i.a_valid & tl_o.a_ready;
    assign d_ack = tl_o.d_valid & tl_i.d_ready;
    assign sram_a_ack = tl_sram_o.a_valid & tl_sram_i.a_ready;
    assign sram_d_ack = tl_sram_i.d_valid & tl_sram_o.d_ready;
    assign wr_txn = (tl_i.a_opcode == PutFullData) | (tl_i.a_opcode == PutPartialData);

    assign byte_req_ack = byte_wr_txn & a_ack & ~error_i;
    assign byte_wr_txn = tl_i.a_valid & ~&tl_i.a_mask & wr_txn;

    // state machine handling
    always_comb begin
      rd_wait = 1'b0;
      stall_host = 1'b0;
      wr_phase = 1'b0;
      rd_phase = 1'b0;
      state_d = state_q;

      unique case (state_q)
        StPassThru: begin
          if (byte_wr_txn) begin
            rd_phase = 1'b1;
            if (byte_req_ack) begin
              state_d = StWaitRd;
            end
          end
        end

        // Due to the way things are serialized, there is no way for the logic to tell which read
        // belongs to the partial read unless it flushes all prior transactions. Hence, we wait
        // here until exactly one outstanding transaction remains (that one is the partial read).
        StWaitRd: begin
          rd_phase = 1'b1;
          stall_host = 1'b1;
          if (pending_txn_cnt == $bits(pending_txn_cnt)'(1)) begin
            rd_wait = 1'b1;
            if (sram_d_ack) begin
              state_d = StWriteCmd;
            end
          end
        end

        StWriteCmd: begin
          stall_host = 1'b1;
          wr_phase = 1'b1;

          if (sram_a_ack) begin
            state_d = StPassThru;
          end
        end

        default:;

      endcase // unique case (state_q)

    end

    // prim fifo for capturing info
    typedef struct packed {
      logic                  [2:0]  a_param;
      logic  [top_pkg::TL_SZW-1:0]  a_size;
      logic  [top_pkg::TL_AIW-1:0]  a_source;
      logic   [top_pkg::TL_AW-1:0]  a_address;
      logic  [top_pkg::TL_DBW-1:0]  a_mask;
      logic   [top_pkg::TL_DW-1:0]  a_data;
      tl_a_user_t                   a_user;
    } tl_txn_data_t;

    tl_txn_data_t txn_data;
    tl_txn_data_t held_data;
    logic fifo_rdy;
    localparam int TxnDataWidth = $bits(tl_txn_data_t);

    assign txn_data = '{
      a_param: tl_i.a_param,
      a_size: tl_i.a_size,
      a_source: tl_i.a_source,
      a_address: tl_i.a_address,
      a_mask: tl_i.a_mask,
      a_data: tl_i.a_data,
      a_user: tl_i.a_user
    };

    prim_fifo_sync #(
      .Width(TxnDataWidth),
      .Pass(1'b0),
      .Depth(1),
      .OutputZeroIfEmpty(1'b0)
    ) u_sync_fifo (
      .clk_i,
      .rst_ni,
      .clr_i(1'b0),
      .wvalid_i(byte_req_ack),
      .wready_o(fifo_rdy),
      .wdata_i(txn_data),
      .rvalid_o(),
      .rready_i(sram_a_ack),
      .rdata_o(held_data),
      .full_o(),
      .depth_o(),
      .err_o()
    );

    // captured read data
    logic [top_pkg::TL_DW-1:0] rsp_data;
    always_ff @(posedge clk_i) begin
      if (sram_d_ack && rd_wait) begin
        rsp_data <= tl_sram_i.d_data;
      end
    end

    // while we could simply not assert a_ready to ensure the host keeps
    // the request lines stable, there is no guarantee the hosts (if there are multiple)
    // do not re-arbitrate on every cycle if its transactions are not accepted.
    // As a result, it is better to capture the transaction attributes.
    logic [top_pkg::TL_DW-1:0] combined_data, unused_data;
    always_comb begin
      for (int i = 0; i < top_pkg::TL_DBW; i++) begin
        combined_data[i*8 +: 8] = held_data.a_mask[i] ?
                                  held_data.a_data[i*8 +: 8] :
                                  rsp_data[i*8 +: 8];
      end
    end

    // Compute updated integrity bits for the data.
    // Note that the CMD integrity does not have to be correct, since it is not consumed nor
    // checked further downstream.
    logic [tlul_pkg::DataIntgWidth-1:0] data_intg;

    tlul_data_integ_enc u_tlul_data_integ_enc (
      .data_i(combined_data),
      .data_intg_o({data_intg, unused_data})
    );

    tl_a_user_t combined_user;
    always_comb begin
      combined_user           = held_data.a_user;
      combined_user.data_intg = data_intg;
    end

    localparam int unsigned AccessSize = $clog2(top_pkg::TL_DBW);
    always_comb begin
      // Pass-through by default
      tl_sram_o = tl_i;
      // if we're waiting for an internal read for RMW, we force this to 1.
      tl_sram_o.d_ready = tl_i.d_ready | rd_wait;

      // We take over the TL-UL bus if there is a pending read or write for the RMW transaction.
      // TL-UL signals are selectively muxed below to reduce complexity and remove long timing
      // paths through the error_i signal. In particular, we avoid creating paths from error_i
      // to the address and data output since these may feed into RAM scrambling logic further
      // downstream.

      // Write transactions for RMW.
      if (wr_phase) begin
        tl_sram_o.a_valid   = 1'b1;
        tl_sram_o.a_opcode  = PutFullData;
        // Since we are performing a read-modify-write operation,
        // we always access the entire word.
        tl_sram_o.a_size    = top_pkg::TL_SZW'(AccessSize);
        tl_sram_o.a_mask    = '{default: '1};
        // override with held / combined data.
        // need to use word aligned addresses here.
        tl_sram_o.a_address = held_data.a_address;
        tl_sram_o.a_address[AccessSize-1:0] = '0;
        tl_sram_o.a_source  = held_data.a_source;
        tl_sram_o.a_param   = held_data.a_param;
        tl_sram_o.a_data    = combined_data;
        tl_sram_o.a_user    = combined_user;
      // Read transactions for RMW.
      end else if (rd_phase) begin
        // need to use word aligned addresses here.
        tl_sram_o.a_address[AccessSize-1:0] = '0;
        // Only override the control signals if there is no error at the input.
        if (!error_i || stall_host) begin
          // Since we are performing a read-modify-write operation,
          // we always access the entire word.
          tl_sram_o.a_size    = top_pkg::TL_SZW'(AccessSize);
          tl_sram_o.a_mask    = '{default: '1};
          // use incoming valid as long as we are not stalling the host
          tl_sram_o.a_valid   = tl_i.a_valid & ~stall_host;
          tl_sram_o.a_opcode  = Get;
        end
      end
    end

    // This assert is necessary for the casting of AccessSize.
    `ASSERT(TlulSramByteTlSize_A, top_pkg::TL_SZW >= $clog2(AccessSize + 1))

    logic unused_held_data;
    assign unused_held_data = ^{held_data.a_address[AccessSize-1:0],
                                held_data.a_user.data_intg,
                                held_data.a_size};

    assign error_o = error_i & ~stall_host;

    logic size_fifo_rdy;
    logic [top_pkg::TL_SZW-1:0] a_size;
    prim_fifo_sync #(
      .Width(top_pkg::TL_SZW),
      .Pass(1'b0),
      .Depth(Outstanding),
      .OutputZeroIfEmpty(1'b1)
    ) u_sync_fifo_a_size (
      .clk_i,
      .rst_ni,
      .clr_i(1'b0),
      .wvalid_i(a_ack),
      .wready_o(size_fifo_rdy),
      .wdata_i(tl_i.a_size),
      .rvalid_o(),
      .rready_i(d_ack),
      .rdata_o(a_size),
      .full_o(),
      .depth_o(pending_txn_cnt),
      .err_o()
    );

    always_comb begin
      tl_o = tl_sram_i;

      // pass a_ready through directly if we are not stalling
      tl_o.a_ready = tl_sram_i.a_ready & ~stall_host & fifo_rdy & size_fifo_rdy;

      // when internal logic has taken over, do not show response to host during
      // read phase.  During write phase, allow the host to see the completion.
      tl_o.d_valid = tl_sram_i.d_valid & ~rd_wait;

      // the size returned by tl_sram_i does not always correspond to the actual
      // transaction size in cases where a read modify write operation is
      // performed. Hence, we always return the registered size here.
      tl_o.d_size  = a_size;
    end // always_comb

    // unused info from tl_sram_i
    // see explanation in above block
    logic unused_tl;
    assign unused_tl = |tl_sram_i.d_size;

    // when byte access detected, go to wait read
    `ASSERT(ByteAccessStateChange_A, a_ack & wr_txn & ~&tl_i.a_mask & ~error_i |=>
      state_q inside {StWaitRd})
    // when in wait for read, a successful response should move to write phase
    `ASSERT(ReadCompleteStateChange_A,
        (state_q == StWaitRd) && (pending_txn_cnt == 1) && sram_d_ack |=> state_q == StWriteCmd)

  end else begin : gen_no_integ_handling
    // In this case we pass everything just through.
    assign tl_sram_o = tl_i;
    assign tl_o = tl_sram_i;
    assign error_o = error_i;
  end

endmodule // tlul_adapter_sram


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL adapter for SRAM-like devices
 *
 * This module handles byte writes for tlul integrity.
 * When a byte write is received, the downstream data is read first
 * to correctly create the integrity constant.
 *
 * A tlul transaction goes through this module.  If required, a
 * tlul read transaction is generated out first.  If not required, the
 * incoming tlul transaction is directly muxed out.
 */
module tlul_sram_byte64 import tlul_pkg::*; #(
  parameter bit EnableIntg  = 0,  // Enable integrity handling at byte level
  parameter int Outstanding = 1
) (
  input clk_i,
  input rst_ni,

  input tl_h2d_t64 tl_i,
  output tl_d2h_t64 tl_o,

  output tl_h2d_t64 tl_sram_o,
  input tl_d2h_t64 tl_sram_i,

  // if incoming transaction already has an error, do not
  // attempt to handle the byte-write access.  Instead treat as
  // feedthrough and allow the system to directly error back.
  // The error indication is also fed through
  input error_i,
  output logic error_o
);

  if (EnableIntg) begin : gen_integ_handling

    // state enumeration
    typedef enum logic [1:0] {
      StPassThru,
      StWaitRd,
      StWriteCmd
    } state_e;

    // state and selection
    logic stall_host;
    logic rd_phase;
    logic rd_wait;
    logic wr_phase;
    state_e state_d, state_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        state_q <= StPassThru;
      end else begin
        state_q <= state_d;
      end
    end

    // transaction qualifying signals
    logic a_ack;  // upstream a channel acknowledgement
    logic d_ack;  // upstream d channel acknowledgement
    logic sram_a_ack; // downstream a channel acknowledgement
    logic sram_d_ack; // downstream d channel acknowledgement
    logic wr_txn;
    logic byte_wr_txn;
    logic byte_req_ack;
    logic [prim_util_pkg::vbits(Outstanding+1)-1:0] pending_txn_cnt;

    assign a_ack = tl_i.a_valid & tl_o.a_ready;
    assign d_ack = tl_o.d_valid & tl_i.d_ready;
    assign sram_a_ack = tl_sram_o.a_valid & tl_sram_i.a_ready;
    assign sram_d_ack = tl_sram_i.d_valid & tl_sram_o.d_ready;
    assign wr_txn = (tl_i.a_opcode == PutFullData) | (tl_i.a_opcode == PutPartialData);

    assign byte_req_ack = byte_wr_txn & a_ack & ~error_i;
    assign byte_wr_txn = tl_i.a_valid & ~&tl_i.a_mask & wr_txn;

    // state machine handling
    always_comb begin
      rd_wait = 1'b0;
      stall_host = 1'b0;
      wr_phase = 1'b0;
      rd_phase = 1'b0;
      state_d = state_q;

      unique case (state_q)
        StPassThru: begin
          if (byte_wr_txn) begin
            rd_phase = 1'b1;
            if (byte_req_ack) begin
              state_d = StWaitRd;
            end
          end
        end

        // Due to the way things are serialized, there is no way for the logic to tell which read
        // belongs to the partial read unless it flushes all prior transactions. Hence, we wait
        // here until exactly one outstanding transaction remains (that one is the partial read).
        StWaitRd: begin
          rd_phase = 1'b1;
          stall_host = 1'b1;
          if (pending_txn_cnt == $bits(pending_txn_cnt)'(1)) begin
            rd_wait = 1'b1;
            if (sram_d_ack) begin
              state_d = StWriteCmd;
            end
          end
        end

        StWriteCmd: begin
          stall_host = 1'b1;
          wr_phase = 1'b1;

          if (sram_a_ack) begin
            state_d = StPassThru;
          end
        end

        default:;

      endcase // unique case (state_q)

    end

    // prim fifo for capturing info
    typedef struct packed {
      logic                  [2:0]  a_param;
      logic  [top_pkg::TL_SZW64-1:0]  a_size;
      logic  [top_pkg::TL_AIW-1:0]  a_source;
      logic   [top_pkg::TL_AW-1:0]  a_address;
      logic  [top_pkg::TL_DBW64-1:0]  a_mask;
      logic   [top_pkg::TL_DW64-1:0]  a_data;
      tl_a_user_t                   a_user;
    } tl_txn_data_t;

    tl_txn_data_t txn_data;
    tl_txn_data_t held_data;
    logic fifo_rdy;
    localparam int TxnDataWidth = $bits(tl_txn_data_t);

    assign txn_data = '{
      a_param: tl_i.a_param,
      a_size: tl_i.a_size,
      a_source: tl_i.a_source,
      a_address: tl_i.a_address,
      a_mask: tl_i.a_mask,
      a_data: tl_i.a_data,
      a_user: tl_i.a_user
    };

    prim_fifo_sync #(
      .Width(TxnDataWidth),
      .Pass(1'b0),
      .Depth(1),
      .OutputZeroIfEmpty(1'b0)
    ) u_sync_fifo (
      .clk_i,
      .rst_ni,
      .clr_i(1'b0),
      .wvalid_i(byte_req_ack),
      .wready_o(fifo_rdy),
      .wdata_i(txn_data),
      .rvalid_o(),
      .rready_i(sram_a_ack),
      .rdata_o(held_data),
      .full_o(),
      .depth_o(),
      .err_o()
    );

    // captured read data
    logic [top_pkg::TL_DW64-1:0] rsp_data;
    always_ff @(posedge clk_i) begin
      if (sram_d_ack && rd_wait) begin
        rsp_data <= tl_sram_i.d_data;
      end
    end

    // while we could simply not assert a_ready to ensure the host keeps
    // the request lines stable, there is no guarantee the hosts (if there are multiple)
    // do not re-arbitrate on every cycle if its transactions are not accepted.
    // As a result, it is better to capture the transaction attributes.
    logic [top_pkg::TL_DW64-1:0] combined_data, unused_data;
    always_comb begin
      for (int i = 0; i < top_pkg::TL_DBW64; i++) begin
        combined_data[i*8 +: 8] = held_data.a_mask[i] ?
                                  held_data.a_data[i*8 +: 8] :
                                  rsp_data[i*8 +: 8];
      end
    end

    // Compute updated integrity bits for the data.
    // Note that the CMD integrity does not have to be correct, since it is not consumed nor
    // checked further downstream.
    logic [tlul_pkg::DataIntgWidth-1:0] data_intg;

    tlul_data_integ_enc u_tlul_data_integ_enc (
      .data_i(combined_data),
      .data_intg_o({data_intg, unused_data})
    );

    tl_a_user_t combined_user;
    always_comb begin
      combined_user           = held_data.a_user;
      combined_user.data_intg = data_intg;
    end

    localparam int unsigned AccessSize = $clog2(top_pkg::TL_DBW64);
    always_comb begin
      // Pass-through by default
      tl_sram_o = tl_i;
      // if we're waiting for an internal read for RMW, we force this to 1.
      tl_sram_o.d_ready = tl_i.d_ready | rd_wait;

      // We take over the TL-UL bus if there is a pending read or write for the RMW transaction.
      // TL-UL signals are selectively muxed below to reduce complexity and remove long timing
      // paths through the error_i signal. In particular, we avoid creating paths from error_i
      // to the address and data output since these may feed into RAM scrambling logic further
      // downstream.

      // Write transactions for RMW.
      if (wr_phase) begin
        tl_sram_o.a_valid   = 1'b1;
        tl_sram_o.a_opcode  = PutFullData;
        // Since we are performing a read-modify-write operation,
        // we always access the entire word.
        tl_sram_o.a_size    = top_pkg::TL_SZW64'(AccessSize);
        tl_sram_o.a_mask    = '{default: '1};
        // override with held / combined data.
        // need to use word aligned addresses here.
        tl_sram_o.a_address = held_data.a_address;
        tl_sram_o.a_address[AccessSize-1:0] = '0;
        tl_sram_o.a_source  = held_data.a_source;
        tl_sram_o.a_param   = held_data.a_param;
        tl_sram_o.a_data    = combined_data;
        tl_sram_o.a_user    = combined_user;
      // Read transactions for RMW.
      end else if (rd_phase) begin
        // need to use word aligned addresses here.
        tl_sram_o.a_address[AccessSize-1:0] = '0;
        // Only override the control signals if there is no error at the input.
        if (!error_i || stall_host) begin
          // Since we are performing a read-modify-write operation,
          // we always access the entire word.
          tl_sram_o.a_size    = top_pkg::TL_SZW64'(AccessSize);
          tl_sram_o.a_mask    = '{default: '1};
          // use incoming valid as long as we are not stalling the host
          tl_sram_o.a_valid   = tl_i.a_valid & ~stall_host;
          tl_sram_o.a_opcode  = Get;
        end
      end
    end

    // This assert is necessary for the casting of AccessSize.
    `ASSERT(TlulSramByteTlSize_A, top_pkg::TL_SZW64 >= $clog2(AccessSize + 1))

    logic unused_held_data;
    assign unused_held_data = ^{held_data.a_address[AccessSize-1:0],
                                held_data.a_user.data_intg,
                                held_data.a_size};

    assign error_o = error_i & ~stall_host;

    logic size_fifo_rdy;
    logic [top_pkg::TL_SZW64-1:0] a_size;
    prim_fifo_sync #(
      .Width(top_pkg::TL_SZW64),
      .Pass(1'b0),
      .Depth(Outstanding),
      .OutputZeroIfEmpty(1'b1)
    ) u_sync_fifo_a_size (
      .clk_i,
      .rst_ni,
      .clr_i(1'b0),
      .wvalid_i(a_ack),
      .wready_o(size_fifo_rdy),
      .wdata_i(tl_i.a_size),
      .rvalid_o(),
      .rready_i(d_ack),
      .rdata_o(a_size),
      .full_o(),
      .depth_o(pending_txn_cnt),
      .err_o()
    );

    always_comb begin
      tl_o = tl_sram_i;

      // pass a_ready through directly if we are not stalling
      tl_o.a_ready = tl_sram_i.a_ready & ~stall_host & fifo_rdy & size_fifo_rdy;

      // when internal logic has taken over, do not show response to host during
      // read phase.  During write phase, allow the host to see the completion.
      tl_o.d_valid = tl_sram_i.d_valid & ~rd_wait;

      // the size returned by tl_sram_i does not always correspond to the actual
      // transaction size in cases where a read modify write operation is
      // performed. Hence, we always return the registered size here.
      tl_o.d_size  = a_size;
    end // always_comb

    // unused info from tl_sram_i
    // see explanation in above block
    logic unused_tl;
    assign unused_tl = |tl_sram_i.d_size;

    // when byte access detected, go to wait read
    `ASSERT(ByteAccessStateChange_A, a_ack & wr_txn & ~&tl_i.a_mask & ~error_i |=>
      state_q inside {StWaitRd})
    // when in wait for read, a successful response should move to write phase
    `ASSERT(ReadCompleteStateChange_A,
        (state_q == StWaitRd) && (pending_txn_cnt == 1) && sram_d_ack |=> state_q == StWriteCmd)

  end else begin : gen_no_integ_handling
    // In this case we pass everything just through.
    assign tl_sram_o = tl_i;
    assign tl_o = tl_sram_i;
    assign error_o = error_i;
  end

endmodule // tlul_adapter_sram


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL adapter for SRAM-like devices
 *
 * - Intentionally omitted BaseAddr in case of multiple memory maps are used in a SoC,
 *   it means that aliasing can happen if target device size in TL-UL crossbar is bigger
 *   than SRAM size
 * - At most one of EnableDataIntgGen / EnableDataIntgPt can be enabled. However it
 *   possible for both to be disabled.
 *   A module can neither generate an integrity response nor pass through any pre-existing
 *   integrity.  This might be the case for non-security critical memories where there is
 *   no stored integrity AND another entity upstream is already generating returning integrity.
 *   There is however no case where EnableDataIntgGen and EnableDataIntgPt are both true.
 */
module tlul_adapter_sram
  import tlul_pkg::*;
  import prim_mubi_pkg::mubi4_t;
#(
  parameter int SramAw            = 12,
  parameter int SramDw            = 32, // Must be multiple of the TL width
  parameter int Outstanding       = 1,  // Only one request is accepted
  parameter bit ByteAccess        = 1,  // 1: Enables sub-word write transactions. Note that this
                                        //    results in read-modify-write operations for integrity
                                        //    re-generation if EnableDataIntgPt is set to 1.
  parameter bit ErrOnWrite        = 0,  // 1: Writes not allowed, automatically error
  parameter bit ErrOnRead         = 0,  // 1: Reads not allowed, automatically error
  parameter bit CmdIntgCheck      = 0,  // 1: Enable command integrity check
  parameter bit EnableRspIntgGen  = 0,  // 1: Generate response integrity
  parameter bit EnableDataIntgGen = 0,  // 1: Generate response data integrity
  parameter bit EnableDataIntgPt  = 0,  // 1: Passthrough command/response data integrity
  parameter bit SecFifoPtr        = 0,  // 1: Duplicated fifo pointers
  localparam int WidthMult        = SramDw / top_pkg::TL_DW,
  localparam int IntgWidth        = tlul_pkg::DataIntgWidth * WidthMult,
  localparam int DataOutW         = EnableDataIntgPt ? SramDw + IntgWidth : SramDw
) (
  input   clk_i,
  input   rst_ni,

  // TL-UL interface
  input   tl_h2d_t          tl_i,
  output  tl_d2h_t          tl_o,

  // control interface
  input   mubi4_t en_ifetch_i,

  // SRAM interface
  output logic                req_o,
  output mubi4_t              req_type_o,
  input                       gnt_i,
  output logic                we_o,
  output logic [SramAw-1:0]   addr_o,
  output logic [DataOutW-1:0] wdata_o,
  output logic [DataOutW-1:0] wmask_o,
  output logic                intg_error_o,
  input        [DataOutW-1:0] rdata_i,
  input                       rvalid_i,
  input        [1:0]          rerror_i // 2 bit error [1]: Uncorrectable, [0]: Correctable
);

  localparam int SramByte = SramDw/8;
  localparam int DataBitWidth = prim_util_pkg::vbits(SramByte);
  localparam int WoffsetWidth = (SramByte == top_pkg::TL_DBW) ? 1 :
                                DataBitWidth - prim_util_pkg::vbits(top_pkg::TL_DBW);

  logic error_det; // Internal protocol error checker
  logic error_internal; // Internal protocol error checker
  logic wr_attr_error;
  logic instr_error;
  logic wr_vld_error;
  logic rd_vld_error;
  logic rsp_fifo_error;
  logic intg_error;
  logic tlul_error;

  // integrity check
  if (CmdIntgCheck) begin : gen_cmd_intg_check
    tlul_cmd_intg_chk u_cmd_intg_chk (
      .tl_i(tl_i),
      .err_o (intg_error)
    );
  end else begin : gen_no_cmd_intg_check
    assign intg_error = '0;
  end

  // permanently latch integrity error until reset
  logic intg_error_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      intg_error_q <= '0;
    end else if (intg_error || rsp_fifo_error) begin
      intg_error_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // or other downstream effects
  assign intg_error_o = intg_error | rsp_fifo_error | intg_error_q;

  // wr_attr_error: Check if the request size, mask are permitted.
  //    Basic check of size, mask, addr align is done in tlul_err module.
  //    Here it checks any partial write if ByteAccess isn't allowed.
  assign wr_attr_error = (tl_i.a_opcode == PutFullData || tl_i.a_opcode == PutPartialData)
                         ? ((ByteAccess == 0) ?
                           (tl_i.a_mask != '1 || tl_i.a_size != 2'h2) : 1'b0)
                           : 1'b0;

  // An instruction type transaction is only valid if en_ifetch is enabled
  // If the instruction type is completely invalid, also considered an instruction error
  assign instr_error = prim_mubi_pkg::mubi4_test_invalid(tl_i.a_user.instr_type) |
                       (prim_mubi_pkg::mubi4_test_true_strict(tl_i.a_user.instr_type) &
                        prim_mubi_pkg::mubi4_test_false_loose(en_ifetch_i));

  if (ErrOnWrite == 1) begin : gen_no_writes
    assign wr_vld_error = tl_i.a_opcode != Get;
  end else begin : gen_writes_allowed
    assign wr_vld_error = 1'b0;
  end

  if (ErrOnRead == 1) begin: gen_no_reads
    assign rd_vld_error = tl_i.a_opcode == Get;
  end else begin : gen_reads_allowed
    assign rd_vld_error = 1'b0;
  end

  // tlul protocol check
  tlul_err u_err (
    .clk_i,
    .rst_ni,
    .tl_i(tl_i),
    .err_o (tlul_error)
  );

  // error return is transactional and thus does not used the "latched" intg_err signal
  assign error_det = wr_attr_error | wr_vld_error | rd_vld_error | instr_error |
                     tlul_error    | intg_error;

  // from sram_byte to adapter logic
  tl_h2d_t tl_i_int;
  // from adapter logic to sram_byte
  tl_d2h_t tl_o_int;
  // from sram_byte to rsp_gen
  tl_d2h_t tl_out;

  // not all parts of tl_i_int are used
  logic unused_tl_i_int;
  assign unused_tl_i_int = ^tl_i_int;

  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(EnableRspIntgGen),
    .EnableDataIntgGen(EnableDataIntgGen)
  ) u_rsp_gen (
    .tl_i(tl_out),
    .tl_o
  );

  // byte handling for integrity
  tlul_sram_byte #(
    .EnableIntg(ByteAccess & EnableDataIntgPt & !ErrOnWrite),
    .Outstanding(Outstanding)
  ) u_sram_byte (
    .clk_i,
    .rst_ni,
    .tl_i,
    .tl_o(tl_out),
    .tl_sram_o(tl_i_int),
    .tl_sram_i(tl_o_int),
    .error_i(error_det),
    .error_o(error_internal)
  );

  typedef struct packed {
    logic [top_pkg::TL_DBW-1:0] mask ; // Byte mask within the TL-UL word
    logic [WoffsetWidth-1:0]    woffset ; // Offset of the TL-UL word within the SRAM word
  } sram_req_t ;

  typedef enum logic [1:0] {
    OpWrite,
    OpRead,
    OpUnknown
  } req_op_e ;

  typedef struct packed {
    req_op_e                    op ;
    logic                       error ;
    prim_mubi_pkg::mubi4_t      instr_type;
    logic [top_pkg::TL_SZW-1:0] size ;
    logic [top_pkg::TL_AIW-1:0] source ;
  } req_t ;

  typedef struct packed {
    logic [top_pkg::TL_DW-1:0] data ;
    logic [DataIntgWidth-1:0]  data_intg ;
    logic                      error ;
  } rsp_t ;

  localparam int SramReqFifoWidth = $bits(sram_req_t) ;
  localparam int ReqFifoWidth = $bits(req_t) ;
  localparam int RspFifoWidth = $bits(rsp_t) ;

  // FIFO signal in case OutStand is greater than 1
  // If request is latched, {write, source} is pushed to req fifo.
  // Req fifo is popped when D channel is acknowledged (v & r)
  // D channel valid is asserted if it is write request or rsp fifo not empty if read.
  logic reqfifo_wvalid, reqfifo_wready;
  logic reqfifo_rvalid, reqfifo_rready;
  req_t reqfifo_wdata,  reqfifo_rdata;

  logic sramreqfifo_wvalid, sramreqfifo_wready;
  logic sramreqfifo_rready;
  sram_req_t sramreqfifo_wdata, sramreqfifo_rdata;

  logic rspfifo_wvalid, rspfifo_wready;
  logic rspfifo_rvalid, rspfifo_rready;
  rsp_t rspfifo_wdata,  rspfifo_rdata;

  logic a_ack, d_ack, sram_ack;
  assign a_ack    = tl_i_int.a_valid & tl_o_int.a_ready ;
  assign d_ack    = tl_o_int.d_valid & tl_i_int.d_ready ;
  assign sram_ack = req_o        & gnt_i ;

  // Valid handling
  logic d_valid, d_error;
  always_comb begin
    d_valid = 1'b0;

    if (reqfifo_rvalid) begin
      if (reqfifo_rdata.error) begin
        // Return error response. Assume no request went out to SRAM
        d_valid = 1'b1;
      end else if (reqfifo_rdata.op == OpRead) begin
        d_valid = rspfifo_rvalid;
      end else begin
        // Write without error
        d_valid = 1'b1;
      end
    end else begin
      d_valid = 1'b0;
    end
  end



  always_comb begin
    d_error = 1'b0;

    if (reqfifo_rvalid) begin
      if (reqfifo_rdata.op == OpRead) begin
        d_error = rspfifo_rdata.error | reqfifo_rdata.error;
      end else begin
        d_error = reqfifo_rdata.error;
      end
    end else begin
      d_error = 1'b0;
    end
  end

  logic vld_rd_rsp;
  assign vld_rd_rsp = d_valid & reqfifo_rvalid & rspfifo_rvalid & (reqfifo_rdata.op == OpRead);
  // If the response data is not valid, we set it to an illegal blanking value which is determined
  // by whether the current transaction is an instruction fetch or a regular read operation.
  logic [top_pkg::TL_DW-1:0] error_blanking_data;
  assign error_blanking_data = (prim_mubi_pkg::mubi4_test_true_strict(reqfifo_rdata.instr_type)) ?
                                 DataWhenInstrError :
                                 DataWhenError;

  // Since DataWhenInstrError and DataWhenError can be arbitrary parameters
  // we statically calculate the correct integrity values for these parameters here so that
  // they do not have to be supplied externally.
  logic [top_pkg::TL_DW-1:0] unused_instr, unused_data;
  logic [DataIntgWidth-1:0] error_instr_integ, error_data_integ;
  tlul_data_integ_enc u_tlul_data_integ_enc_instr (
    .data_i(DataMaxWidth'(DataWhenInstrError)),
    .data_intg_o({error_instr_integ, unused_instr})
  );
  tlul_data_integ_enc u_tlul_data_integ_enc_data (
    .data_i(DataMaxWidth'(DataWhenError)),
    .data_intg_o({error_data_integ, unused_data})
  );

  logic [DataIntgWidth-1:0] error_blanking_integ;
  assign error_blanking_integ = (prim_mubi_pkg::mubi4_test_true_strict(reqfifo_rdata.instr_type)) ?
                                 error_instr_integ :
                                 error_data_integ;

  logic [top_pkg::TL_DW-1:0] d_data;
  assign d_data = (vld_rd_rsp & ~d_error) ? rspfifo_rdata.data   // valid read
                                          : error_blanking_data; // write or TL-UL error

  // If this a write response with data fields set to 0, we have to set all ECC bits correctly
  // since we are using an inverted Hsiao code.
  logic [DataIntgWidth-1:0] data_intg;
  assign data_intg = (vld_rd_rsp && reqfifo_rdata.error) ? error_blanking_integ    : // TL-UL error
                     (vld_rd_rsp)                        ? rspfifo_rdata.data_intg : // valid read
                     prim_secded_pkg::SecdedInv3932ZeroEcc;                          // valid write

  assign tl_o_int = '{
      d_valid  : d_valid ,
      d_opcode : (d_valid && reqfifo_rdata.op != OpRead) ? AccessAck : AccessAckData,
      d_param  : '0,
      d_size   : (d_valid) ? reqfifo_rdata.size : '0,
      d_source : (d_valid) ? reqfifo_rdata.source : '0,
      d_sink   : 1'b0,
      d_data   : d_data,
      d_user   : '{default: '0, data_intg: data_intg},
      d_error  : d_valid && d_error,
      a_ready  : (gnt_i | error_internal) & reqfifo_wready & sramreqfifo_wready
  };

  // a_ready depends on the FIFO full condition and grant from SRAM (or SRAM arbiter)
  // assemble response, including read response, write response, and error for unsupported stuff

  // Output to SRAM:
  //    Generate request only when no internal error occurs. If error occurs, the request should be
  //    dropped and returned error response to the host. So, error to be pushed to reqfifo.
  //    In this case, it is assumed the request is granted (may cause ordering issue later?)
  assign req_o      = tl_i_int.a_valid & reqfifo_wready & ~error_internal;
  assign req_type_o = tl_i_int.a_user.instr_type;
  assign we_o       = tl_i_int.a_valid & (tl_i_int.a_opcode inside {PutFullData, PutPartialData});
  assign addr_o     = (tl_i_int.a_valid) ? tl_i_int.a_address[DataBitWidth+:SramAw] : '0;

  // Support SRAMs wider than the TL-UL word width by mapping the parts of the
  // TL-UL address which are more fine-granular than the SRAM width to the
  // SRAM write mask.
  logic [WoffsetWidth-1:0] woffset;
  if (top_pkg::TL_DW != SramDw) begin : gen_wordwidthadapt
    assign woffset = tl_i_int.a_address[DataBitWidth-1:prim_util_pkg::vbits(top_pkg::TL_DBW)];
  end else begin : gen_no_wordwidthadapt
    assign woffset = '0;
  end

  // The size of the data/wmask depends on whether passthrough integrity is enabled.
  // If passthrough integrity is enabled, the data is concatenated with the integrity passed through
  // the user bits.  Otherwise, it is the data only.
  localparam int DataWidth = EnableDataIntgPt ? top_pkg::TL_DW + DataIntgWidth : top_pkg::TL_DW;

  // Final combined wmask / wdata
  logic [WidthMult-1:0][DataWidth-1:0] wmask_combined;
  logic [WidthMult-1:0][DataWidth-1:0] wdata_combined;

  // Original tlul portion
  logic [WidthMult-1:0][top_pkg::TL_DW-1:0] wmask_int;
  logic [WidthMult-1:0][top_pkg::TL_DW-1:0] wdata_int;

  // Integrity portion
  logic [WidthMult-1:0][DataIntgWidth-1:0] wmask_intg;
  logic [WidthMult-1:0][DataIntgWidth-1:0] wdata_intg;

  always_comb begin
    wmask_int = '0;
    wdata_int = '0;

    if (tl_i_int.a_valid) begin
      for (int i = 0 ; i < top_pkg::TL_DW/8 ; i++) begin
        wmask_int[woffset][8*i +: 8] = {8{tl_i_int.a_mask[i]}};
        wdata_int[woffset][8*i +: 8] = (tl_i_int.a_mask[i] && we_o) ? tl_i_int.a_data[8*i+:8] : '0;
      end
    end
  end

  always_comb begin
    wmask_intg  = '0;
    wdata_intg  = '0;

    if (tl_i_int.a_valid) begin
      wmask_intg[woffset] = {DataIntgWidth{1'b1}};
      wdata_intg[woffset] = tl_i_int.a_user.data_intg;
    end
  end

  for (genvar i = 0; i < WidthMult; i++) begin : gen_write_output
    if (EnableDataIntgPt) begin : gen_combined_output
      assign wmask_combined[i] = {wmask_intg[i], wmask_int[i]};
      assign wdata_combined[i] = {wdata_intg[i], wdata_int[i]};
    end else begin : gen_ft_output
      logic unused_w;
      assign wmask_combined[i] = wmask_int[i];
      assign wdata_combined[i] = wdata_int[i];
      assign unused_w = |wmask_intg & |wdata_intg;
    end
  end

  assign wmask_o = wmask_combined;
  assign wdata_o = wdata_combined;

  assign reqfifo_wvalid = a_ack ; // Push to FIFO only when granted
  assign reqfifo_wdata  = '{
    op:     (tl_i_int.a_opcode != Get) ? OpWrite : OpRead, // To return AccessAck for opcode error
    error:  error_internal,
    instr_type: tl_i_int.a_user.instr_type,
    size:   tl_i_int.a_size,
    source: tl_i_int.a_source
  }; // Store the request only. Doesn't have to store data
  assign reqfifo_rready = d_ack ;

  // push together with ReqFIFO, pop upon returning read
  assign sramreqfifo_wdata = '{
    mask    : tl_i_int.a_mask,
    woffset : woffset
  };
  assign sramreqfifo_wvalid = sram_ack & ~we_o;
  assign sramreqfifo_rready = rspfifo_wvalid;

  assign rspfifo_wvalid = rvalid_i & reqfifo_rvalid;

  // Make sure only requested bytes are forwarded
  logic [WidthMult-1:0][DataWidth-1:0] rdata_reshaped;
  logic [DataWidth-1:0] rdata_tlword;

  // This just changes the array format so that the correct word can be selected by indexing.
  assign rdata_reshaped = rdata_i;

  if (EnableDataIntgPt) begin : gen_no_rmask
    always_comb begin
      // If the read mask is set to zero, all read data is zeroed out by the mask.
      // We have to set the ECC bits accordingly since we are using an inverted Hsiao code.
      rdata_tlword = prim_secded_pkg::SecdedInv3932ZeroWord;
      // Otherwise, if at least one mask bit is nonzero, we are passing through the integrity.
      // In that case we need to feed back the entire word since otherwise the integrity
      // will not calculate correctly.
      if (|sramreqfifo_rdata.mask) begin
        // Select correct word.
        rdata_tlword = rdata_reshaped[sramreqfifo_rdata.woffset];
      end
    end
  end else begin : gen_rmask
    logic [DataWidth-1:0] rmask;
    always_comb begin
      rmask = '0;
      for (int i = 0 ; i < top_pkg::TL_DW/8 ; i++) begin
        rmask[8*i +: 8] = {8{sramreqfifo_rdata.mask[i]}};
      end
    end
    // Select correct word and mask it.
    assign rdata_tlword = rdata_reshaped[sramreqfifo_rdata.woffset] & rmask;
  end

  assign rspfifo_wdata  = '{
    data      : rdata_tlword[top_pkg::TL_DW-1:0],
    data_intg : EnableDataIntgPt ? rdata_tlword[DataWidth-1 -: DataIntgWidth] : '0,
    error     : rerror_i[1] // Only care for Uncorrectable error
  };
  assign rspfifo_rready = (reqfifo_rdata.op == OpRead & ~reqfifo_rdata.error)
                        ? reqfifo_rready : 1'b0 ;

  // This module only cares about uncorrectable errors.
  logic unused_rerror;
  assign unused_rerror = rerror_i[0];

  // FIFO instance: REQ, RSP

  // ReqFIFO is to store the Access type to match to the Response data.
  //    For instance, SRAM accepts the write request but doesn't return the
  //    acknowledge. In this case, it may be hard to determine when the D
  //    response for the write data should send out if reads/writes are
  //    interleaved. So, to make it in-order (even TL-UL allows out-of-order
  //    responses), storing the request is necessary. And if the read entry
  //    is write op, it is safe to return the response right away. If it is
  //    read reqeust, then D response is waiting until read data arrives.
  prim_fifo_sync #(
    .Width   (ReqFifoWidth),
    .Pass    (1'b0),
    .Depth   (Outstanding)
  ) u_reqfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),
    .wvalid_i(reqfifo_wvalid),
    .wready_o(reqfifo_wready),
    .wdata_i (reqfifo_wdata),
    .rvalid_o(reqfifo_rvalid),
    .rready_i(reqfifo_rready),
    .rdata_o (reqfifo_rdata),
    .full_o  (),
    .depth_o (),
    .err_o   ()
  );

  // sramreqfifo:
  //    While the ReqFIFO holds the request until it is sent back via TL-UL, the
  //    sramreqfifo only needs to hold the mask and word offset until the read
  //    data returns from memory.
  prim_fifo_sync #(
    .Width   (SramReqFifoWidth),
    .Pass    (1'b0),
    .Depth   (Outstanding)
  ) u_sramreqfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),
    .wvalid_i(sramreqfifo_wvalid),
    .wready_o(sramreqfifo_wready),
    .wdata_i (sramreqfifo_wdata),
    .rvalid_o(),
    .rready_i(sramreqfifo_rready),
    .rdata_o (sramreqfifo_rdata),
    .full_o  (),
    .depth_o (),
    .err_o   ()
  );

  // Rationale having #Outstanding depth in response FIFO.
  //    In normal case, if the host or the crossbar accepts the response data,
  //    response FIFO isn't needed. But if in any case it has a chance to be
  //    back pressured, the response FIFO should store the returned data not to
  //    lose the data from the SRAM interface. Remember, SRAM interface doesn't
  //    have back-pressure signal such as read_ready.
  prim_fifo_sync #(
    .Width   (RspFifoWidth),
    .Pass    (1'b1),
    .Depth   (Outstanding),
    .Secure  (SecFifoPtr)
  ) u_rspfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),
    .wvalid_i(rspfifo_wvalid),
    .wready_o(rspfifo_wready),
    .wdata_i (rspfifo_wdata),
    .rvalid_o(rspfifo_rvalid),
    .rready_i(rspfifo_rready),
    .rdata_o (rspfifo_rdata),
    .full_o  (),
    .depth_o (),
    .err_o   (rsp_fifo_error)
  );

  // below assertion fails when SRAM rvalid is asserted even though ReqFifo is empty
  `ASSERT(rvalidHighReqFifoEmpty, rvalid_i |-> reqfifo_rvalid)

  // below assertion fails when outstanding value is too small (SRAM rvalid is asserted
  // even though the RspFifo is full)
  `ASSERT(rvalidHighWhenRspFifoFull, rvalid_i |-> rspfifo_wready)

  // If both ErrOnWrite and ErrOnRead are set, this block is useless
  `ASSERT_INIT(adapterNoReadOrWrite, (ErrOnWrite & ErrOnRead) == 0)

  `ASSERT_INIT(SramDwHasByteGranularity_A, SramDw % 8 == 0)
  `ASSERT_INIT(SramDwIsMultipleOfTlulWidth_A, SramDw % top_pkg::TL_DW == 0)

  // These parameter options cannot both be true at the same time
  `ASSERT_INIT(DataIntgOptions_A, ~(EnableDataIntgGen & EnableDataIntgPt))

  // make sure outputs are defined
  `ASSERT_KNOWN(TlOutKnown_A,    tl_o.d_valid)
  `ASSERT_KNOWN_IF(TlOutPayloadKnown_A, tl_o, tl_o.d_valid)
  `ASSERT_KNOWN(ReqOutKnown_A,   req_o  )
  `ASSERT_KNOWN(WeOutKnown_A,    we_o   )
  `ASSERT_KNOWN(AddrOutKnown_A,  addr_o )
  `ASSERT_KNOWN(WdataOutKnown_A, wdata_o)
  `ASSERT_KNOWN(WmaskOutKnown_A, wmask_o)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * Tile-Link UL adapter for SRAM-like devices
 *
 * - Intentionally omitted BaseAddr in case of multiple memory maps are used in a SoC,
 *   it means that aliasing can happen if target device size in TL-UL crossbar is bigger
 *   than SRAM size
 * - At most one of EnableDataIntgGen / EnableDataIntgPt can be enabled. However it
 *   possible for both to be disabled.
 *   A module can neither generate an integrity response nor pass through any pre-existing
 *   integrity.  This might be the case for non-security critical memories where there is
 *   no stored integrity AND another entity upstream is already generating returning integrity.
 *   There is however no case where EnableDataIntgGen and EnableDataIntgPt are both true.
 */
module tlul_adapter_sram64
  import tlul_pkg::*;
  import prim_mubi_pkg::mubi4_t;
#(
  parameter int SramAw            = 12,
  parameter int SramDw            = 64, // Must be multiple of the TL width
  parameter int Outstanding       = 1,  // Only one request is accepted
  parameter bit ByteAccess        = 1,  // 1: Enables sub-word write transactions. Note that this
                                        //    results in read-modify-write operations for integrity
                                        //    re-generation if EnableDataIntgPt is set to 1.
  parameter bit ErrOnWrite        = 0,  // 1: Writes not allowed, automatically error
  parameter bit ErrOnRead         = 0,  // 1: Reads not allowed, automatically error
  parameter bit CmdIntgCheck      = 0,  // 1: Enable command integrity check
  parameter bit EnableRspIntgGen  = 0,  // 1: Generate response integrity
  parameter bit EnableDataIntgGen = 0,  // 1: Generate response data integrity
  parameter bit EnableDataIntgPt  = 0,  // 1: Passthrough command/response data integrity
  parameter bit SecFifoPtr        = 0,  // 1: Duplicated fifo pointers
  localparam int WidthMult        = SramDw / top_pkg::TL_DW64,
  localparam int IntgWidth        = tlul_pkg::DataIntgWidth * WidthMult,
  localparam int DataOutW         = EnableDataIntgPt ? SramDw + IntgWidth : SramDw
) (
  input   clk_i,
  input   rst_ni,

  // TL-UL interface
  input   tl_h2d_t64          tl_i,
  output  tl_d2h_t64          tl_o,

  // control interface
  input   mubi4_t en_ifetch_i,

  // SRAM interface
  output logic                req_o,
  output mubi4_t              req_type_o,
  input                       gnt_i,
  output logic                we_o,
  output logic [SramAw-1:0]   addr_o,
  output logic [DataOutW-1:0] wdata_o,
  output logic [DataOutW-1:0] wmask_o,
  output logic                intg_error_o,
  input        [DataOutW-1:0] rdata_i,
  input                       rvalid_i,
  input        [1:0]          rerror_i // 2 bit error [1]: Uncorrectable, [0]: Correctable
);

  localparam int SramByte = SramDw/8;
  localparam int DataBitWidth = prim_util_pkg::vbits(SramByte);
  localparam int WoffsetWidth = (SramByte == top_pkg::TL_DBW64) ? 1 :
                                DataBitWidth - prim_util_pkg::vbits(top_pkg::TL_DBW64);

  logic error_det; // Internal protocol error checker
  logic error_internal; // Internal protocol error checker
  logic wr_attr_error;
  logic instr_error;
  logic wr_vld_error;
  logic rd_vld_error;
  logic rsp_fifo_error;
  logic intg_error;
  logic tlul_error;

  // integrity check
  if (CmdIntgCheck) begin : gen_cmd_intg_check
    tlul_cmd_intg_chk u_cmd_intg_chk (
      .tl_i(tl_i),
      .err_o (intg_error)
    );
  end else begin : gen_no_cmd_intg_check
    assign intg_error = '0;
  end

  // permanently latch integrity error until reset
  logic intg_error_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      intg_error_q <= '0;
    end else if (intg_error || rsp_fifo_error) begin
      intg_error_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // or other downstream effects
  assign intg_error_o = intg_error | rsp_fifo_error | intg_error_q;

  // wr_attr_error: Check if the request size, mask are permitted.
  //    Basic check of size, mask, addr align is done in tlul_err module.
  //    Here it checks any partial write if ByteAccess isn't allowed.
  assign wr_attr_error = (tl_i.a_opcode == PutFullData || tl_i.a_opcode == PutPartialData)
                         ? ((ByteAccess == 0) ?
                           (tl_i.a_mask != '1 || tl_i.a_size != 2'h2) : 1'b0)
                           : 1'b0;

  // An instruction type transaction is only valid if en_ifetch is enabled
  // If the instruction type is completely invalid, also considered an instruction error
  assign instr_error = prim_mubi_pkg::mubi4_test_invalid(tl_i.a_user.instr_type) |
                       (prim_mubi_pkg::mubi4_test_true_strict(tl_i.a_user.instr_type) &
                        prim_mubi_pkg::mubi4_test_false_loose(en_ifetch_i));

  if (ErrOnWrite == 1) begin : gen_no_writes
    assign wr_vld_error = tl_i.a_opcode != Get;
  end else begin : gen_writes_allowed
    assign wr_vld_error = 1'b0;
  end

  if (ErrOnRead == 1) begin: gen_no_reads
    assign rd_vld_error = tl_i.a_opcode == Get;
  end else begin : gen_reads_allowed
    assign rd_vld_error = 1'b0;
  end

  // tlul protocol check
  // tlul_err u_err (
  //   .clk_i,
  //   .rst_ni,
  //   .tl_i(tl_i),
  //   .err_o (tlul_error)
  // );

  //zdr: del tlul err for only support 32bit DW
  logic tlul_error64;
  // assign tlul_error64 = tlul_error? 1'b0 : 1'b0;
  assign tlul_error64 = 1'b0;
  
  // error return is transactional and thus does not used the "latched" intg_err signal
  assign error_det = wr_attr_error | wr_vld_error | rd_vld_error | instr_error |
                     tlul_error64    | intg_error;

  // from sram_byte to adapter logic
  tl_h2d_t64 tl_i_int;
  // from adapter logic to sram_byte
  tl_d2h_t64 tl_o_int;
  // from sram_byte to rsp_gen
  tl_d2h_t64 tl_out;

  // not all parts of tl_i_int are used
  logic unused_tl_i_int;
  assign unused_tl_i_int = ^tl_i_int;

  //zdr: del tlul_rsp_intg_gen
  // tlul_rsp_intg_gen #(
  //   .EnableRspIntgGen(EnableRspIntgGen),
  //   .EnableDataIntgGen(EnableDataIntgGen)
  // ) u_rsp_gen (
  //   .tl_i(tl_out),
  //   .tl_o
  // );
  assign tl_o = tl_out;

  // byte handling for integrity
  tlul_sram_byte64 #(
    .EnableIntg(ByteAccess & EnableDataIntgPt & !ErrOnWrite),
    .Outstanding(Outstanding)
  ) u_sram_byte (
    .clk_i,
    .rst_ni,
    .tl_i,
    .tl_o(tl_out),
    .tl_sram_o(tl_i_int),
    .tl_sram_i(tl_o_int),
    .error_i(error_det),
    .error_o(error_internal)
  );

  typedef struct packed {
    logic [top_pkg::TL_DBW64-1:0] mask ; // Byte mask within the TL-UL word
    logic [WoffsetWidth-1:0]    woffset ; // Offset of the TL-UL word within the SRAM word
  } sram_req_t ;

  typedef enum logic [1:0] {
    OpWrite,
    OpRead,
    OpUnknown
  } req_op_e ;

  typedef struct packed {
    req_op_e                    op ;
    logic                       error ;
    prim_mubi_pkg::mubi4_t      instr_type;
    logic [top_pkg::TL_SZW64-1:0] size ;
    logic [top_pkg::TL_AIW-1:0] source ;
  } req_t ;

  typedef struct packed {
    logic [top_pkg::TL_DW64-1:0] data ;
    logic [DataIntgWidth-1:0]  data_intg ;
    logic                      error ;
  } rsp_t ;

  localparam int SramReqFifoWidth = $bits(sram_req_t) ;
  localparam int ReqFifoWidth = $bits(req_t) ;
  localparam int RspFifoWidth = $bits(rsp_t) ;

  // FIFO signal in case OutStand is greater than 1
  // If request is latched, {write, source} is pushed to req fifo.
  // Req fifo is popped when D channel is acknowledged (v & r)
  // D channel valid is asserted if it is write request or rsp fifo not empty if read.
  logic reqfifo_wvalid, reqfifo_wready;
  logic reqfifo_rvalid, reqfifo_rready;
  req_t reqfifo_wdata,  reqfifo_rdata;

  logic sramreqfifo_wvalid, sramreqfifo_wready;
  logic sramreqfifo_rready;
  sram_req_t sramreqfifo_wdata, sramreqfifo_rdata;

  logic rspfifo_wvalid, rspfifo_wready;
  logic rspfifo_rvalid, rspfifo_rready;
  rsp_t rspfifo_wdata,  rspfifo_rdata;

  logic a_ack, d_ack, sram_ack;
  assign a_ack    = tl_i_int.a_valid & tl_o_int.a_ready ;
  assign d_ack    = tl_o_int.d_valid & tl_i_int.d_ready ;
  assign sram_ack = req_o        & gnt_i ;

  // Valid handling
  logic d_valid, d_error;
  always_comb begin
    d_valid = 1'b0;

    if (reqfifo_rvalid) begin
      if (reqfifo_rdata.error) begin
        // Return error response. Assume no request went out to SRAM
        d_valid = 1'b1;
      end else if (reqfifo_rdata.op == OpRead) begin
        d_valid = rspfifo_rvalid;
      end else begin
        // Write without error
        d_valid = 1'b1;
      end
    end else begin
      d_valid = 1'b0;
    end
  end



  always_comb begin
    d_error = 1'b0;

    if (reqfifo_rvalid) begin
      if (reqfifo_rdata.op == OpRead) begin
        d_error = rspfifo_rdata.error | reqfifo_rdata.error;
      end else begin
        d_error = reqfifo_rdata.error;
      end
    end else begin
      d_error = 1'b0;
    end
  end

  logic vld_rd_rsp;
  assign vld_rd_rsp = d_valid & reqfifo_rvalid & rspfifo_rvalid & (reqfifo_rdata.op == OpRead);
  // If the response data is not valid, we set it to an illegal blanking value which is determined
  // by whether the current transaction is an instruction fetch or a regular read operation.
  logic [top_pkg::TL_DW64-1:0] error_blanking_data;
  assign error_blanking_data = (prim_mubi_pkg::mubi4_test_true_strict(reqfifo_rdata.instr_type)) ?
                                 DataWhenInstrError :
                                 DataWhenError;

  // Since DataWhenInstrError and DataWhenError can be arbitrary parameters
  // we statically calculate the correct integrity values for these parameters here so that
  // they do not have to be supplied externally.
  logic [top_pkg::TL_DW64-1:0] unused_instr, unused_data;
  // logic [DataIntgWidth-1:0] error_instr_integ, error_data_integ;
  // tlul_data_integ_enc u_tlul_data_integ_enc_instr (
  //   .data_i(DataMaxWidth'(DataWhenInstrError)),
  //   .data_intg_o({error_instr_integ, unused_instr})
  // );
  // tlul_data_integ_enc u_tlul_data_integ_enc_data (
  //   .data_i(DataMaxWidth'(DataWhenError)),
  //   .data_intg_o({error_data_integ, unused_data})
  // );
  logic [DataIntgWidth-1:0] error_instr_integ = '0;
  logic [DataIntgWidth-1:0]  error_data_integ = '0;

  logic [DataIntgWidth-1:0] error_blanking_integ = '0;
  // assign error_blanking_integ = (prim_mubi_pkg::mubi4_test_true_strict(reqfifo_rdata.instr_type)) ?
  //                                error_instr_integ :
  //                                error_data_integ;

  logic [top_pkg::TL_DW64-1:0] d_data;
  assign d_data = (vld_rd_rsp & ~d_error) ? rspfifo_rdata.data   // valid read
                                          : error_blanking_data; // write or TL-UL error

  // If this a write response with data fields set to 0, we have to set all ECC bits correctly
  // since we are using an inverted Hsiao code.
  logic [DataIntgWidth-1:0] data_intg;
  assign data_intg = (vld_rd_rsp && reqfifo_rdata.error) ? '0    : // TL-UL error
                     (vld_rd_rsp)                        ? rspfifo_rdata.data_intg : // valid read
                     prim_secded_pkg::SecdedInv3932ZeroEcc;                          // valid write

  assign tl_o_int = '{
      d_valid  : d_valid ,
      d_opcode : (d_valid && reqfifo_rdata.op != OpRead) ? AccessAck : AccessAckData,
      d_param  : '0,
      d_size   : (d_valid) ? reqfifo_rdata.size : '0,
      d_source : (d_valid) ? reqfifo_rdata.source : '0,
      d_sink   : 1'b0,
      d_data   : d_data,
      d_user   : '{default: '0, data_intg: data_intg},
      d_error  : d_valid && d_error,
      a_ready  : (gnt_i | error_internal) & reqfifo_wready & sramreqfifo_wready
  };

  // a_ready depends on the FIFO full condition and grant from SRAM (or SRAM arbiter)
  // assemble response, including read response, write response, and error for unsupported stuff

  // Output to SRAM:
  //    Generate request only when no internal error occurs. If error occurs, the request should be
  //    dropped and returned error response to the host. So, error to be pushed to reqfifo.
  //    In this case, it is assumed the request is granted (may cause ordering issue later?)
  assign req_o      = tl_i_int.a_valid & reqfifo_wready & ~error_internal;
  assign req_type_o = tl_i_int.a_user.instr_type;
  assign we_o       = tl_i_int.a_valid & (tl_i_int.a_opcode inside {PutFullData, PutPartialData});
  //zdr: addr gen change
  assign addr_o     = (tl_i_int.a_valid) ? tl_i_int.a_address[DataBitWidth+:SramAw] : '0;

  // Support SRAMs wider than the TL-UL word width by mapping the parts of the
  // TL-UL address which are more fine-granular than the SRAM width to the
  // SRAM write mask.
  logic [WoffsetWidth-1:0] woffset;
  if (top_pkg::TL_DW64 != SramDw) begin : gen_wordwidthadapt
    assign woffset = tl_i_int.a_address[DataBitWidth-1:prim_util_pkg::vbits(top_pkg::TL_DBW64)];
  end else begin : gen_no_wordwidthadapt
    assign woffset = '0;
  end

  // The size of the data/wmask depends on whether passthrough integrity is enabled.
  // If passthrough integrity is enabled, the data is concatenated with the integrity passed through
  // the user bits.  Otherwise, it is the data only.
  localparam int DataWidth = EnableDataIntgPt ? top_pkg::TL_DW64 + DataIntgWidth : top_pkg::TL_DW64;

  // Final combined wmask / wdata
  logic [WidthMult-1:0][DataWidth-1:0] wmask_combined;
  logic [WidthMult-1:0][DataWidth-1:0] wdata_combined;

  // Original tlul portion
  logic [WidthMult-1:0][top_pkg::TL_DW64-1:0] wmask_int;
  logic [WidthMult-1:0][top_pkg::TL_DW64-1:0] wdata_int;

  // Integrity portion
  logic [WidthMult-1:0][DataIntgWidth-1:0] wmask_intg;
  logic [WidthMult-1:0][DataIntgWidth-1:0] wdata_intg;

  always_comb begin
    wmask_int = '0;
    wdata_int = '0;

    if (tl_i_int.a_valid) begin
      for (int i = 0 ; i < top_pkg::TL_DW64/8 ; i++) begin
        wmask_int[woffset][8*i +: 8] = {8{tl_i_int.a_mask[i]}};
        wdata_int[woffset][8*i +: 8] = (tl_i_int.a_mask[i] && we_o) ? tl_i_int.a_data[8*i+:8] : '0;
      end
    end
  end

  always_comb begin
    wmask_intg  = '0;
    wdata_intg  = '0;

    if (tl_i_int.a_valid) begin
      wmask_intg[woffset] = {DataIntgWidth{1'b1}};
      wdata_intg[woffset] = tl_i_int.a_user.data_intg;
    end
  end

  for (genvar i = 0; i < WidthMult; i++) begin : gen_write_output
    if (EnableDataIntgPt) begin : gen_combined_output
      assign wmask_combined[i] = {wmask_intg[i], wmask_int[i]};
      assign wdata_combined[i] = {wdata_intg[i], wdata_int[i]};
    end else begin : gen_ft_output
      logic unused_w;
      assign wmask_combined[i] = wmask_int[i];
      assign wdata_combined[i] = wdata_int[i];
      assign unused_w = |wmask_intg & |wdata_intg;
    end
  end

  assign wmask_o = wmask_combined;
  assign wdata_o = wdata_combined;

  assign reqfifo_wvalid = a_ack ; // Push to FIFO only when granted
  assign reqfifo_wdata  = '{
    op:     (tl_i_int.a_opcode != Get) ? OpWrite : OpRead, // To return AccessAck for opcode error
    error:  error_internal,
    instr_type: tl_i_int.a_user.instr_type,
    size:   tl_i_int.a_size,
    source: tl_i_int.a_source
  }; // Store the request only. Doesn't have to store data
  assign reqfifo_rready = d_ack ;

  // push together with ReqFIFO, pop upon returning read
  assign sramreqfifo_wdata = '{
    mask    : tl_i_int.a_mask,
    woffset : woffset
  };
  assign sramreqfifo_wvalid = sram_ack & ~we_o;
  assign sramreqfifo_rready = rspfifo_wvalid;

  assign rspfifo_wvalid = rvalid_i & reqfifo_rvalid;

  // Make sure only requested bytes are forwarded
  logic [WidthMult-1:0][DataWidth-1:0] rdata_reshaped;
  logic [DataWidth-1:0] rdata_tlword;

  // This just changes the array format so that the correct word can be selected by indexing.
  assign rdata_reshaped = rdata_i;

  if (EnableDataIntgPt) begin : gen_no_rmask
    always_comb begin
      // If the read mask is set to zero, all read data is zeroed out by the mask.
      // We have to set the ECC bits accordingly since we are using an inverted Hsiao code.
      rdata_tlword = prim_secded_pkg::SecdedInv3932ZeroWord;
      // Otherwise, if at least one mask bit is nonzero, we are passing through the integrity.
      // In that case we need to feed back the entire word since otherwise the integrity
      // will not calculate correctly.
      if (|sramreqfifo_rdata.mask) begin
        // Select correct word.
        rdata_tlword = rdata_reshaped[sramreqfifo_rdata.woffset];
      end
    end
  end else begin : gen_rmask
    logic [DataWidth-1:0] rmask;
    always_comb begin
      rmask = '0;
      for (int i = 0 ; i < top_pkg::TL_DW64/8 ; i++) begin
        rmask[8*i +: 8] = {8{sramreqfifo_rdata.mask[i]}};
      end
    end
    // Select correct word and mask it.
    assign rdata_tlword = rdata_reshaped[sramreqfifo_rdata.woffset] & rmask;
  end

  assign rspfifo_wdata  = '{
    data      : rdata_tlword[top_pkg::TL_DW64-1:0],
    data_intg : EnableDataIntgPt ? rdata_tlword[DataWidth-1 -: DataIntgWidth] : '0,
    error     : rerror_i[1] // Only care for Uncorrectable error
  };
  assign rspfifo_rready = (reqfifo_rdata.op == OpRead & ~reqfifo_rdata.error)
                        ? reqfifo_rready : 1'b0 ;

  // This module only cares about uncorrectable errors.
  logic unused_rerror;
  assign unused_rerror = rerror_i[0];

  // FIFO instance: REQ, RSP

  // ReqFIFO is to store the Access type to match to the Response data.
  //    For instance, SRAM accepts the write request but doesn't return the
  //    acknowledge. In this case, it may be hard to determine when the D
  //    response for the write data should send out if reads/writes are
  //    interleaved. So, to make it in-order (even TL-UL allows out-of-order
  //    responses), storing the request is necessary. And if the read entry
  //    is write op, it is safe to return the response right away. If it is
  //    read reqeust, then D response is waiting until read data arrives.
  prim_fifo_sync #(
    .Width   (ReqFifoWidth),
    .Pass    (1'b0),
    .Depth   (Outstanding)
  ) u_reqfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),
    .wvalid_i(reqfifo_wvalid),
    .wready_o(reqfifo_wready),
    .wdata_i (reqfifo_wdata),
    .rvalid_o(reqfifo_rvalid),
    .rready_i(reqfifo_rready),
    .rdata_o (reqfifo_rdata),
    .full_o  (),
    .depth_o (),
    .err_o   ()
  );

  // sramreqfifo:
  //    While the ReqFIFO holds the request until it is sent back via TL-UL, the
  //    sramreqfifo only needs to hold the mask and word offset until the read
  //    data returns from memory.
  prim_fifo_sync #(
    .Width   (SramReqFifoWidth),
    .Pass    (1'b0),
    .Depth   (Outstanding)
  ) u_sramreqfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),
    .wvalid_i(sramreqfifo_wvalid),
    .wready_o(sramreqfifo_wready),
    .wdata_i (sramreqfifo_wdata),
    .rvalid_o(),
    .rready_i(sramreqfifo_rready),
    .rdata_o (sramreqfifo_rdata),
    .full_o  (),
    .depth_o (),
    .err_o   ()
  );

  // Rationale having #Outstanding depth in response FIFO.
  //    In normal case, if the host or the crossbar accepts the response data,
  //    response FIFO isn't needed. But if in any case it has a chance to be
  //    back pressured, the response FIFO should store the returned data not to
  //    lose the data from the SRAM interface. Remember, SRAM interface doesn't
  //    have back-pressure signal such as read_ready.
  prim_fifo_sync #(
    .Width   (RspFifoWidth),
    .Pass    (1'b1),
    .Depth   (Outstanding),
    .Secure  (SecFifoPtr)
  ) u_rspfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),
    .wvalid_i(rspfifo_wvalid),
    .wready_o(rspfifo_wready),
    .wdata_i (rspfifo_wdata),
    .rvalid_o(rspfifo_rvalid),
    .rready_i(rspfifo_rready),
    .rdata_o (rspfifo_rdata),
    .full_o  (),
    .depth_o (),
    .err_o   (rsp_fifo_error)
  );

  // below assertion fails when SRAM rvalid is asserted even though ReqFifo is empty
  `ASSERT(rvalidHighReqFifoEmpty, rvalid_i |-> reqfifo_rvalid)

  // below assertion fails when outstanding value is too small (SRAM rvalid is asserted
  // even though the RspFifo is full)
  `ASSERT(rvalidHighWhenRspFifoFull, rvalid_i |-> rspfifo_wready)

  // If both ErrOnWrite and ErrOnRead are set, this block is useless
  `ASSERT_INIT(adapterNoReadOrWrite, (ErrOnWrite & ErrOnRead) == 0)

  `ASSERT_INIT(SramDwHasByteGranularity_A, SramDw % 8 == 0)
  `ASSERT_INIT(SramDwIsMultipleOfTlulWidth_A, SramDw % top_pkg::TL_DW64 == 0)

  // These parameter options cannot both be true at the same time
  `ASSERT_INIT(DataIntgOptions_A, ~(EnableDataIntgGen & EnableDataIntgPt))

  // make sure outputs are defined
  `ASSERT_KNOWN(TlOutKnown_A,    tl_o.d_valid)
  `ASSERT_KNOWN_IF(TlOutPayloadKnown_A, tl_o, tl_o.d_valid)
  `ASSERT_KNOWN(ReqOutKnown_A,   req_o  )
  `ASSERT_KNOWN(WeOutKnown_A,    we_o   )
  `ASSERT_KNOWN(AddrOutKnown_A,  addr_o )
  `ASSERT_KNOWN(WdataOutKnown_A, wdata_o)
  `ASSERT_KNOWN(WmaskOutKnown_A, wmask_o)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Life cycle gating module for TL-UL protocol.
// Transactions are passed through when lc_en_i == ON.
// In all other cases (lc_en_i != ON) incoming transactions return a bus error.
//
// Note that the lc_en_i should be synchronized and buffered outside of this module using
// an instance of prim_lc_sync.

module tlul_lc_gate
  import tlul_pkg::*;
  import lc_ctrl_pkg::*;
#(
  // Number of LC gating muxes in each direction.
  // It is recommended to set this parameter to 2, which results
  // in a total of 4 gating muxes.
  parameter int NumGatesPerDirection = 2
) (
  input clk_i,
  input rst_ni,

  // To host
  input  tl_h2d_t tl_h2d_i,
  output tl_d2h_t tl_d2h_o,

  // To device
  output tl_h2d_t tl_h2d_o,
  input  tl_d2h_t tl_d2h_i,

  // Flush control signaling
  input flush_req_i,
  output logic flush_ack_o,

  // Indicates whether there are pending responses on the device side.
  output logic resp_pending_o,

  // LC control signal
  input  lc_tx_t  lc_en_i,
  output logic err_o
);

  //////////////////
  // Access Gates //
  //////////////////

  lc_tx_t err_en;
  lc_tx_t [NumGatesPerDirection-1:0] err_en_buf;

  prim_lc_sync #(
    .NumCopies(NumGatesPerDirection),
    .AsyncOn(0)
  ) u_err_en_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i(err_en),
    .lc_en_o(err_en_buf)
  );

  tl_h2d_t tl_h2d_int [NumGatesPerDirection+1];
  tl_d2h_t tl_d2h_int [NumGatesPerDirection+1];
  for (genvar k = 0; k < NumGatesPerDirection; k++) begin : gen_lc_gating_muxes
    // H -> D path.
    prim_blanker #(
      .Width($bits(tl_h2d_t))
    ) u_prim_blanker_h2d (
      .in_i(tl_h2d_int[k]),
      .en_i(lc_tx_test_false_strict(err_en_buf[k])),
      .out_o(tl_h2d_int[k+1])
    );

    // D -> H path.
    prim_blanker #(
      .Width($bits(tl_d2h_t))
    ) u_prim_blanker_d2h (
      .in_i(tl_d2h_int[k+1]),
      .en_i(lc_tx_test_false_strict(err_en_buf[k])),
      .out_o(tl_d2h_int[k])
    );
  end

  // Assign signals on the device side.
  assign tl_h2d_o = tl_h2d_int[NumGatesPerDirection];
  assign tl_d2h_int[NumGatesPerDirection] = tl_d2h_i;

  ///////////////////////////
  // Host Side Interposing //
  ///////////////////////////

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 4 -n 8 \
  //      -s 3379253306 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||||||| (66.67%)
  //  6: |||||||||| (33.33%)
  //  7: --
  //  8: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 6
  // Minimum Hamming weight: 3
  // Maximum Hamming weight: 5
  //
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 5 -n 9 \
  //      -s 686407169 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||||||| (60.00%)
  //  6: ||||||||||||| (40.00%)
  //  7: --
  //  8: --
  //  9: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 6
  // Minimum Hamming weight: 3
  // Maximum Hamming weight: 6
  //
  localparam int StateWidth = 9;
  typedef enum logic [StateWidth-1:0] {
    StActive = 9'b100100001,
    StOutstanding = 9'b011100111,
    StFlush = 9'b001001100,
    StError = 9'b010111010,
    StErrorOutstanding = 9'b100010110
  } state_e;

  state_e state_d, state_q;
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, StError)

  logic [1:0] outstanding_txn;
  logic a_ack;
  logic d_ack;
  assign a_ack = tl_h2d_i.a_valid & tl_d2h_o.a_ready;
  assign d_ack = tl_h2d_i.d_ready & tl_d2h_o.d_valid;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      outstanding_txn <= '0;
    end else if (a_ack && !d_ack) begin
      outstanding_txn <= outstanding_txn + 1'b1;
    end else if (d_ack && !a_ack) begin
      outstanding_txn <= outstanding_txn - 1'b1;
    end
  end

  logic block_cmd;
  always_comb begin
    block_cmd = '0;
    state_d = state_q;
    err_en = Off;
    err_o = '0;
    flush_ack_o = '0;
    resp_pending_o = 1'b0;

    unique case (state_q)
      StActive: begin
        if (lc_tx_test_false_loose(lc_en_i) || flush_req_i) begin
          state_d = StOutstanding;
        end
        if (outstanding_txn != '0) begin
          resp_pending_o = 1'b1;
        end
      end

      StOutstanding: begin
        block_cmd = 1'b1;
        if (outstanding_txn == '0) begin
          state_d = lc_tx_test_false_loose(lc_en_i) ? StError : StFlush;
        end else begin
          resp_pending_o = 1'b1;
        end
      end

      StFlush: begin
        block_cmd = 1'b1;
        flush_ack_o = 1'b1;
        if (lc_tx_test_false_loose(lc_en_i)) begin
          state_d = StError;
        end else if (!flush_req_i) begin
          state_d = StActive;
        end
      end

      StError: begin
        err_en = On;
        if (lc_tx_test_true_strict(lc_en_i)) begin
          state_d = StErrorOutstanding;
        end
      end

      StErrorOutstanding: begin
        err_en = On;
        block_cmd = 1'b1;
        if (outstanding_txn == '0) begin
          state_d = StActive;
        end
      end

      default: begin
        err_o = 1'b1;
        err_en = On;
      end

    endcase // unique case (state_q)
  end


  // At the host side, we interpose the ready / valid signals so that we can return a bus error
  // in case the lc signal is not set to ON. Note that this logic does not have to be duplicated
  // since erroring back is considered a convenience feature so that the bus does not lock up.
  tl_h2d_t tl_h2d_error;
  tl_d2h_t tl_d2h_error;
  always_comb begin
    tl_h2d_int[0] = tl_h2d_i;
    tl_d2h_o      = tl_d2h_int[0];
    tl_h2d_error  = '0;

    if (lc_tx_test_true_loose(err_en)) begin
      tl_h2d_error  = tl_h2d_i;
      tl_d2h_o      = tl_d2h_error;
    end

    if (block_cmd) begin
      tl_d2h_o.a_ready = 1'b0;
      tl_h2d_int[0].a_valid = 1'b0;
      tl_h2d_error.a_valid = 1'b0;
    end
  end

  tlul_err_resp u_tlul_err_resp (
    .clk_i,
    .rst_ni,
    .tl_h_i(tl_h2d_error),
    .tl_h_o(tl_d2h_error)
  );

  // Add assertion
  `ASSERT(OutStandingOvfl_A, &outstanding_txn |-> ~a_ack)

endmodule : tlul_lc_gate


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// TL-UL error responder module, used by tlul_socket_1n to help response
// to requests to no correct address space. Responses are always one cycle
// after request with no stalling unless response is stuck on the way out.

module tlul_err_resp (
  input                     clk_i,
  input                     rst_ni,
  input  tlul_pkg::tl_h2d_t tl_h_i,
  output tlul_pkg::tl_d2h_t tl_h_o
);
  import tlul_pkg::*;
  import prim_mubi_pkg::*;

  tl_a_op_e                          err_opcode;
  logic [$bits(tl_h_i.a_source)-1:0] err_source;
  logic [$bits(tl_h_i.a_size)-1:0]   err_size;
  logic                              err_req_pending, err_rsp_pending;
  mubi4_t                            err_instr_type;
  tlul_pkg::tl_d2h_t                 tl_h_o_int;

  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_intg_gen (
    .tl_i(tl_h_o_int),
    .tl_o(tl_h_o)
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_req_pending <= 1'b0;
      err_source      <= {top_pkg::TL_AIW{1'b0}};
      err_opcode      <= Get;
      err_size        <= '0;
      err_instr_type  <= MuBi4False;
    end else if (tl_h_i.a_valid && tl_h_o_int.a_ready) begin
      err_req_pending <= 1'b1;
      err_source      <= tl_h_i.a_source;
      err_opcode      <= tl_h_i.a_opcode;
      err_size        <= tl_h_i.a_size;
      err_instr_type  <= tl_h_i.a_user.instr_type;
    end else if (!err_rsp_pending) begin
      err_req_pending <= 1'b0;
    end
  end

  assign tl_h_o_int.a_ready  = ~err_rsp_pending & ~(err_req_pending & ~tl_h_i.d_ready);
  assign tl_h_o_int.d_valid  = err_req_pending | err_rsp_pending;
  assign tl_h_o_int.d_data   = (mubi4_test_true_strict(err_instr_type)) ? DataWhenInstrError :
                                                                          DataWhenError;
  assign tl_h_o_int.d_source = err_source;
  assign tl_h_o_int.d_sink   = '0;
  assign tl_h_o_int.d_param  = '0;
  assign tl_h_o_int.d_size   = err_size;
  assign tl_h_o_int.d_opcode = (err_opcode == Get) ? AccessAckData : AccessAck;
  assign tl_h_o_int.d_user   = '0;
  assign tl_h_o_int.d_error  = 1'b1;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_rsp_pending <= 1'b0;
    end else if ((err_req_pending || err_rsp_pending) && !tl_h_i.d_ready) begin
      err_rsp_pending <= 1'b1;
    end else begin
      err_rsp_pending <= 1'b0;
    end
  end

  // Waive unused bits of tl_h_i
  logic unused_tl_h;
  assign unused_tl_h = ^tl_h_i;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// TL-UL socket 1:N module
//
// configuration settings
//   device_count: 4
//
// Verilog parameters
//   HReqPass:      if 1 then host requests can pass through on empty fifo,
//                  default 1
//   HRspPass:      if 1 then host responses can pass through on empty fifo,
//                  default 1
//   DReqPass:      (one per device_count) if 1 then device i requests can
//                  pass through on empty fifo, default 1
//   DRspPass:      (one per device_count) if 1 then device i responses can
//                  pass through on empty fifo, default 1
//   HReqDepth:     Depth of host request FIFO, default 2
//   HRspDepth:     Depth of host response FIFO, default 2
//   DReqDepth:     (one per device_count) Depth of device i request FIFO,
//                  default 2
//   DRspDepth:     (one per device_count) Depth of device i response FIFO,
//                  default 2
//   ExplicitErrs:  This module always returns a request error if dev_select_i
//                  is greater than N-1. If ExplicitErrs is set then the width
//                  of the dev_select_i signal will be chosen to make sure that
//                  this is possible. This only makes a difference if N is a
//                  power of 2.
//
// Requests must stall to one device until all responses from other devices
// have returned.  Need to keep a counter of all outstanding requests and
// wait until that counter is zero before switching devices.
//
// This module will return a request error if the input value of 'dev_select_i'
// is not within the range 0..N-1. Thus the instantiator of the socket
// can indicate error by any illegal value of dev_select_i. 4'b1111 is
// recommended for visibility
//
// The maximum value of N is 15

`include "prim_assert.sv"

module tlul_socket_1n #(
  parameter int unsigned  N            = 4,
  parameter bit           HReqPass     = 1'b1,
  parameter bit           HRspPass     = 1'b1,
  parameter bit [N-1:0]   DReqPass     = {N{1'b1}},
  parameter bit [N-1:0]   DRspPass     = {N{1'b1}},
  parameter bit [3:0]     HReqDepth    = 4'h1,
  parameter bit [3:0]     HRspDepth    = 4'h1,
  parameter bit [N*4-1:0] DReqDepth    = {N{4'h1}},
  parameter bit [N*4-1:0] DRspDepth    = {N{4'h1}},
  parameter bit           ExplicitErrs = 1'b1,

  // The width of dev_select_i. We must be able to select any of the N devices
  // (i.e. values 0..N-1). If ExplicitErrs is set, we also need to be able to
  // represent N.
  localparam int unsigned NWD = $clog2(ExplicitErrs ? N+1 : N)
) (
  input                     clk_i,
  input                     rst_ni,
  input  tlul_pkg::tl_h2d_t tl_h_i,
  output tlul_pkg::tl_d2h_t tl_h_o,
  output tlul_pkg::tl_h2d_t tl_d_o    [N],
  input  tlul_pkg::tl_d2h_t tl_d_i    [N],
  input  [NWD-1:0]          dev_select_i
);

  `ASSERT_INIT(maxN, N < 32)

  // Since our steering is done after potential FIFOing, we need to
  // shove our device select bits into spare bits of reqfifo

  // instantiate the host fifo, create intermediate bus 't'

  // FIFO'd version of device select
  logic [NWD-1:0] dev_select_t;

  tlul_pkg::tl_h2d_t   tl_t_o;
  tlul_pkg::tl_d2h_t   tl_t_i;

  tlul_fifo_sync #(
    .ReqPass(HReqPass),
    .RspPass(HRspPass),
    .ReqDepth(HReqDepth),
    .RspDepth(HRspDepth),
    .SpareReqW(NWD)
  ) fifo_h (
    .clk_i,
    .rst_ni,
    .tl_h_i,
    .tl_h_o,
    .tl_d_o     (tl_t_o),
    .tl_d_i     (tl_t_i),
    .spare_req_i (dev_select_i),
    .spare_req_o (dev_select_t),
    .spare_rsp_i (1'b0),
    .spare_rsp_o ());


  // We need to keep track of how many requests are outstanding,
  // and to which device. New requests are compared to this and
  // stall until that number is zero.
  localparam int MaxOutstanding = 2**top_pkg::TL_AIW; // Up to 256 ounstanding
  localparam int OutstandingW = $clog2(MaxOutstanding+1);
  logic [OutstandingW-1:0] num_req_outstanding;
  logic [NWD-1:0]          dev_select_outstanding;
  logic                    hold_all_requests;
  logic                    accept_t_req, accept_t_rsp;

  assign  accept_t_req = tl_t_o.a_valid & tl_t_i.a_ready;
  assign  accept_t_rsp = tl_t_i.d_valid & tl_t_o.d_ready;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      num_req_outstanding <= '0;
      dev_select_outstanding <= '0;
    end else if (accept_t_req) begin
      if (!accept_t_rsp) begin
        `ASSERT_I(NotOverflowed_A, num_req_outstanding <= MaxOutstanding)
        num_req_outstanding <= num_req_outstanding + 1'b1;
      end
      dev_select_outstanding <= dev_select_t;
    end else if (accept_t_rsp) begin
      num_req_outstanding <= num_req_outstanding - 1'b1;
    end
  end

  assign hold_all_requests =
      (num_req_outstanding != '0) &
      (dev_select_t != dev_select_outstanding);

  // Make N copies of 't' request side with modified reqvalid, call
  // them 'u[0]' .. 'u[n-1]'.

  tlul_pkg::tl_h2d_t   tl_u_o [N+1];
  tlul_pkg::tl_d2h_t   tl_u_i [N+1];

  // ensure that when a device is not selected, both command
  // data integrity can never match
  tlul_pkg::tl_a_user_t blanked_auser;
  assign blanked_auser = '{
    rsvd: tl_t_o.a_user.rsvd,
    instr_type: tl_t_o.a_user.instr_type,
    cmd_intg: tlul_pkg::get_bad_cmd_intg(tl_t_o),
    data_intg: tlul_pkg::get_bad_data_intg(tlul_pkg::BlankedAData)
  };

  // if a host is not selected, or if requests are held off, blank the bus
  for (genvar i = 0 ; i < N ; i++) begin : gen_u_o
    logic dev_select;
    assign dev_select = dev_select_t == NWD'(i) & ~hold_all_requests;

    assign tl_u_o[i].a_valid   = tl_t_o.a_valid & dev_select;
    assign tl_u_o[i].a_opcode  = tl_t_o.a_opcode;
    assign tl_u_o[i].a_param   = tl_t_o.a_param;
    assign tl_u_o[i].a_size    = tl_t_o.a_size;
    assign tl_u_o[i].a_source  = tl_t_o.a_source;
    assign tl_u_o[i].a_address = tl_t_o.a_address;
    assign tl_u_o[i].a_mask    = tl_t_o.a_mask;
    assign tl_u_o[i].a_data    = dev_select ?
                                 tl_t_o.a_data :
                                 tlul_pkg::BlankedAData;
    assign tl_u_o[i].a_user    = dev_select ?
                                 tl_t_o.a_user :
                                 blanked_auser;

    assign tl_u_o[i].d_ready   = tl_t_o.d_ready;
  end


  tlul_pkg::tl_d2h_t tl_t_p ;

  // for the returning reqready, only look at the device we're addressing
  logic hfifo_reqready;
  always_comb begin
    hfifo_reqready = tl_u_i[N].a_ready; // default to error
    for (int idx = 0 ; idx < N ; idx++) begin
      //if (dev_select_outstanding == NWD'(idx)) hfifo_reqready = tl_u_i[idx].a_ready;
      if (dev_select_t == NWD'(idx)) hfifo_reqready = tl_u_i[idx].a_ready;
    end
    if (hold_all_requests) hfifo_reqready = 1'b0;
  end
  // Adding a_valid as a qualifier. This prevents the a_ready from having unknown value
  // when the address is unknown and the Host TL-UL FIFO is bypass mode.
  assign tl_t_i.a_ready = tl_t_o.a_valid & hfifo_reqready;

  always_comb begin
    tl_t_p = tl_u_i[N];
    for (int idx = 0 ; idx < N ; idx++) begin
      if (dev_select_outstanding == NWD'(idx)) tl_t_p = tl_u_i[idx];
    end
  end
  assign tl_t_i.d_valid  = tl_t_p.d_valid ;
  assign tl_t_i.d_opcode = tl_t_p.d_opcode;
  assign tl_t_i.d_param  = tl_t_p.d_param ;
  assign tl_t_i.d_size   = tl_t_p.d_size  ;
  assign tl_t_i.d_source = tl_t_p.d_source;
  assign tl_t_i.d_sink   = tl_t_p.d_sink  ;
  assign tl_t_i.d_data   = tl_t_p.d_data  ;
  assign tl_t_i.d_user   = tl_t_p.d_user  ;
  assign tl_t_i.d_error  = tl_t_p.d_error ;

  // Instantiate all the device FIFOs
  for (genvar i = 0 ; i < N ; i++) begin : gen_dfifo
    tlul_fifo_sync #(
      .ReqPass(DReqPass[i]),
      .RspPass(DRspPass[i]),
      .ReqDepth(DReqDepth[i*4+:4]),
      .RspDepth(DRspDepth[i*4+:4])
    ) fifo_d (
      .clk_i,
      .rst_ni,
      .tl_h_i      (tl_u_o[i]),
      .tl_h_o      (tl_u_i[i]),
      .tl_d_o      (tl_d_o[i]),
      .tl_d_i      (tl_d_i[i]),
      .spare_req_i (1'b0),
      .spare_req_o (),
      .spare_rsp_i (1'b0),
      .spare_rsp_o ());
  end

  // Instantiate the error responder. It's only needed if a value greater than
  // N-1 is actually representable in NWD bits.
  if ($clog2(N+1) <= NWD) begin : gen_err_resp
    assign tl_u_o[N].d_ready     = tl_t_o.d_ready;
    assign tl_u_o[N].a_valid     = tl_t_o.a_valid &
                                   (dev_select_t >= NWD'(N)) &
                                   ~hold_all_requests;
    assign tl_u_o[N].a_opcode    = tl_t_o.a_opcode;
    assign tl_u_o[N].a_param     = tl_t_o.a_param;
    assign tl_u_o[N].a_size      = tl_t_o.a_size;
    assign tl_u_o[N].a_source    = tl_t_o.a_source;
    assign tl_u_o[N].a_address   = tl_t_o.a_address;
    assign tl_u_o[N].a_mask      = tl_t_o.a_mask;
    assign tl_u_o[N].a_data      = tl_t_o.a_data;
    assign tl_u_o[N].a_user      = tl_t_o.a_user;
    tlul_err_resp err_resp (
      .clk_i,
      .rst_ni,
      .tl_h_i     (tl_u_o[N]),
      .tl_h_o     (tl_u_i[N])
    );
  end else begin : gen_no_err_resp // block: gen_err_resp
    assign tl_u_o[N] = '0;
    assign tl_u_i[N] = '0;
    logic unused_sig;
    assign unused_sig = ^tl_u_o[N];
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// TL-UL socket M:1 module
//
// Verilog parameters
//   M:             Number of host ports.
//   HReqPass:      M bit array to allow requests to pass through the host i
//                  FIFO with no clock delay if the request FIFO is empty. If
//                  1'b0, at least one clock cycle of latency is created.
//                  Default is 1'b1.
//   HRspPass:      Same as HReqPass but for host response FIFO.
//   HReqDepth:     Mx4 bit array. bit[i*4+:4] is depth of host i request FIFO.
//                  Depth of zero is allowed if ReqPass is true. A maximum value
//                  of 16 is allowed, default is 2.
//   HRspDepth:     Same as HReqDepth but for host response FIFO.
//   DReqPass:      Same as HReqPass but for device request FIFO.
//   DRspPass:      Same as HReqPass but for device response FIFO.
//   DReqDepth:     Same as HReqDepth but for device request FIFO.
//   DRspDepth:     Same as HReqDepth but for device response FIFO.

`include "prim_assert.sv"

module tlul_socket_m1 #(
  parameter int unsigned  M         = 4,
  parameter bit [M-1:0]   HReqPass  = {M{1'b1}},
  parameter bit [M-1:0]   HRspPass  = {M{1'b1}},
  parameter bit [M*4-1:0] HReqDepth = {M{4'h1}},
  parameter bit [M*4-1:0] HRspDepth = {M{4'h1}},
  parameter bit           DReqPass  = 1'b1,
  parameter bit           DRspPass  = 1'b1,
  parameter bit [3:0]     DReqDepth = 4'h1,
  parameter bit [3:0]     DRspDepth = 4'h1
) (
  input                     clk_i,
  input                     rst_ni,

  input  tlul_pkg::tl_h2d_t tl_h_i [M],
  output tlul_pkg::tl_d2h_t tl_h_o [M],

  output tlul_pkg::tl_h2d_t tl_d_o,
  input  tlul_pkg::tl_d2h_t tl_d_i
);

  `ASSERT_INIT(maxM, M < 16)


  // Signals
  //
  //  tl_h_i/o[0] |  tl_h_i/o[1] | ... |  tl_h_i/o[M-1]
  //      |              |                    |
  // u_hostfifo[0]  u_hostfifo[1]        u_hostfifo[M-1]
  //      |              |                    |
  //       hreq_fifo_o(i) / hrsp_fifo_i(i)
  //     ---------------------------------------
  //     |       request/grant/req_data        |
  //     |                                     |
  //     |           PRIM_ARBITER              |
  //     |                                     |
  //     |  arb_valid / arb_ready / arb_data   |
  //     ---------------------------------------
  //                     |
  //                dreq_fifo_i / drsp_fifo_o
  //                     |
  //                u_devicefifo
  //                     |
  //                  tl_d_o/i
  //
  // Required ID width to distinguish between host ports
  //  Used in response steering
  localparam int unsigned IDW   = top_pkg::TL_AIW;
  // localparam int unsigned STIDW = $clog2(M);
  localparam int unsigned STIDW = 1;

  tlul_pkg::tl_h2d_t hreq_fifo_o [M];
  tlul_pkg::tl_d2h_t hrsp_fifo_i [M];

  logic [M-1:0] hrequest;
  logic [M-1:0] hgrant;

  tlul_pkg::tl_h2d_t dreq_fifo_i;
  tlul_pkg::tl_d2h_t drsp_fifo_o;

  logic arb_valid;
  logic arb_ready;
  tlul_pkg::tl_h2d_t arb_data;

  // Host Req/Rsp FIFO
  for (genvar i = 0 ; i < M ; i++) begin : gen_host_fifo
    tlul_pkg::tl_h2d_t hreq_fifo_i;

    // ID Shifting
    logic [STIDW-1:0] reqid_sub;
    logic [IDW-1:0] shifted_id;
    assign reqid_sub = i;   // can cause conversion error?
    assign shifted_id = {
      tl_h_i[i].a_source[0+:(IDW-STIDW)],
      reqid_sub
    };

  `ASSERT(idInRange, tl_h_i[i].a_valid |-> tl_h_i[i].a_source[IDW-1 -:STIDW] == '0)

    // assign not connected bits to nc_* signal to make lint happy
    logic [IDW-1 : IDW-STIDW] unused_tl_h_source;
    assign unused_tl_h_source = tl_h_i[i].a_source[IDW-1 -: STIDW];

    // Put shifted ID
    assign hreq_fifo_i = '{
      a_valid:    tl_h_i[i].a_valid,
      a_opcode:   tl_h_i[i].a_opcode,
      a_param:    tl_h_i[i].a_param,
      a_size:     tl_h_i[i].a_size,
      a_source:   shifted_id,
      a_address:  tl_h_i[i].a_address,
      a_mask:     tl_h_i[i].a_mask,
      a_data:     tl_h_i[i].a_data,
      a_user:     tl_h_i[i].a_user,
      d_ready:    tl_h_i[i].d_ready
    };

    tlul_fifo_sync #(
      .ReqPass    (HReqPass[i]),
      .RspPass    (HRspPass[i]),
      .ReqDepth   (HReqDepth[i*4+:4]),
      .RspDepth   (HRspDepth[i*4+:4]),
      .SpareReqW  (1)
    ) u_hostfifo (
      .clk_i,
      .rst_ni,
      .tl_h_i      (hreq_fifo_i),
      .tl_h_o      (tl_h_o[i]),
      .tl_d_o      (hreq_fifo_o[i]),
      .tl_d_i      (hrsp_fifo_i[i]),
      .spare_req_i (1'b0),
      .spare_req_o (),
      .spare_rsp_i (1'b0),
      .spare_rsp_o ()
    );
  end

  // Device Req/Rsp FIFO
  tlul_fifo_sync #(
    .ReqPass    (DReqPass),
    .RspPass    (DRspPass),
    .ReqDepth   (DReqDepth),
    .RspDepth   (DRspDepth),
    .SpareReqW  (1)
  ) u_devicefifo (
    .clk_i,
    .rst_ni,
    .tl_h_i      (dreq_fifo_i),
    .tl_h_o      (drsp_fifo_o),
    .tl_d_o      (tl_d_o),
    .tl_d_i      (tl_d_i),
    .spare_req_i (1'b0),
    .spare_req_o (),
    .spare_rsp_i (1'b0),
    .spare_rsp_o ()
  );

  // Request Arbiter
  for (genvar i = 0 ; i < M ; i++) begin : gen_arbreqgnt
    assign hrequest[i] = hreq_fifo_o[i].a_valid;
  end

  assign arb_ready = drsp_fifo_o.a_ready;

  if (tlul_pkg::ArbiterImpl == "PPC") begin : gen_arb_ppc
    prim_arbiter_ppc #(
      .N          (M),
      .DW         ($bits(tlul_pkg::tl_h2d_t))
    ) u_reqarb (
      .clk_i,
      .rst_ni,
      .req_chk_i ( 1'b0        ), // TL-UL allows dropping valid without ready. See #3354.
      .req_i     ( hrequest    ),
      .data_i    ( hreq_fifo_o ),
      .gnt_o     ( hgrant      ),
      .idx_o     (             ),
      .valid_o   ( arb_valid   ),
      .data_o    ( arb_data    ),
      .ready_i   ( arb_ready   )
    );
  end else if (tlul_pkg::ArbiterImpl == "BINTREE") begin : gen_tree_arb
    prim_arbiter_tree #(
      .N          (M),
      .DW         ($bits(tlul_pkg::tl_h2d_t))
    ) u_reqarb (
      .clk_i,
      .rst_ni,
      .req_chk_i ( 1'b0        ), // TL-UL allows dropping valid without ready. See #3354.
      .req_i     ( hrequest    ),
      .data_i    ( hreq_fifo_o ),
      .gnt_o     ( hgrant      ),
      .idx_o     (             ),
      .valid_o   ( arb_valid   ),
      .data_o    ( arb_data    ),
      .ready_i   ( arb_ready   )
    );
  end else begin : gen_unknown
    `ASSERT_INIT(UnknownArbImpl_A, 0)
  end

  logic [  M-1:0] hfifo_rspvalid;
  logic [  M-1:0] dfifo_rspready;
  logic [IDW-1:0] hfifo_rspid;
  logic dfifo_rspready_merged;

  // arb_data --> dreq_fifo_i
  //   dreq_fifo_i.hd_rspready <= dfifo_rspready

  assign dfifo_rspready_merged = |dfifo_rspready;
  assign dreq_fifo_i = '{
    a_valid:   arb_valid,
    a_opcode:  arb_data.a_opcode,
    a_param:   arb_data.a_param,
    a_size:    arb_data.a_size,
    a_source:  arb_data.a_source,
    a_address: arb_data.a_address,
    a_mask:    arb_data.a_mask,
    a_data:    arb_data.a_data,
    a_user:    arb_data.a_user,

    d_ready:   dfifo_rspready_merged
  };

  // Response ID steering
  // drsp_fifo_o --> hrsp_fifo_i[i]

  // Response ID shifting before put into host fifo
  assign hfifo_rspid = {
    {STIDW{1'b0}},
    drsp_fifo_o.d_source[IDW-1:STIDW]
  };
  for (genvar i = 0 ; i < M ; i++) begin : gen_idrouting
    assign hfifo_rspvalid[i] = drsp_fifo_o.d_valid &
                               (drsp_fifo_o.d_source[0+:STIDW] == i);
    assign dfifo_rspready[i] = hreq_fifo_o[i].d_ready                &
                               (drsp_fifo_o.d_source[0+:STIDW] == i) &
                              drsp_fifo_o.d_valid;

    assign hrsp_fifo_i[i] = '{
      d_valid:  hfifo_rspvalid[i],
      d_opcode: drsp_fifo_o.d_opcode,
      d_param:  drsp_fifo_o.d_param,
      d_size:   drsp_fifo_o.d_size,
      d_source: hfifo_rspid,
      d_sink:   drsp_fifo_o.d_sink,
      d_data:   drsp_fifo_o.d_data,
      d_user:   drsp_fifo_o.d_user,
      d_error:  drsp_fifo_o.d_error,
      a_ready:  hgrant[i]
    };
  end

  // this assertion fails when rspid[0+:STIDW] not in [0..M-1]
  `ASSERT(rspIdInRange, drsp_fifo_o.d_valid |->
      drsp_fifo_o.d_source[0+:STIDW] >= 0 && drsp_fifo_o.d_source[0+:STIDW] < M)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SRAM interface to TL-UL converter
//      Current version only supports if TL-UL width and SRAM width are same
//      If SRAM interface requests more than MaxOutstanding cap, it generates
//      error in simulation but not in Silicon.

`include "prim_assert.sv"

module sram2tlul #(
  parameter int                        SramAw = 12,
  parameter int                        SramDw = 32,
  parameter logic [top_pkg::TL_AW-1:0] TlBaseAddr = 'h0  // Base address of SRAM request
) (
  input clk_i,
  input rst_ni,

  output tlul_pkg::tl_h2d_t tl_o,
  input  tlul_pkg::tl_d2h_t tl_i,

  // SRAM
  input                     mem_req_i,
  input                     mem_write_i,
  input        [SramAw-1:0] mem_addr_i,
  input        [SramDw-1:0] mem_wdata_i,
  output logic              mem_rvalid_o,
  output logic [SramDw-1:0] mem_rdata_o,
  output logic        [1:0] mem_error_o
);

  import tlul_pkg::*;

  `ASSERT_INIT(wrongSramDw, SramDw == top_pkg::TL_DW)

  localparam int unsigned SRAM_DWB = $clog2(SramDw/8);

  assign tl_o.a_valid   = mem_req_i;
  assign tl_o.a_opcode  = (mem_write_i) ? PutFullData : Get;
  assign tl_o.a_param   = '0;
  assign tl_o.a_size    = top_pkg::TL_SZW'(SRAM_DWB); // Max Size always
  assign tl_o.a_source  = '0;
  assign tl_o.a_address = TlBaseAddr |
                          {{(top_pkg::TL_AW-SramAw-SRAM_DWB){1'b0}},mem_addr_i,{(SRAM_DWB){1'b0}}};
  assign tl_o.a_mask    = '1;
  assign tl_o.a_data    = mem_wdata_i;
  assign tl_o.a_user    = '0;

  assign tl_o.d_ready   = 1'b1;

  assign mem_rvalid_o   = tl_i.d_valid && (tl_i.d_opcode == AccessAckData);
  assign mem_rdata_o    = tl_i.d_data;
  assign mem_error_o    = {2{tl_i.d_error}};

  // below assertion fails when TL-UL doesn't accept request in a cycle,
  // which is currently not supported by sram2tlul
  `ASSERT(validNotReady, tl_o.a_valid |-> tl_i.a_ready)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package aes_reg_pkg;

  // Param list
  parameter int NumRegsKey = 8;
  parameter int NumRegsIv = 4;
  parameter int NumRegsData = 4;
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 8;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_ctrl_update_err;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_fault;
  } aes_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } aes_reg2hw_key_share0_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } aes_reg2hw_key_share1_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } aes_reg2hw_iv_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } aes_reg2hw_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        re;
  } aes_reg2hw_data_out_mreg_t;

  typedef struct packed {
    struct packed {
      logic [1:0]  q;
      logic        qe;
      logic        re;
    } operation;
    struct packed {
      logic [5:0]  q;
      logic        qe;
      logic        re;
    } mode;
    struct packed {
      logic [2:0]  q;
      logic        qe;
      logic        re;
    } key_len;
    struct packed {
      logic        q;
      logic        qe;
      logic        re;
    } sideload;
    struct packed {
      logic [2:0]  q;
      logic        qe;
      logic        re;
    } prng_reseed_rate;
    struct packed {
      logic        q;
      logic        qe;
      logic        re;
    } manual_operation;
  } aes_reg2hw_ctrl_shadowed_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } key_touch_forces_reseed;
    struct packed {
      logic        q;
    } force_masks;
  } aes_reg2hw_ctrl_aux_shadowed_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } start;
    struct packed {
      logic        q;
    } key_iv_data_in_clear;
    struct packed {
      logic        q;
    } data_out_clear;
    struct packed {
      logic        q;
    } prng_reseed;
  } aes_reg2hw_trigger_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } idle;
    struct packed {
      logic        q;
    } output_lost;
  } aes_reg2hw_status_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } aes_hw2reg_key_share0_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } aes_hw2reg_key_share1_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } aes_hw2reg_iv_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } aes_hw2reg_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } aes_hw2reg_data_out_mreg_t;

  typedef struct packed {
    struct packed {
      logic [1:0]  d;
    } operation;
    struct packed {
      logic [5:0]  d;
    } mode;
    struct packed {
      logic [2:0]  d;
    } key_len;
    struct packed {
      logic        d;
    } sideload;
    struct packed {
      logic [2:0]  d;
    } prng_reseed_rate;
    struct packed {
      logic        d;
    } manual_operation;
  } aes_hw2reg_ctrl_shadowed_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } start;
    struct packed {
      logic        d;
      logic        de;
    } key_iv_data_in_clear;
    struct packed {
      logic        d;
      logic        de;
    } data_out_clear;
    struct packed {
      logic        d;
      logic        de;
    } prng_reseed;
  } aes_hw2reg_trigger_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } idle;
    struct packed {
      logic        d;
      logic        de;
    } stall;
    struct packed {
      logic        d;
      logic        de;
    } output_lost;
    struct packed {
      logic        d;
      logic        de;
    } output_valid;
    struct packed {
      logic        d;
      logic        de;
    } input_ready;
    struct packed {
      logic        d;
      logic        de;
    } alert_recov_ctrl_update_err;
    struct packed {
      logic        d;
      logic        de;
    } alert_fatal_fault;
  } aes_hw2reg_status_reg_t;

  // Register -> HW type
  typedef struct packed {
    aes_reg2hw_alert_test_reg_t alert_test; // [957:954]
    aes_reg2hw_key_share0_mreg_t [7:0] key_share0; // [953:690]
    aes_reg2hw_key_share1_mreg_t [7:0] key_share1; // [689:426]
    aes_reg2hw_iv_mreg_t [3:0] iv; // [425:294]
    aes_reg2hw_data_in_mreg_t [3:0] data_in; // [293:162]
    aes_reg2hw_data_out_mreg_t [3:0] data_out; // [161:30]
    aes_reg2hw_ctrl_shadowed_reg_t ctrl_shadowed; // [29:8]
    aes_reg2hw_ctrl_aux_shadowed_reg_t ctrl_aux_shadowed; // [7:6]
    aes_reg2hw_trigger_reg_t trigger; // [5:2]
    aes_reg2hw_status_reg_t status; // [1:0]
  } aes_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    aes_hw2reg_key_share0_mreg_t [7:0] key_share0; // [937:682]
    aes_hw2reg_key_share1_mreg_t [7:0] key_share1; // [681:426]
    aes_hw2reg_iv_mreg_t [3:0] iv; // [425:298]
    aes_hw2reg_data_in_mreg_t [3:0] data_in; // [297:166]
    aes_hw2reg_data_out_mreg_t [3:0] data_out; // [165:38]
    aes_hw2reg_ctrl_shadowed_reg_t ctrl_shadowed; // [37:22]
    aes_hw2reg_trigger_reg_t trigger; // [21:14]
    aes_hw2reg_status_reg_t status; // [13:0]
  } aes_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] AES_ALERT_TEST_OFFSET = 8'h 0;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_0_OFFSET = 8'h 4;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_1_OFFSET = 8'h 8;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_2_OFFSET = 8'h c;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_3_OFFSET = 8'h 10;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_4_OFFSET = 8'h 14;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_5_OFFSET = 8'h 18;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_6_OFFSET = 8'h 1c;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE0_7_OFFSET = 8'h 20;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_0_OFFSET = 8'h 24;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_1_OFFSET = 8'h 28;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_2_OFFSET = 8'h 2c;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_3_OFFSET = 8'h 30;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_4_OFFSET = 8'h 34;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_5_OFFSET = 8'h 38;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_6_OFFSET = 8'h 3c;
  parameter logic [BlockAw-1:0] AES_KEY_SHARE1_7_OFFSET = 8'h 40;
  parameter logic [BlockAw-1:0] AES_IV_0_OFFSET = 8'h 44;
  parameter logic [BlockAw-1:0] AES_IV_1_OFFSET = 8'h 48;
  parameter logic [BlockAw-1:0] AES_IV_2_OFFSET = 8'h 4c;
  parameter logic [BlockAw-1:0] AES_IV_3_OFFSET = 8'h 50;
  parameter logic [BlockAw-1:0] AES_DATA_IN_0_OFFSET = 8'h 54;
  parameter logic [BlockAw-1:0] AES_DATA_IN_1_OFFSET = 8'h 58;
  parameter logic [BlockAw-1:0] AES_DATA_IN_2_OFFSET = 8'h 5c;
  parameter logic [BlockAw-1:0] AES_DATA_IN_3_OFFSET = 8'h 60;
  parameter logic [BlockAw-1:0] AES_DATA_OUT_0_OFFSET = 8'h 64;
  parameter logic [BlockAw-1:0] AES_DATA_OUT_1_OFFSET = 8'h 68;
  parameter logic [BlockAw-1:0] AES_DATA_OUT_2_OFFSET = 8'h 6c;
  parameter logic [BlockAw-1:0] AES_DATA_OUT_3_OFFSET = 8'h 70;
  parameter logic [BlockAw-1:0] AES_CTRL_SHADOWED_OFFSET = 8'h 74;
  parameter logic [BlockAw-1:0] AES_CTRL_AUX_SHADOWED_OFFSET = 8'h 78;
  parameter logic [BlockAw-1:0] AES_CTRL_AUX_REGWEN_OFFSET = 8'h 7c;
  parameter logic [BlockAw-1:0] AES_TRIGGER_OFFSET = 8'h 80;
  parameter logic [BlockAw-1:0] AES_STATUS_OFFSET = 8'h 84;

  // Reset values for hwext registers and their fields
  parameter logic [1:0] AES_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] AES_ALERT_TEST_RECOV_CTRL_UPDATE_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] AES_ALERT_TEST_FATAL_FAULT_RESVAL = 1'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_0_KEY_SHARE0_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_1_KEY_SHARE0_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_2_KEY_SHARE0_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_3_KEY_SHARE0_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_4_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_4_KEY_SHARE0_4_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_5_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_5_KEY_SHARE0_5_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_6_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_6_KEY_SHARE0_6_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_7_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE0_7_KEY_SHARE0_7_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_0_KEY_SHARE1_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_1_KEY_SHARE1_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_2_KEY_SHARE1_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_3_KEY_SHARE1_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_4_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_4_KEY_SHARE1_4_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_5_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_5_KEY_SHARE1_5_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_6_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_6_KEY_SHARE1_6_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_7_RESVAL = 32'h 0;
  parameter logic [31:0] AES_KEY_SHARE1_7_KEY_SHARE1_7_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_0_IV_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_1_IV_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_2_IV_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_IV_3_IV_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_0_DATA_OUT_0_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_1_DATA_OUT_1_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_2_DATA_OUT_2_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_3_RESVAL = 32'h 0;
  parameter logic [31:0] AES_DATA_OUT_3_DATA_OUT_3_RESVAL = 32'h 0;
  parameter logic [15:0] AES_CTRL_SHADOWED_RESVAL = 16'h 1181;
  parameter logic [1:0] AES_CTRL_SHADOWED_OPERATION_RESVAL = 2'h 1;
  parameter logic [5:0] AES_CTRL_SHADOWED_MODE_RESVAL = 6'h 20;
  parameter logic [2:0] AES_CTRL_SHADOWED_KEY_LEN_RESVAL = 3'h 1;
  parameter logic [0:0] AES_CTRL_SHADOWED_SIDELOAD_RESVAL = 1'h 0;
  parameter logic [2:0] AES_CTRL_SHADOWED_PRNG_RESEED_RATE_RESVAL = 3'h 1;
  parameter logic [0:0] AES_CTRL_SHADOWED_MANUAL_OPERATION_RESVAL = 1'h 0;

  // Register index
  typedef enum int {
    AES_ALERT_TEST,
    AES_KEY_SHARE0_0,
    AES_KEY_SHARE0_1,
    AES_KEY_SHARE0_2,
    AES_KEY_SHARE0_3,
    AES_KEY_SHARE0_4,
    AES_KEY_SHARE0_5,
    AES_KEY_SHARE0_6,
    AES_KEY_SHARE0_7,
    AES_KEY_SHARE1_0,
    AES_KEY_SHARE1_1,
    AES_KEY_SHARE1_2,
    AES_KEY_SHARE1_3,
    AES_KEY_SHARE1_4,
    AES_KEY_SHARE1_5,
    AES_KEY_SHARE1_6,
    AES_KEY_SHARE1_7,
    AES_IV_0,
    AES_IV_1,
    AES_IV_2,
    AES_IV_3,
    AES_DATA_IN_0,
    AES_DATA_IN_1,
    AES_DATA_IN_2,
    AES_DATA_IN_3,
    AES_DATA_OUT_0,
    AES_DATA_OUT_1,
    AES_DATA_OUT_2,
    AES_DATA_OUT_3,
    AES_CTRL_SHADOWED,
    AES_CTRL_AUX_SHADOWED,
    AES_CTRL_AUX_REGWEN,
    AES_TRIGGER,
    AES_STATUS
  } aes_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] AES_PERMIT [34] = '{
    4'b 0001, // index[ 0] AES_ALERT_TEST
    4'b 1111, // index[ 1] AES_KEY_SHARE0_0
    4'b 1111, // index[ 2] AES_KEY_SHARE0_1
    4'b 1111, // index[ 3] AES_KEY_SHARE0_2
    4'b 1111, // index[ 4] AES_KEY_SHARE0_3
    4'b 1111, // index[ 5] AES_KEY_SHARE0_4
    4'b 1111, // index[ 6] AES_KEY_SHARE0_5
    4'b 1111, // index[ 7] AES_KEY_SHARE0_6
    4'b 1111, // index[ 8] AES_KEY_SHARE0_7
    4'b 1111, // index[ 9] AES_KEY_SHARE1_0
    4'b 1111, // index[10] AES_KEY_SHARE1_1
    4'b 1111, // index[11] AES_KEY_SHARE1_2
    4'b 1111, // index[12] AES_KEY_SHARE1_3
    4'b 1111, // index[13] AES_KEY_SHARE1_4
    4'b 1111, // index[14] AES_KEY_SHARE1_5
    4'b 1111, // index[15] AES_KEY_SHARE1_6
    4'b 1111, // index[16] AES_KEY_SHARE1_7
    4'b 1111, // index[17] AES_IV_0
    4'b 1111, // index[18] AES_IV_1
    4'b 1111, // index[19] AES_IV_2
    4'b 1111, // index[20] AES_IV_3
    4'b 1111, // index[21] AES_DATA_IN_0
    4'b 1111, // index[22] AES_DATA_IN_1
    4'b 1111, // index[23] AES_DATA_IN_2
    4'b 1111, // index[24] AES_DATA_IN_3
    4'b 1111, // index[25] AES_DATA_OUT_0
    4'b 1111, // index[26] AES_DATA_OUT_1
    4'b 1111, // index[27] AES_DATA_OUT_2
    4'b 1111, // index[28] AES_DATA_OUT_3
    4'b 0011, // index[29] AES_CTRL_SHADOWED
    4'b 0001, // index[30] AES_CTRL_AUX_SHADOWED
    4'b 0001, // index[31] AES_CTRL_AUX_REGWEN
    4'b 0001, // index[32] AES_TRIGGER
    4'b 0001  // index[33] AES_STATUS
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES package

package aes_pkg;

// If this parameter is set, fatal alerts clear all status and trigger bits to zero. By
// default, it's not set, i.e., no clearing is happening, in order to simplify debugging.
parameter bit ClearStatusOnFatalAlert = 1'b0;

// The initial key is always provided in two shares, independently whether the cipher core is
// masked or not.
parameter int unsigned NumSharesKey = 2;

// Software updates IV in chunks of 32 bits, the counter updates 16 bits at a time.
parameter int unsigned SliceSizeCtr = 16;
parameter int unsigned NumSlicesCtr = aes_reg_pkg::NumRegsIv * 32 / SliceSizeCtr;
parameter int unsigned SliceIdxWidth = prim_util_pkg::vbits(NumSlicesCtr);

// Widths of signals carrying pseudo-random data for clearing
parameter int unsigned WidthPRDClearing = 64;
parameter int unsigned NumChunksPRDClearing128 = 128/WidthPRDClearing;
parameter int unsigned NumChunksPRDClearing256 = 256/WidthPRDClearing;

// Widths of signals carrying pseudo-random data for masking
parameter int unsigned WidthPRDSBox     = 8;  // Number PRD bits per S-Box. This includes the
                                              // 8 bits for the output mask when using any of the
                                              // masked Canright S-Box implementations.
parameter int unsigned WidthPRDData     = 16*WidthPRDSBox; // 16 S-Boxes for the data path
parameter int unsigned WidthPRDKey      = 4*WidthPRDSBox;  // 4 S-Boxes for the key expand
parameter int unsigned WidthPRDMasking  = WidthPRDData + WidthPRDKey;

parameter int unsigned ChunkSizePRDMasking = WidthPRDMasking/5;

// Clearing PRNG default LFSR seed and permutation
// These LFSR parameters have been generated with
// $ util/design/gen-lfsr-seed.py --width 64 --seed 31468618 --prefix "Clearing"
parameter int ClearingLfsrWidth = 64;
typedef logic [ClearingLfsrWidth-1:0] clearing_lfsr_seed_t;
typedef logic [ClearingLfsrWidth-1:0][$clog2(ClearingLfsrWidth)-1:0] clearing_lfsr_perm_t;
parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeedDefault = 64'hc32d580f74f1713a;
parameter clearing_lfsr_perm_t RndCnstClearingLfsrPermDefault = {
  128'hb33fdfc81deb6292c21f8a3102585067,
  256'h9c2f4be1bbe937b4b7c9d7f4e57568d99c8ae291a899143e0d8459d31b143223
};
// A second permutation is needed for the second share.
parameter clearing_lfsr_perm_t RndCnstClearingSharePermDefault = {
  128'hf66fd61b27847edc2286706fb3a2e900,
  256'h9736b95ac3f3b5205caf8dc536aad73605d393c8dd94476e830e97891d4828d0
};

// Masking PRNG default LFSR seed and permutation
// We use a single seed that is split down into chunks internally.
// These LFSR parameters have been generated with
// $ util/design/gen-lfsr-seed.py --width 160 --seed 31468618 --prefix "Masking"
parameter int MaskingLfsrWidth = 160; // = WidthPRDMasking = WidthPRDSBox * (16 + 4)
typedef logic [MaskingLfsrWidth-1:0] masking_lfsr_seed_t;
typedef logic [MaskingLfsrWidth-1:0][$clog2(MaskingLfsrWidth)-1:0] masking_lfsr_perm_t;
parameter masking_lfsr_seed_t RndCnstMaskingLfsrSeedDefault =
  160'hc132b5723c5a4cf4743b3c7c32d580f74f1713a;
parameter masking_lfsr_perm_t RndCnstMaskingLfsrPermDefault = {
  256'h17261943423e4c5c03872194050c7e5f8497081d96666d406f4b606473303469,
  256'h8e7c721c8832471f59919e0b128f067b25622768462e554d8970815d490d7f44,
  256'h048c867d907a239b20220f6c79071a852d76485452189f14091b1e744e396737,
  256'h4f785b772b352f6550613c58130a8b104a3f28019c9a380233956b00563a512c,
  256'h808d419d63982a16995e0e3b57826a36718a9329452492533d83115a75316e15
};

typedef enum integer {
  SBoxImplLut,                   // Unmasked LUT-based S-Box
  SBoxImplCanright,              // Unmasked Canright S-Box, see aes_sbox_canright.sv
  SBoxImplCanrightMasked,        // First-order masked Canright S-Box
                                 // see aes_sbox_canright_masked.sv
  SBoxImplCanrightMaskedNoreuse, // First-order masked Canright S-Box without mask reuse,
                                 // see aes_sbox_canright_masked_noreuse.sv
  SBoxImplDom                    // First-order masked S-Box using domain-oriented masking,
                                 // see aes_sbox_canright_dom.sv
} sbox_impl_e;


// Parameters used for controlgroups in the coverage
parameter int AES_OP_WIDTH             = 2;
parameter int AES_MODE_WIDTH           = 6;
parameter int AES_KEYLEN_WIDTH         = 3;
parameter int AES_PRNGRESEEDRATE_WIDTH = 3;

// SEC_CM: MAIN.CONFIG.SPARSE
typedef enum logic [AES_OP_WIDTH-1:0] {
  AES_ENC = 2'b01,
  AES_DEC = 2'b10
} aes_op_e;

// SEC_CM: MAIN.CONFIG.SPARSE
typedef enum logic [AES_MODE_WIDTH-1:0] {
  AES_ECB  = 6'b00_0001,
  AES_CBC  = 6'b00_0010,
  AES_CFB  = 6'b00_0100,
  AES_OFB  = 6'b00_1000,
  AES_CTR  = 6'b01_0000,
  AES_NONE = 6'b10_0000
} aes_mode_e;

typedef enum logic [AES_OP_WIDTH-1:0] {
  CIPH_FWD = 2'b01,
  CIPH_INV = 2'b10
} ciph_op_e;

// SEC_CM: MAIN.CONFIG.SPARSE
typedef enum logic [AES_KEYLEN_WIDTH-1:0] {
  AES_128 = 3'b001,
  AES_192 = 3'b010,
  AES_256 = 3'b100
} key_len_e;

// SEC_CM: MAIN.CONFIG.SPARSE
typedef enum logic [AES_PRNGRESEEDRATE_WIDTH-1:0] {
  PER_1  = 3'b001,
  PER_64 = 3'b010,
  PER_8K = 3'b100
} prs_rate_e;
parameter int unsigned BlockCtrWidth = 13;

typedef struct packed {
  logic [31:7] unused;
  logic        alert_fatal_fault;
  logic        alert_recov_ctrl_update_err;
  logic        input_ready;
  logic        output_valid;
  logic        output_lost;
  logic        stall;
  logic        idle;
} status_t;

typedef struct packed {
  logic        recov_ctrl_update_err;
  logic        fatal_fault;
} alert_test_t;

  // Sparse state encodings

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 8 -n 6 \
  //      -s 31468618 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (57.14%)
  //  4: ||||||||||||||| (42.86%)
  //  5: --
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 5
  //
  localparam int CipherCtrlStateWidth = 6;
  typedef enum logic [CipherCtrlStateWidth-1:0] {
    CIPHER_CTRL_IDLE        = 6'b001001,
    CIPHER_CTRL_INIT        = 6'b100011,
    CIPHER_CTRL_ROUND       = 6'b111101,
    CIPHER_CTRL_FINISH      = 6'b010000,
    CIPHER_CTRL_PRNG_RESEED = 6'b100100,
    CIPHER_CTRL_CLEAR_S     = 6'b111010,
    CIPHER_CTRL_CLEAR_KD    = 6'b001110,
    CIPHER_CTRL_ERROR       = 6'b010111
  } aes_cipher_ctrl_e;

  // $ ./sparse-fsm-encode.py -d 3 -m 3 -n 5 \
  //      -s 31468618 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (66.67%)
  //  4: |||||||||| (33.33%)
  //  5: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  //
  localparam int CtrStateWidth = 5;
  typedef enum logic [CtrStateWidth-1:0] {
    CTR_IDLE  = 5'b01110,
    CTR_INCR  = 5'b11000,
    CTR_ERROR = 5'b00001
  } aes_ctr_e;

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 8 -n 6 \
  //      -s 31468618 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (57.14%)
  //  4: ||||||||||||||| (42.86%)
  //  5: --
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 5
  //
  localparam int CtrlStateWidth = 6;
  typedef enum logic [CtrlStateWidth-1:0] {
    CTRL_IDLE        = 6'b001001,
    CTRL_LOAD        = 6'b100011,
    CTRL_PRNG_UPDATE = 6'b111101,
    CTRL_PRNG_RESEED = 6'b010000,
    CTRL_FINISH      = 6'b100100,
    CTRL_CLEAR_I     = 6'b111010,
    CTRL_CLEAR_CO    = 6'b001110,
    CTRL_ERROR       = 6'b010111
  } aes_ctrl_e;

// Generic, sparse mux selector encodings

// Encoding generated with:
// $ ./util/design/sparse-fsm-encode.py -d 3 -m 2 -n 3 \
//      -s 31468618 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (100.00%)
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 3
// Minimum Hamming weight: 1
// Maximum Hamming weight: 2
//
parameter int Mux2SelWidth = 3;
typedef enum logic [Mux2SelWidth-1:0] {
  MUX2_SEL_0 = 3'b011,
  MUX2_SEL_1 = 3'b100
} mux2_sel_e;

// Encoding generated with:
// $ ./sparse-fsm-encode.py -d 3 -m 3 -n 5 \
//      -s 31468618 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (66.67%)
//  4: |||||||||| (33.33%)
//  5: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 4
//
parameter int Mux3SelWidth = 5;
typedef enum logic [Mux3SelWidth-1:0] {
  MUX3_SEL_0 = 5'b01110,
  MUX3_SEL_1 = 5'b11000,
  MUX3_SEL_2 = 5'b00001
} mux3_sel_e;

// Encoding generated with:
// $ ./sparse-fsm-encode.py -d 3 -m 4 -n 5 \
//      -s 31468618 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (66.67%)
//  4: |||||||||| (33.33%)
//  5: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 4
//
parameter int Mux4SelWidth = 5;
typedef enum logic [Mux4SelWidth-1:0] {
  MUX4_SEL_0 = 5'b01110,
  MUX4_SEL_1 = 5'b11000,
  MUX4_SEL_2 = 5'b00001,
  MUX4_SEL_3 = 5'b10111
} mux4_sel_e;

// $ ./sparse-fsm-encode.py -d 3 -m 6 -n 6 \
//      -s 31468618 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (53.33%)
//  4: ||||||||||||||| (40.00%)
//  5: || (6.67%)
//  6: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 5
//
parameter int Mux6SelWidth = 6;
typedef enum logic [Mux6SelWidth-1:0] {
  MUX6_SEL_0 = 6'b011101,
  MUX6_SEL_1 = 6'b110000,
  MUX6_SEL_2 = 6'b001000,
  MUX6_SEL_3 = 6'b000011,
  MUX6_SEL_4 = 6'b111110,
  MUX6_SEL_5 = 6'b100101
} mux6_sel_e;

// Mux selector signal types. These use the generic types defined above.

parameter int DIPSelNum = 2;
parameter int DIPSelWidth = Mux2SelWidth;
typedef enum logic [DIPSelWidth-1:0] {
  DIP_DATA_IN = MUX2_SEL_0,
  DIP_CLEAR   = MUX2_SEL_1
} dip_sel_e;

parameter int SISelNum = 2;
parameter int SISelWidth = Mux2SelWidth;
typedef enum logic [SISelWidth-1:0] {
  SI_ZERO = MUX2_SEL_0,
  SI_DATA = MUX2_SEL_1
} si_sel_e;

parameter int AddSISelNum = 2;
parameter int AddSISelWidth = Mux2SelWidth;
typedef enum logic [AddSISelWidth-1:0] {
  ADD_SI_ZERO = MUX2_SEL_0,
  ADD_SI_IV   = MUX2_SEL_1
} add_si_sel_e;

parameter int StateSelNum = 3;
parameter int StateSelWidth = Mux3SelWidth;
typedef enum logic [StateSelWidth-1:0] {
  STATE_INIT  = MUX3_SEL_0,
  STATE_ROUND = MUX3_SEL_1,
  STATE_CLEAR = MUX3_SEL_2
} state_sel_e;

parameter int AddRKSelNum = 3;
parameter int AddRKSelWidth = Mux3SelWidth;
typedef enum logic [AddRKSelWidth-1:0] {
  ADD_RK_INIT  = MUX3_SEL_0,
  ADD_RK_ROUND = MUX3_SEL_1,
  ADD_RK_FINAL = MUX3_SEL_2
} add_rk_sel_e;

parameter int KeyInitSelNum = 3;
parameter int KeyInitSelWidth = Mux3SelWidth;
typedef enum logic [KeyInitSelWidth-1:0] {
  KEY_INIT_INPUT  = MUX3_SEL_0,
  KEY_INIT_KEYMGR = MUX3_SEL_1,
  KEY_INIT_CLEAR  = MUX3_SEL_2
} key_init_sel_e;

parameter int IVSelNum = 6;
parameter int IVSelWidth = Mux6SelWidth;
typedef enum logic [IVSelWidth-1:0] {
  IV_INPUT        = MUX6_SEL_0,
  IV_DATA_OUT     = MUX6_SEL_1,
  IV_DATA_OUT_RAW = MUX6_SEL_2,
  IV_DATA_IN_PREV = MUX6_SEL_3,
  IV_CTR          = MUX6_SEL_4,
  IV_CLEAR        = MUX6_SEL_5
} iv_sel_e;

parameter int KeyFullSelNum = 4;
parameter int KeyFullSelWidth = Mux4SelWidth;
typedef enum logic [KeyFullSelWidth-1:0] {
  KEY_FULL_ENC_INIT = MUX4_SEL_0,
  KEY_FULL_DEC_INIT = MUX4_SEL_1,
  KEY_FULL_ROUND    = MUX4_SEL_2,
  KEY_FULL_CLEAR    = MUX4_SEL_3
} key_full_sel_e;

parameter int KeyDecSelNum = 2;
parameter int KeyDecSelWidth = Mux2SelWidth;
typedef enum logic [KeyDecSelWidth-1:0] {
  KEY_DEC_EXPAND = MUX2_SEL_0,
  KEY_DEC_CLEAR  = MUX2_SEL_1
} key_dec_sel_e;

parameter int KeyWordsSelNum = 4;
parameter int KeyWordsSelWidth = Mux4SelWidth;
typedef enum logic [KeyWordsSelWidth-1:0] {
  KEY_WORDS_0123 = MUX4_SEL_0,
  KEY_WORDS_2345 = MUX4_SEL_1,
  KEY_WORDS_4567 = MUX4_SEL_2,
  KEY_WORDS_ZERO = MUX4_SEL_3
} key_words_sel_e;

parameter int RoundKeySelNum = 2;
parameter int RoundKeySelWidth = Mux2SelWidth;
typedef enum logic [RoundKeySelWidth-1:0] {
  ROUND_KEY_DIRECT = MUX2_SEL_0,
  ROUND_KEY_MIXED  = MUX2_SEL_1
} round_key_sel_e;

parameter int AddSOSelNum = 3;
parameter int AddSOSelWidth = Mux3SelWidth;
typedef enum logic [AddSOSelWidth-1:0] {
  ADD_SO_ZERO = MUX3_SEL_0,
  ADD_SO_IV   = MUX3_SEL_1,
  ADD_SO_DIP  = MUX3_SEL_2
} add_so_sel_e;

// Sparse two-value signal type sp2v_e
parameter int Sp2VNum = 2;
parameter int Sp2VWidth = Mux2SelWidth;
typedef enum logic [Sp2VWidth-1:0] {
  SP2V_HIGH = MUX2_SEL_0,
  SP2V_LOW  = MUX2_SEL_1
} sp2v_e;

typedef logic [Sp2VWidth-1:0] sp2v_logic_t;
parameter sp2v_logic_t SP2V_LOGIC_HIGH = {SP2V_HIGH};

// Control register type
typedef struct packed {
  logic      manual_operation;
  prs_rate_e prng_reseed_rate;
  logic      sideload;
  key_len_e  key_len;
  aes_mode_e mode;
  aes_op_e   operation;
} ctrl_reg_t;

parameter ctrl_reg_t CTRL_RESET = '{
  manual_operation: aes_reg_pkg::AES_CTRL_SHADOWED_MANUAL_OPERATION_RESVAL,
  prng_reseed_rate: prs_rate_e'(aes_reg_pkg::AES_CTRL_SHADOWED_PRNG_RESEED_RATE_RESVAL),
  sideload:         aes_reg_pkg::AES_CTRL_SHADOWED_SIDELOAD_RESVAL,
  key_len:          key_len_e'(aes_reg_pkg::AES_CTRL_SHADOWED_KEY_LEN_RESVAL),
  mode:             aes_mode_e'(aes_reg_pkg::AES_CTRL_SHADOWED_MODE_RESVAL),
  operation:        aes_op_e'(aes_reg_pkg::AES_CTRL_SHADOWED_OPERATION_RESVAL)
};

// Multiplication by {02} (i.e. x) on GF(2^8)
// with field generating polynomial {01}{1b} (9'h11b)
// Sometimes also denoted by xtime().
function automatic logic [7:0] aes_mul2(logic [7:0] in);
  logic [7:0] out;
  out[7] = in[6];
  out[6] = in[5];
  out[5] = in[4];
  out[4] = in[3] ^ in[7];
  out[3] = in[2] ^ in[7];
  out[2] = in[1];
  out[1] = in[0] ^ in[7];
  out[0] = in[7];
  return out;
endfunction

// Multiplication by {04} (i.e. x^2) on GF(2^8)
// with field generating polynomial {01}{1b} (9'h11b)
function automatic logic [7:0] aes_mul4(logic [7:0] in);
  return aes_mul2(aes_mul2(in));
endfunction

// Division by {02} (i.e. x) on GF(2^8)
// with field generating polynomial {01}{1b} (9'h11b)
// This is the inverse of aes_mul2() or xtime().
function automatic logic [7:0] aes_div2(logic [7:0] in);
  logic [7:0] out;
  out[7] = in[0];
  out[6] = in[7];
  out[5] = in[6];
  out[4] = in[5];
  out[3] = in[4] ^ in[0];
  out[2] = in[3] ^ in[0];
  out[1] = in[2];
  out[0] = in[1] ^ in[0];
  return out;
endfunction

// Circular byte shift to the left
function automatic logic [31:0] aes_circ_byte_shift(logic [31:0] in, logic [1:0] shift);
  logic [31:0] out;
  logic [31:0] s;
  s = {30'b0,shift};
  out = {in[8*((7-s)%4) +: 8], in[8*((6-s)%4) +: 8],
         in[8*((5-s)%4) +: 8], in[8*((4-s)%4) +: 8]};
  return out;
endfunction

// Transpose state matrix
function automatic logic [3:0][3:0][7:0] aes_transpose(logic [3:0][3:0][7:0] in);
  logic [3:0][3:0][7:0] transpose;
  transpose = '0;
  for (int j = 0; j < 4; j++) begin
    for (int i = 0; i < 4; i++) begin
      transpose[i][j] = in[j][i];
    end
  end
  return transpose;
endfunction

// Extract single column from state matrix
function automatic logic [3:0][7:0] aes_col_get(logic [3:0][3:0][7:0] in, logic [1:0] idx);
  logic [3:0][7:0] out;
  for (int i = 0; i < 4; i++) begin
    out[i] = in[i][idx];
  end
  return out;
endfunction

// Matrix-vector multiplication in GF(2^8): c = A * b
function automatic logic [7:0] aes_mvm(
  logic [7:0] vec_b,
  logic [7:0] mat_a [8]
);
  logic [7:0] vec_c;
  vec_c = '0;
  for (int i = 0; i < 8; i++) begin
    for (int j = 0; j < 8; j++) begin
      vec_c[i] = vec_c[i] ^ (mat_a[j][i] & vec_b[7-j]);
    end
  end
  return vec_c;
endfunction

// Rotate integer indices
function automatic integer aes_rot_int(integer in, integer num);
  integer out;
  if (in == 0) begin
    out = num - 1;
  end else begin
    out = in - 1;
  end
  return out;
endfunction

// Function for extracting LSBs of the per-S-Box pseudo-random data (PRD) from the output of the
// masking PRNG.
//
// The masking PRNG is used for generating both the PRD for the S-Boxes/SubBytes operation as
// well as for the input data masks. When using any of the masked Canright S-Box implementations,
// it is important that the SubBytes input masks (generated by the PRNG in Round X-1) and the
// SubBytes output masks (generated by the PRNG in Round X) are independent. Inside the PRNG,
// this is achieved by using multiple, separately re-seeded LFSR chunks and by selecting the
// separate LFSR chunks in alternating fashion. Since the input data masks become the SubBytes
// input masks in the first round, we select the same 8 bit lanes for the input data masks which
// are also used to form the SubBytes output mask for the masked Canright S-Box implementations,
// i.e., the 8 LSBs of the per S-Box PRD. In particular, we have:
//
// prng_output = { prd_key_expand, ... , sb_prd[4], sb_out_mask[4], sb_prd[0], sb_out_mask[0] }
//
// Where sb_out_mask[x] contains the SubBytes output mask for byte x (when using a masked
// Canright S-Box implementation) and sb_prd[x] contains additional PRD consumed by SubBytes for
// byte x.
//
// When using a masked S-Box implementation other than Canright, we still select the 8 LSBs of
// the per-S-Box PRD to form the input data mask of the corresponding byte. We do this to
// distribute the input data masks over all LFSR chunks of the masking PRNG.

// For one row of the state matrix, extract the 8 LSBs of the per-S-Box PRD from the PRNG output.
// These bits are used as:
// - input data masks, and
// - SubBytes output mask when using a masked Canright S-Box implementation.
function automatic logic [3:0][7:0] aes_prd_get_lsbs(
  logic [(4*WidthPRDSBox)-1:0] in
);
  logic [3:0][7:0] prd_lsbs;
  for (int i = 0; i < 4; i++) begin
    prd_lsbs[i] = in[i*WidthPRDSBox +: 8];
  end
  return prd_lsbs;
endfunction

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module aes_reg_top (
  input clk_i,
  input rst_ni,
  input rst_shadowed_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output aes_reg_pkg::aes_reg2hw_t reg2hw, // Write
  input  aes_reg_pkg::aes_hw2reg_t hw2reg, // Read

  output logic shadowed_storage_err_o,
  output logic shadowed_update_err_o,

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import aes_reg_pkg::* ;

  localparam int AW = 8;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [33:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(34)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic alert_test_we;
  logic alert_test_recov_ctrl_update_err_wd;
  logic alert_test_fatal_fault_wd;
  logic key_share0_0_we;
  logic [31:0] key_share0_0_wd;
  logic key_share0_1_we;
  logic [31:0] key_share0_1_wd;
  logic key_share0_2_we;
  logic [31:0] key_share0_2_wd;
  logic key_share0_3_we;
  logic [31:0] key_share0_3_wd;
  logic key_share0_4_we;
  logic [31:0] key_share0_4_wd;
  logic key_share0_5_we;
  logic [31:0] key_share0_5_wd;
  logic key_share0_6_we;
  logic [31:0] key_share0_6_wd;
  logic key_share0_7_we;
  logic [31:0] key_share0_7_wd;
  logic key_share1_0_we;
  logic [31:0] key_share1_0_wd;
  logic key_share1_1_we;
  logic [31:0] key_share1_1_wd;
  logic key_share1_2_we;
  logic [31:0] key_share1_2_wd;
  logic key_share1_3_we;
  logic [31:0] key_share1_3_wd;
  logic key_share1_4_we;
  logic [31:0] key_share1_4_wd;
  logic key_share1_5_we;
  logic [31:0] key_share1_5_wd;
  logic key_share1_6_we;
  logic [31:0] key_share1_6_wd;
  logic key_share1_7_we;
  logic [31:0] key_share1_7_wd;
  logic iv_0_re;
  logic iv_0_we;
  logic [31:0] iv_0_qs;
  logic [31:0] iv_0_wd;
  logic iv_1_re;
  logic iv_1_we;
  logic [31:0] iv_1_qs;
  logic [31:0] iv_1_wd;
  logic iv_2_re;
  logic iv_2_we;
  logic [31:0] iv_2_qs;
  logic [31:0] iv_2_wd;
  logic iv_3_re;
  logic iv_3_we;
  logic [31:0] iv_3_qs;
  logic [31:0] iv_3_wd;
  logic data_in_0_we;
  logic [31:0] data_in_0_wd;
  logic data_in_1_we;
  logic [31:0] data_in_1_wd;
  logic data_in_2_we;
  logic [31:0] data_in_2_wd;
  logic data_in_3_we;
  logic [31:0] data_in_3_wd;
  logic data_out_0_re;
  logic [31:0] data_out_0_qs;
  logic data_out_1_re;
  logic [31:0] data_out_1_qs;
  logic data_out_2_re;
  logic [31:0] data_out_2_qs;
  logic data_out_3_re;
  logic [31:0] data_out_3_qs;
  logic ctrl_shadowed_re;
  logic ctrl_shadowed_we;
  logic [1:0] ctrl_shadowed_operation_qs;
  logic [1:0] ctrl_shadowed_operation_wd;
  logic [5:0] ctrl_shadowed_mode_qs;
  logic [5:0] ctrl_shadowed_mode_wd;
  logic [2:0] ctrl_shadowed_key_len_qs;
  logic [2:0] ctrl_shadowed_key_len_wd;
  logic ctrl_shadowed_sideload_qs;
  logic ctrl_shadowed_sideload_wd;
  logic [2:0] ctrl_shadowed_prng_reseed_rate_qs;
  logic [2:0] ctrl_shadowed_prng_reseed_rate_wd;
  logic ctrl_shadowed_manual_operation_qs;
  logic ctrl_shadowed_manual_operation_wd;
  logic ctrl_aux_shadowed_re;
  logic ctrl_aux_shadowed_we;
  logic ctrl_aux_shadowed_key_touch_forces_reseed_qs;
  logic ctrl_aux_shadowed_key_touch_forces_reseed_wd;
  logic ctrl_aux_shadowed_key_touch_forces_reseed_storage_err;
  logic ctrl_aux_shadowed_key_touch_forces_reseed_update_err;
  logic ctrl_aux_shadowed_force_masks_qs;
  logic ctrl_aux_shadowed_force_masks_wd;
  logic ctrl_aux_shadowed_force_masks_storage_err;
  logic ctrl_aux_shadowed_force_masks_update_err;
  logic ctrl_aux_regwen_we;
  logic ctrl_aux_regwen_qs;
  logic ctrl_aux_regwen_wd;
  logic trigger_we;
  logic trigger_start_wd;
  logic trigger_key_iv_data_in_clear_wd;
  logic trigger_data_out_clear_wd;
  logic trigger_prng_reseed_wd;
  logic status_idle_qs;
  logic status_stall_qs;
  logic status_output_lost_qs;
  logic status_output_valid_qs;
  logic status_input_ready_qs;
  logic status_alert_recov_ctrl_update_err_qs;
  logic status_alert_fatal_fault_qs;

  // Register instances
  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[recov_ctrl_update_err]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov_ctrl_update_err (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_ctrl_update_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.recov_ctrl_update_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov_ctrl_update_err.qe = alert_test_qe;

  //   F[fatal_fault]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal_fault (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_fault_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.fatal_fault.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal_fault.qe = alert_test_qe;


  // Subregister 0 of Multireg key_share0
  // R[key_share0_0]: V(True)
  logic key_share0_0_qe;
  logic [0:0] key_share0_0_flds_we;
  assign key_share0_0_qe = &key_share0_0_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_0 (
    .re     (1'b0),
    .we     (key_share0_0_we),
    .wd     (key_share0_0_wd),
    .d      (hw2reg.key_share0[0].d),
    .qre    (),
    .qe     (key_share0_0_flds_we[0]),
    .q      (reg2hw.key_share0[0].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[0].qe = key_share0_0_qe;


  // Subregister 1 of Multireg key_share0
  // R[key_share0_1]: V(True)
  logic key_share0_1_qe;
  logic [0:0] key_share0_1_flds_we;
  assign key_share0_1_qe = &key_share0_1_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_1 (
    .re     (1'b0),
    .we     (key_share0_1_we),
    .wd     (key_share0_1_wd),
    .d      (hw2reg.key_share0[1].d),
    .qre    (),
    .qe     (key_share0_1_flds_we[0]),
    .q      (reg2hw.key_share0[1].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[1].qe = key_share0_1_qe;


  // Subregister 2 of Multireg key_share0
  // R[key_share0_2]: V(True)
  logic key_share0_2_qe;
  logic [0:0] key_share0_2_flds_we;
  assign key_share0_2_qe = &key_share0_2_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_2 (
    .re     (1'b0),
    .we     (key_share0_2_we),
    .wd     (key_share0_2_wd),
    .d      (hw2reg.key_share0[2].d),
    .qre    (),
    .qe     (key_share0_2_flds_we[0]),
    .q      (reg2hw.key_share0[2].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[2].qe = key_share0_2_qe;


  // Subregister 3 of Multireg key_share0
  // R[key_share0_3]: V(True)
  logic key_share0_3_qe;
  logic [0:0] key_share0_3_flds_we;
  assign key_share0_3_qe = &key_share0_3_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_3 (
    .re     (1'b0),
    .we     (key_share0_3_we),
    .wd     (key_share0_3_wd),
    .d      (hw2reg.key_share0[3].d),
    .qre    (),
    .qe     (key_share0_3_flds_we[0]),
    .q      (reg2hw.key_share0[3].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[3].qe = key_share0_3_qe;


  // Subregister 4 of Multireg key_share0
  // R[key_share0_4]: V(True)
  logic key_share0_4_qe;
  logic [0:0] key_share0_4_flds_we;
  assign key_share0_4_qe = &key_share0_4_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_4 (
    .re     (1'b0),
    .we     (key_share0_4_we),
    .wd     (key_share0_4_wd),
    .d      (hw2reg.key_share0[4].d),
    .qre    (),
    .qe     (key_share0_4_flds_we[0]),
    .q      (reg2hw.key_share0[4].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[4].qe = key_share0_4_qe;


  // Subregister 5 of Multireg key_share0
  // R[key_share0_5]: V(True)
  logic key_share0_5_qe;
  logic [0:0] key_share0_5_flds_we;
  assign key_share0_5_qe = &key_share0_5_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_5 (
    .re     (1'b0),
    .we     (key_share0_5_we),
    .wd     (key_share0_5_wd),
    .d      (hw2reg.key_share0[5].d),
    .qre    (),
    .qe     (key_share0_5_flds_we[0]),
    .q      (reg2hw.key_share0[5].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[5].qe = key_share0_5_qe;


  // Subregister 6 of Multireg key_share0
  // R[key_share0_6]: V(True)
  logic key_share0_6_qe;
  logic [0:0] key_share0_6_flds_we;
  assign key_share0_6_qe = &key_share0_6_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_6 (
    .re     (1'b0),
    .we     (key_share0_6_we),
    .wd     (key_share0_6_wd),
    .d      (hw2reg.key_share0[6].d),
    .qre    (),
    .qe     (key_share0_6_flds_we[0]),
    .q      (reg2hw.key_share0[6].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[6].qe = key_share0_6_qe;


  // Subregister 7 of Multireg key_share0
  // R[key_share0_7]: V(True)
  logic key_share0_7_qe;
  logic [0:0] key_share0_7_flds_we;
  assign key_share0_7_qe = &key_share0_7_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_7 (
    .re     (1'b0),
    .we     (key_share0_7_we),
    .wd     (key_share0_7_wd),
    .d      (hw2reg.key_share0[7].d),
    .qre    (),
    .qe     (key_share0_7_flds_we[0]),
    .q      (reg2hw.key_share0[7].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[7].qe = key_share0_7_qe;


  // Subregister 0 of Multireg key_share1
  // R[key_share1_0]: V(True)
  logic key_share1_0_qe;
  logic [0:0] key_share1_0_flds_we;
  assign key_share1_0_qe = &key_share1_0_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_0 (
    .re     (1'b0),
    .we     (key_share1_0_we),
    .wd     (key_share1_0_wd),
    .d      (hw2reg.key_share1[0].d),
    .qre    (),
    .qe     (key_share1_0_flds_we[0]),
    .q      (reg2hw.key_share1[0].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[0].qe = key_share1_0_qe;


  // Subregister 1 of Multireg key_share1
  // R[key_share1_1]: V(True)
  logic key_share1_1_qe;
  logic [0:0] key_share1_1_flds_we;
  assign key_share1_1_qe = &key_share1_1_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_1 (
    .re     (1'b0),
    .we     (key_share1_1_we),
    .wd     (key_share1_1_wd),
    .d      (hw2reg.key_share1[1].d),
    .qre    (),
    .qe     (key_share1_1_flds_we[0]),
    .q      (reg2hw.key_share1[1].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[1].qe = key_share1_1_qe;


  // Subregister 2 of Multireg key_share1
  // R[key_share1_2]: V(True)
  logic key_share1_2_qe;
  logic [0:0] key_share1_2_flds_we;
  assign key_share1_2_qe = &key_share1_2_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_2 (
    .re     (1'b0),
    .we     (key_share1_2_we),
    .wd     (key_share1_2_wd),
    .d      (hw2reg.key_share1[2].d),
    .qre    (),
    .qe     (key_share1_2_flds_we[0]),
    .q      (reg2hw.key_share1[2].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[2].qe = key_share1_2_qe;


  // Subregister 3 of Multireg key_share1
  // R[key_share1_3]: V(True)
  logic key_share1_3_qe;
  logic [0:0] key_share1_3_flds_we;
  assign key_share1_3_qe = &key_share1_3_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_3 (
    .re     (1'b0),
    .we     (key_share1_3_we),
    .wd     (key_share1_3_wd),
    .d      (hw2reg.key_share1[3].d),
    .qre    (),
    .qe     (key_share1_3_flds_we[0]),
    .q      (reg2hw.key_share1[3].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[3].qe = key_share1_3_qe;


  // Subregister 4 of Multireg key_share1
  // R[key_share1_4]: V(True)
  logic key_share1_4_qe;
  logic [0:0] key_share1_4_flds_we;
  assign key_share1_4_qe = &key_share1_4_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_4 (
    .re     (1'b0),
    .we     (key_share1_4_we),
    .wd     (key_share1_4_wd),
    .d      (hw2reg.key_share1[4].d),
    .qre    (),
    .qe     (key_share1_4_flds_we[0]),
    .q      (reg2hw.key_share1[4].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[4].qe = key_share1_4_qe;


  // Subregister 5 of Multireg key_share1
  // R[key_share1_5]: V(True)
  logic key_share1_5_qe;
  logic [0:0] key_share1_5_flds_we;
  assign key_share1_5_qe = &key_share1_5_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_5 (
    .re     (1'b0),
    .we     (key_share1_5_we),
    .wd     (key_share1_5_wd),
    .d      (hw2reg.key_share1[5].d),
    .qre    (),
    .qe     (key_share1_5_flds_we[0]),
    .q      (reg2hw.key_share1[5].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[5].qe = key_share1_5_qe;


  // Subregister 6 of Multireg key_share1
  // R[key_share1_6]: V(True)
  logic key_share1_6_qe;
  logic [0:0] key_share1_6_flds_we;
  assign key_share1_6_qe = &key_share1_6_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_6 (
    .re     (1'b0),
    .we     (key_share1_6_we),
    .wd     (key_share1_6_wd),
    .d      (hw2reg.key_share1[6].d),
    .qre    (),
    .qe     (key_share1_6_flds_we[0]),
    .q      (reg2hw.key_share1[6].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[6].qe = key_share1_6_qe;


  // Subregister 7 of Multireg key_share1
  // R[key_share1_7]: V(True)
  logic key_share1_7_qe;
  logic [0:0] key_share1_7_flds_we;
  assign key_share1_7_qe = &key_share1_7_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_7 (
    .re     (1'b0),
    .we     (key_share1_7_we),
    .wd     (key_share1_7_wd),
    .d      (hw2reg.key_share1[7].d),
    .qre    (),
    .qe     (key_share1_7_flds_we[0]),
    .q      (reg2hw.key_share1[7].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[7].qe = key_share1_7_qe;


  // Subregister 0 of Multireg iv
  // R[iv_0]: V(True)
  logic iv_0_qe;
  logic [0:0] iv_0_flds_we;
  assign iv_0_qe = &iv_0_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_iv_0 (
    .re     (iv_0_re),
    .we     (iv_0_we),
    .wd     (iv_0_wd),
    .d      (hw2reg.iv[0].d),
    .qre    (),
    .qe     (iv_0_flds_we[0]),
    .q      (reg2hw.iv[0].q),
    .ds     (),
    .qs     (iv_0_qs)
  );
  assign reg2hw.iv[0].qe = iv_0_qe;


  // Subregister 1 of Multireg iv
  // R[iv_1]: V(True)
  logic iv_1_qe;
  logic [0:0] iv_1_flds_we;
  assign iv_1_qe = &iv_1_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_iv_1 (
    .re     (iv_1_re),
    .we     (iv_1_we),
    .wd     (iv_1_wd),
    .d      (hw2reg.iv[1].d),
    .qre    (),
    .qe     (iv_1_flds_we[0]),
    .q      (reg2hw.iv[1].q),
    .ds     (),
    .qs     (iv_1_qs)
  );
  assign reg2hw.iv[1].qe = iv_1_qe;


  // Subregister 2 of Multireg iv
  // R[iv_2]: V(True)
  logic iv_2_qe;
  logic [0:0] iv_2_flds_we;
  assign iv_2_qe = &iv_2_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_iv_2 (
    .re     (iv_2_re),
    .we     (iv_2_we),
    .wd     (iv_2_wd),
    .d      (hw2reg.iv[2].d),
    .qre    (),
    .qe     (iv_2_flds_we[0]),
    .q      (reg2hw.iv[2].q),
    .ds     (),
    .qs     (iv_2_qs)
  );
  assign reg2hw.iv[2].qe = iv_2_qe;


  // Subregister 3 of Multireg iv
  // R[iv_3]: V(True)
  logic iv_3_qe;
  logic [0:0] iv_3_flds_we;
  assign iv_3_qe = &iv_3_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_iv_3 (
    .re     (iv_3_re),
    .we     (iv_3_we),
    .wd     (iv_3_wd),
    .d      (hw2reg.iv[3].d),
    .qre    (),
    .qe     (iv_3_flds_we[0]),
    .q      (reg2hw.iv[3].q),
    .ds     (),
    .qs     (iv_3_qs)
  );
  assign reg2hw.iv[3].qe = iv_3_qe;


  // Subregister 0 of Multireg data_in
  // R[data_in_0]: V(False)
  logic data_in_0_qe;
  logic [0:0] data_in_0_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_0_flds_we),
    .q_o(data_in_0_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (32'h0)
  ) u_data_in_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_0_we),
    .wd     (data_in_0_wd),

    // from internal hardware
    .de     (hw2reg.data_in[0].de),
    .d      (hw2reg.data_in[0].d),

    // to internal hardware
    .qe     (data_in_0_flds_we[0]),
    .q      (reg2hw.data_in[0].q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );
  assign reg2hw.data_in[0].qe = data_in_0_qe;


  // Subregister 1 of Multireg data_in
  // R[data_in_1]: V(False)
  logic data_in_1_qe;
  logic [0:0] data_in_1_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in1_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_1_flds_we),
    .q_o(data_in_1_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (32'h0)
  ) u_data_in_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_1_we),
    .wd     (data_in_1_wd),

    // from internal hardware
    .de     (hw2reg.data_in[1].de),
    .d      (hw2reg.data_in[1].d),

    // to internal hardware
    .qe     (data_in_1_flds_we[0]),
    .q      (reg2hw.data_in[1].q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );
  assign reg2hw.data_in[1].qe = data_in_1_qe;


  // Subregister 2 of Multireg data_in
  // R[data_in_2]: V(False)
  logic data_in_2_qe;
  logic [0:0] data_in_2_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in2_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_2_flds_we),
    .q_o(data_in_2_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (32'h0)
  ) u_data_in_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_2_we),
    .wd     (data_in_2_wd),

    // from internal hardware
    .de     (hw2reg.data_in[2].de),
    .d      (hw2reg.data_in[2].d),

    // to internal hardware
    .qe     (data_in_2_flds_we[0]),
    .q      (reg2hw.data_in[2].q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );
  assign reg2hw.data_in[2].qe = data_in_2_qe;


  // Subregister 3 of Multireg data_in
  // R[data_in_3]: V(False)
  logic data_in_3_qe;
  logic [0:0] data_in_3_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in3_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_3_flds_we),
    .q_o(data_in_3_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (32'h0)
  ) u_data_in_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_3_we),
    .wd     (data_in_3_wd),

    // from internal hardware
    .de     (hw2reg.data_in[3].de),
    .d      (hw2reg.data_in[3].d),

    // to internal hardware
    .qe     (data_in_3_flds_we[0]),
    .q      (reg2hw.data_in[3].q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );
  assign reg2hw.data_in[3].qe = data_in_3_qe;


  // Subregister 0 of Multireg data_out
  // R[data_out_0]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_data_out_0 (
    .re     (data_out_0_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.data_out[0].d),
    .qre    (reg2hw.data_out[0].re),
    .qe     (),
    .q      (reg2hw.data_out[0].q),
    .ds     (),
    .qs     (data_out_0_qs)
  );


  // Subregister 1 of Multireg data_out
  // R[data_out_1]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_data_out_1 (
    .re     (data_out_1_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.data_out[1].d),
    .qre    (reg2hw.data_out[1].re),
    .qe     (),
    .q      (reg2hw.data_out[1].q),
    .ds     (),
    .qs     (data_out_1_qs)
  );


  // Subregister 2 of Multireg data_out
  // R[data_out_2]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_data_out_2 (
    .re     (data_out_2_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.data_out[2].d),
    .qre    (reg2hw.data_out[2].re),
    .qe     (),
    .q      (reg2hw.data_out[2].q),
    .ds     (),
    .qs     (data_out_2_qs)
  );


  // Subregister 3 of Multireg data_out
  // R[data_out_3]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_data_out_3 (
    .re     (data_out_3_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.data_out[3].d),
    .qre    (reg2hw.data_out[3].re),
    .qe     (),
    .q      (reg2hw.data_out[3].q),
    .ds     (),
    .qs     (data_out_3_qs)
  );


  // R[ctrl_shadowed]: V(True)
  logic ctrl_shadowed_qe;
  logic [5:0] ctrl_shadowed_flds_we;
  assign ctrl_shadowed_qe = &ctrl_shadowed_flds_we;
  //   F[operation]: 1:0
  prim_subreg_ext #(
    .DW    (2)
  ) u_ctrl_shadowed_operation (
    .re     (ctrl_shadowed_re),
    .we     (ctrl_shadowed_we),
    .wd     (ctrl_shadowed_operation_wd),
    .d      (hw2reg.ctrl_shadowed.operation.d),
    .qre    (reg2hw.ctrl_shadowed.operation.re),
    .qe     (ctrl_shadowed_flds_we[0]),
    .q      (reg2hw.ctrl_shadowed.operation.q),
    .ds     (),
    .qs     (ctrl_shadowed_operation_qs)
  );
  assign reg2hw.ctrl_shadowed.operation.qe = ctrl_shadowed_qe;

  //   F[mode]: 7:2
  prim_subreg_ext #(
    .DW    (6)
  ) u_ctrl_shadowed_mode (
    .re     (ctrl_shadowed_re),
    .we     (ctrl_shadowed_we),
    .wd     (ctrl_shadowed_mode_wd),
    .d      (hw2reg.ctrl_shadowed.mode.d),
    .qre    (reg2hw.ctrl_shadowed.mode.re),
    .qe     (ctrl_shadowed_flds_we[1]),
    .q      (reg2hw.ctrl_shadowed.mode.q),
    .ds     (),
    .qs     (ctrl_shadowed_mode_qs)
  );
  assign reg2hw.ctrl_shadowed.mode.qe = ctrl_shadowed_qe;

  //   F[key_len]: 10:8
  prim_subreg_ext #(
    .DW    (3)
  ) u_ctrl_shadowed_key_len (
    .re     (ctrl_shadowed_re),
    .we     (ctrl_shadowed_we),
    .wd     (ctrl_shadowed_key_len_wd),
    .d      (hw2reg.ctrl_shadowed.key_len.d),
    .qre    (reg2hw.ctrl_shadowed.key_len.re),
    .qe     (ctrl_shadowed_flds_we[2]),
    .q      (reg2hw.ctrl_shadowed.key_len.q),
    .ds     (),
    .qs     (ctrl_shadowed_key_len_qs)
  );
  assign reg2hw.ctrl_shadowed.key_len.qe = ctrl_shadowed_qe;

  //   F[sideload]: 11:11
  prim_subreg_ext #(
    .DW    (1)
  ) u_ctrl_shadowed_sideload (
    .re     (ctrl_shadowed_re),
    .we     (ctrl_shadowed_we),
    .wd     (ctrl_shadowed_sideload_wd),
    .d      (hw2reg.ctrl_shadowed.sideload.d),
    .qre    (reg2hw.ctrl_shadowed.sideload.re),
    .qe     (ctrl_shadowed_flds_we[3]),
    .q      (reg2hw.ctrl_shadowed.sideload.q),
    .ds     (),
    .qs     (ctrl_shadowed_sideload_qs)
  );
  assign reg2hw.ctrl_shadowed.sideload.qe = ctrl_shadowed_qe;

  //   F[prng_reseed_rate]: 14:12
  prim_subreg_ext #(
    .DW    (3)
  ) u_ctrl_shadowed_prng_reseed_rate (
    .re     (ctrl_shadowed_re),
    .we     (ctrl_shadowed_we),
    .wd     (ctrl_shadowed_prng_reseed_rate_wd),
    .d      (hw2reg.ctrl_shadowed.prng_reseed_rate.d),
    .qre    (reg2hw.ctrl_shadowed.prng_reseed_rate.re),
    .qe     (ctrl_shadowed_flds_we[4]),
    .q      (reg2hw.ctrl_shadowed.prng_reseed_rate.q),
    .ds     (),
    .qs     (ctrl_shadowed_prng_reseed_rate_qs)
  );
  assign reg2hw.ctrl_shadowed.prng_reseed_rate.qe = ctrl_shadowed_qe;

  //   F[manual_operation]: 15:15
  prim_subreg_ext #(
    .DW    (1)
  ) u_ctrl_shadowed_manual_operation (
    .re     (ctrl_shadowed_re),
    .we     (ctrl_shadowed_we),
    .wd     (ctrl_shadowed_manual_operation_wd),
    .d      (hw2reg.ctrl_shadowed.manual_operation.d),
    .qre    (reg2hw.ctrl_shadowed.manual_operation.re),
    .qe     (ctrl_shadowed_flds_we[5]),
    .q      (reg2hw.ctrl_shadowed.manual_operation.q),
    .ds     (),
    .qs     (ctrl_shadowed_manual_operation_qs)
  );
  assign reg2hw.ctrl_shadowed.manual_operation.qe = ctrl_shadowed_qe;


  // R[ctrl_aux_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic ctrl_aux_shadowed_gated_we;
  assign ctrl_aux_shadowed_gated_we = ctrl_aux_shadowed_we & ctrl_aux_regwen_qs;
  //   F[key_touch_forces_reseed]: 0:0
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h1)
  ) u_ctrl_aux_shadowed_key_touch_forces_reseed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (ctrl_aux_shadowed_re),
    .we     (ctrl_aux_shadowed_gated_we),
    .wd     (ctrl_aux_shadowed_key_touch_forces_reseed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl_aux_shadowed.key_touch_forces_reseed.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_aux_shadowed_key_touch_forces_reseed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (ctrl_aux_shadowed_key_touch_forces_reseed_update_err),
    .err_storage (ctrl_aux_shadowed_key_touch_forces_reseed_storage_err)
  );

  //   F[force_masks]: 1:1
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_aux_shadowed_force_masks (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (ctrl_aux_shadowed_re),
    .we     (ctrl_aux_shadowed_gated_we),
    .wd     (ctrl_aux_shadowed_force_masks_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl_aux_shadowed.force_masks.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_aux_shadowed_force_masks_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (ctrl_aux_shadowed_force_masks_update_err),
    .err_storage (ctrl_aux_shadowed_force_masks_storage_err)
  );


  // R[ctrl_aux_regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_ctrl_aux_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_aux_regwen_we),
    .wd     (ctrl_aux_regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_aux_regwen_qs)
  );


  // R[trigger]: V(False)
  //   F[start]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (1'h0)
  ) u_trigger_start (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (trigger_we),
    .wd     (trigger_start_wd),

    // from internal hardware
    .de     (hw2reg.trigger.start.de),
    .d      (hw2reg.trigger.start.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.trigger.start.q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );

  //   F[key_iv_data_in_clear]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (1'h1)
  ) u_trigger_key_iv_data_in_clear (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (trigger_we),
    .wd     (trigger_key_iv_data_in_clear_wd),

    // from internal hardware
    .de     (hw2reg.trigger.key_iv_data_in_clear.de),
    .d      (hw2reg.trigger.key_iv_data_in_clear.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.trigger.key_iv_data_in_clear.q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );

  //   F[data_out_clear]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (1'h1)
  ) u_trigger_data_out_clear (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (trigger_we),
    .wd     (trigger_data_out_clear_wd),

    // from internal hardware
    .de     (hw2reg.trigger.data_out_clear.de),
    .d      (hw2reg.trigger.data_out_clear.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.trigger.data_out_clear.q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );

  //   F[prng_reseed]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (1'h1)
  ) u_trigger_prng_reseed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (trigger_we),
    .wd     (trigger_prng_reseed_wd),

    // from internal hardware
    .de     (hw2reg.trigger.prng_reseed.de),
    .d      (hw2reg.trigger.prng_reseed.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.trigger.prng_reseed.q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );


  // R[status]: V(False)
  //   F[idle]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_idle (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.idle.de),
    .d      (hw2reg.status.idle.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.status.idle.q),
    .ds     (),

    // to register interface (read)
    .qs     (status_idle_qs)
  );

  //   F[stall]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_stall (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.stall.de),
    .d      (hw2reg.status.stall.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (status_stall_qs)
  );

  //   F[output_lost]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_output_lost (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.output_lost.de),
    .d      (hw2reg.status.output_lost.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.status.output_lost.q),
    .ds     (),

    // to register interface (read)
    .qs     (status_output_lost_qs)
  );

  //   F[output_valid]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_output_valid (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.output_valid.de),
    .d      (hw2reg.status.output_valid.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (status_output_valid_qs)
  );

  //   F[input_ready]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_input_ready (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.input_ready.de),
    .d      (hw2reg.status.input_ready.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (status_input_ready_qs)
  );

  //   F[alert_recov_ctrl_update_err]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_alert_recov_ctrl_update_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.alert_recov_ctrl_update_err.de),
    .d      (hw2reg.status.alert_recov_ctrl_update_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (status_alert_recov_ctrl_update_err_qs)
  );

  //   F[alert_fatal_fault]: 6:6
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_status_alert_fatal_fault (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.alert_fatal_fault.de),
    .d      (hw2reg.status.alert_fatal_fault.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (status_alert_fatal_fault_qs)
  );



  logic [33:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == AES_ALERT_TEST_OFFSET);
    addr_hit[ 1] = (reg_addr == AES_KEY_SHARE0_0_OFFSET);
    addr_hit[ 2] = (reg_addr == AES_KEY_SHARE0_1_OFFSET);
    addr_hit[ 3] = (reg_addr == AES_KEY_SHARE0_2_OFFSET);
    addr_hit[ 4] = (reg_addr == AES_KEY_SHARE0_3_OFFSET);
    addr_hit[ 5] = (reg_addr == AES_KEY_SHARE0_4_OFFSET);
    addr_hit[ 6] = (reg_addr == AES_KEY_SHARE0_5_OFFSET);
    addr_hit[ 7] = (reg_addr == AES_KEY_SHARE0_6_OFFSET);
    addr_hit[ 8] = (reg_addr == AES_KEY_SHARE0_7_OFFSET);
    addr_hit[ 9] = (reg_addr == AES_KEY_SHARE1_0_OFFSET);
    addr_hit[10] = (reg_addr == AES_KEY_SHARE1_1_OFFSET);
    addr_hit[11] = (reg_addr == AES_KEY_SHARE1_2_OFFSET);
    addr_hit[12] = (reg_addr == AES_KEY_SHARE1_3_OFFSET);
    addr_hit[13] = (reg_addr == AES_KEY_SHARE1_4_OFFSET);
    addr_hit[14] = (reg_addr == AES_KEY_SHARE1_5_OFFSET);
    addr_hit[15] = (reg_addr == AES_KEY_SHARE1_6_OFFSET);
    addr_hit[16] = (reg_addr == AES_KEY_SHARE1_7_OFFSET);
    addr_hit[17] = (reg_addr == AES_IV_0_OFFSET);
    addr_hit[18] = (reg_addr == AES_IV_1_OFFSET);
    addr_hit[19] = (reg_addr == AES_IV_2_OFFSET);
    addr_hit[20] = (reg_addr == AES_IV_3_OFFSET);
    addr_hit[21] = (reg_addr == AES_DATA_IN_0_OFFSET);
    addr_hit[22] = (reg_addr == AES_DATA_IN_1_OFFSET);
    addr_hit[23] = (reg_addr == AES_DATA_IN_2_OFFSET);
    addr_hit[24] = (reg_addr == AES_DATA_IN_3_OFFSET);
    addr_hit[25] = (reg_addr == AES_DATA_OUT_0_OFFSET);
    addr_hit[26] = (reg_addr == AES_DATA_OUT_1_OFFSET);
    addr_hit[27] = (reg_addr == AES_DATA_OUT_2_OFFSET);
    addr_hit[28] = (reg_addr == AES_DATA_OUT_3_OFFSET);
    addr_hit[29] = (reg_addr == AES_CTRL_SHADOWED_OFFSET);
    addr_hit[30] = (reg_addr == AES_CTRL_AUX_SHADOWED_OFFSET);
    addr_hit[31] = (reg_addr == AES_CTRL_AUX_REGWEN_OFFSET);
    addr_hit[32] = (reg_addr == AES_TRIGGER_OFFSET);
    addr_hit[33] = (reg_addr == AES_STATUS_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(AES_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(AES_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(AES_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(AES_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(AES_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(AES_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(AES_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(AES_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(AES_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(AES_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(AES_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(AES_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(AES_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(AES_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(AES_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(AES_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(AES_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(AES_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(AES_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(AES_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(AES_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(AES_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(AES_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(AES_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(AES_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(AES_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(AES_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(AES_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(AES_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(AES_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(AES_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(AES_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(AES_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(AES_PERMIT[33] & ~reg_be)))));
  end

  // Generate write-enables
  assign alert_test_we = addr_hit[0] & reg_we & !reg_error;

  assign alert_test_recov_ctrl_update_err_wd = reg_wdata[0];

  assign alert_test_fatal_fault_wd = reg_wdata[1];
  assign key_share0_0_we = addr_hit[1] & reg_we & !reg_error;

  assign key_share0_0_wd = reg_wdata[31:0];
  assign key_share0_1_we = addr_hit[2] & reg_we & !reg_error;

  assign key_share0_1_wd = reg_wdata[31:0];
  assign key_share0_2_we = addr_hit[3] & reg_we & !reg_error;

  assign key_share0_2_wd = reg_wdata[31:0];
  assign key_share0_3_we = addr_hit[4] & reg_we & !reg_error;

  assign key_share0_3_wd = reg_wdata[31:0];
  assign key_share0_4_we = addr_hit[5] & reg_we & !reg_error;

  assign key_share0_4_wd = reg_wdata[31:0];
  assign key_share0_5_we = addr_hit[6] & reg_we & !reg_error;

  assign key_share0_5_wd = reg_wdata[31:0];
  assign key_share0_6_we = addr_hit[7] & reg_we & !reg_error;

  assign key_share0_6_wd = reg_wdata[31:0];
  assign key_share0_7_we = addr_hit[8] & reg_we & !reg_error;

  assign key_share0_7_wd = reg_wdata[31:0];
  assign key_share1_0_we = addr_hit[9] & reg_we & !reg_error;

  assign key_share1_0_wd = reg_wdata[31:0];
  assign key_share1_1_we = addr_hit[10] & reg_we & !reg_error;

  assign key_share1_1_wd = reg_wdata[31:0];
  assign key_share1_2_we = addr_hit[11] & reg_we & !reg_error;

  assign key_share1_2_wd = reg_wdata[31:0];
  assign key_share1_3_we = addr_hit[12] & reg_we & !reg_error;

  assign key_share1_3_wd = reg_wdata[31:0];
  assign key_share1_4_we = addr_hit[13] & reg_we & !reg_error;

  assign key_share1_4_wd = reg_wdata[31:0];
  assign key_share1_5_we = addr_hit[14] & reg_we & !reg_error;

  assign key_share1_5_wd = reg_wdata[31:0];
  assign key_share1_6_we = addr_hit[15] & reg_we & !reg_error;

  assign key_share1_6_wd = reg_wdata[31:0];
  assign key_share1_7_we = addr_hit[16] & reg_we & !reg_error;

  assign key_share1_7_wd = reg_wdata[31:0];
  assign iv_0_re = addr_hit[17] & reg_re & !reg_error;
  assign iv_0_we = addr_hit[17] & reg_we & !reg_error;

  assign iv_0_wd = reg_wdata[31:0];
  assign iv_1_re = addr_hit[18] & reg_re & !reg_error;
  assign iv_1_we = addr_hit[18] & reg_we & !reg_error;

  assign iv_1_wd = reg_wdata[31:0];
  assign iv_2_re = addr_hit[19] & reg_re & !reg_error;
  assign iv_2_we = addr_hit[19] & reg_we & !reg_error;

  assign iv_2_wd = reg_wdata[31:0];
  assign iv_3_re = addr_hit[20] & reg_re & !reg_error;
  assign iv_3_we = addr_hit[20] & reg_we & !reg_error;

  assign iv_3_wd = reg_wdata[31:0];
  assign data_in_0_we = addr_hit[21] & reg_we & !reg_error;

  assign data_in_0_wd = reg_wdata[31:0];
  assign data_in_1_we = addr_hit[22] & reg_we & !reg_error;

  assign data_in_1_wd = reg_wdata[31:0];
  assign data_in_2_we = addr_hit[23] & reg_we & !reg_error;

  assign data_in_2_wd = reg_wdata[31:0];
  assign data_in_3_we = addr_hit[24] & reg_we & !reg_error;

  assign data_in_3_wd = reg_wdata[31:0];
  assign data_out_0_re = addr_hit[25] & reg_re & !reg_error;
  assign data_out_1_re = addr_hit[26] & reg_re & !reg_error;
  assign data_out_2_re = addr_hit[27] & reg_re & !reg_error;
  assign data_out_3_re = addr_hit[28] & reg_re & !reg_error;
  assign ctrl_shadowed_re = addr_hit[29] & reg_re & !reg_error;
  assign ctrl_shadowed_we = addr_hit[29] & reg_we & !reg_error;

  assign ctrl_shadowed_operation_wd = reg_wdata[1:0];

  assign ctrl_shadowed_mode_wd = reg_wdata[7:2];

  assign ctrl_shadowed_key_len_wd = reg_wdata[10:8];

  assign ctrl_shadowed_sideload_wd = reg_wdata[11];

  assign ctrl_shadowed_prng_reseed_rate_wd = reg_wdata[14:12];

  assign ctrl_shadowed_manual_operation_wd = reg_wdata[15];
  assign ctrl_aux_shadowed_re = addr_hit[30] & reg_re & !reg_error;
  assign ctrl_aux_shadowed_we = addr_hit[30] & reg_we & !reg_error;

  assign ctrl_aux_shadowed_key_touch_forces_reseed_wd = reg_wdata[0];

  assign ctrl_aux_shadowed_force_masks_wd = reg_wdata[1];
  assign ctrl_aux_regwen_we = addr_hit[31] & reg_we & !reg_error;

  assign ctrl_aux_regwen_wd = reg_wdata[0];
  assign trigger_we = addr_hit[32] & reg_we & !reg_error;

  assign trigger_start_wd = reg_wdata[0];

  assign trigger_key_iv_data_in_clear_wd = reg_wdata[1];

  assign trigger_data_out_clear_wd = reg_wdata[2];

  assign trigger_prng_reseed_wd = reg_wdata[3];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = alert_test_we;
    reg_we_check[1] = key_share0_0_we;
    reg_we_check[2] = key_share0_1_we;
    reg_we_check[3] = key_share0_2_we;
    reg_we_check[4] = key_share0_3_we;
    reg_we_check[5] = key_share0_4_we;
    reg_we_check[6] = key_share0_5_we;
    reg_we_check[7] = key_share0_6_we;
    reg_we_check[8] = key_share0_7_we;
    reg_we_check[9] = key_share1_0_we;
    reg_we_check[10] = key_share1_1_we;
    reg_we_check[11] = key_share1_2_we;
    reg_we_check[12] = key_share1_3_we;
    reg_we_check[13] = key_share1_4_we;
    reg_we_check[14] = key_share1_5_we;
    reg_we_check[15] = key_share1_6_we;
    reg_we_check[16] = key_share1_7_we;
    reg_we_check[17] = iv_0_we;
    reg_we_check[18] = iv_1_we;
    reg_we_check[19] = iv_2_we;
    reg_we_check[20] = iv_3_we;
    reg_we_check[21] = data_in_0_we;
    reg_we_check[22] = data_in_1_we;
    reg_we_check[23] = data_in_2_we;
    reg_we_check[24] = data_in_3_we;
    reg_we_check[25] = 1'b0;
    reg_we_check[26] = 1'b0;
    reg_we_check[27] = 1'b0;
    reg_we_check[28] = 1'b0;
    reg_we_check[29] = ctrl_shadowed_we;
    reg_we_check[30] = ctrl_aux_shadowed_gated_we;
    reg_we_check[31] = ctrl_aux_regwen_we;
    reg_we_check[32] = trigger_we;
    reg_we_check[33] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[1]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = iv_0_qs;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = iv_1_qs;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = iv_2_qs;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = iv_3_qs;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = data_out_0_qs;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = data_out_1_qs;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = data_out_2_qs;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = data_out_3_qs;
      end

      addr_hit[29]: begin
        reg_rdata_next[1:0] = ctrl_shadowed_operation_qs;
        reg_rdata_next[7:2] = ctrl_shadowed_mode_qs;
        reg_rdata_next[10:8] = ctrl_shadowed_key_len_qs;
        reg_rdata_next[11] = ctrl_shadowed_sideload_qs;
        reg_rdata_next[14:12] = ctrl_shadowed_prng_reseed_rate_qs;
        reg_rdata_next[15] = ctrl_shadowed_manual_operation_qs;
      end

      addr_hit[30]: begin
        reg_rdata_next[0] = ctrl_aux_shadowed_key_touch_forces_reseed_qs;
        reg_rdata_next[1] = ctrl_aux_shadowed_force_masks_qs;
      end

      addr_hit[31]: begin
        reg_rdata_next[0] = ctrl_aux_regwen_qs;
      end

      addr_hit[32]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
        reg_rdata_next[2] = '0;
        reg_rdata_next[3] = '0;
      end

      addr_hit[33]: begin
        reg_rdata_next[0] = status_idle_qs;
        reg_rdata_next[1] = status_stall_qs;
        reg_rdata_next[2] = status_output_lost_qs;
        reg_rdata_next[3] = status_output_valid_qs;
        reg_rdata_next[4] = status_input_ready_qs;
        reg_rdata_next[5] = status_alert_recov_ctrl_update_err_qs;
        reg_rdata_next[6] = status_alert_fatal_fault_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  logic rst_done;
  logic shadow_rst_done;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rst_done <= '0;
    end else begin
      rst_done <= 1'b1;
    end
  end

  always_ff @(posedge clk_i or negedge rst_shadowed_ni) begin
    if (!rst_shadowed_ni) begin
      shadow_rst_done <= '0;
    end else begin
      shadow_rst_done <= 1'b1;
    end
  end

  // both shadow and normal resets have been released
  assign shadow_busy = ~(rst_done & shadow_rst_done);

  // Collect up storage and update errors
  assign shadowed_storage_err_o = |{
    ctrl_aux_shadowed_key_touch_forces_reseed_storage_err,
    ctrl_aux_shadowed_force_masks_storage_err
  };
  assign shadowed_update_err_o = |{
    ctrl_aux_shadowed_key_touch_forces_reseed_update_err,
    ctrl_aux_shadowed_force_masks_update_err
  };

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES shadowed control register
//
// This module implements the AES shadowed control register. The main differences compared
// to implementing the register as part of the auto-generated aes_reg_top.sv are:
//
// 1. The hardware can block updates to the control register from software.
//    Whenever the module is busy, control register writes are ignored.
// 2. Invalid values written by software are resolved to valid configurations.

`include "prim_assert.sv"

module aes_ctrl_reg_shadowed
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit AES192Enable = 1
) (
  input  logic clk_i,
  input  logic rst_ni,
  input  logic rst_shadowed_ni,
  // Main control
  output logic      qe_o, // software wants to write
  input  logic      we_i, // hardware grants software write
  output logic      phase_o,
  output aes_op_e   operation_o,
  output aes_mode_e mode_o,
  output key_len_e  key_len_o,
  output logic      sideload_o,
  output prs_rate_e prng_reseed_rate_o,
  output logic      manual_operation_o,

  // Alerts
  output logic err_update_o,
  output logic err_storage_o,

  // Bus interface
  input  aes_reg2hw_ctrl_shadowed_reg_t reg2hw_ctrl_i,
  output aes_hw2reg_ctrl_shadowed_reg_t hw2reg_ctrl_o
);

  // Signals
  ctrl_reg_t ctrl_wd;
  aes_op_e   op;
  aes_mode_e mode;
  key_len_e  key_len;
  prs_rate_e prng_reseed_rate;
  logic      phase_operation;
  logic      phase_mode;
  logic      phase_key_len;
  logic      phase_key_sideload;
  logic      phase_prng_reseed_rate;
  logic      phase_manual_operation;
  logic      err_update_operation;
  logic      err_update_mode;
  logic      err_update_key_len;
  logic      err_update_sideload;
  logic      err_update_prng_reseed_rate;
  logic      err_update_manual_operation;
  logic      err_storage_operation;
  logic      err_storage_mode;
  logic      err_storage_key_len;
  logic      err_storage_sideload;
  logic      err_storage_prng_reseed_rate;
  logic      err_storage_manual_operation;

  // Get and forward write enable. Writes are only allowed if the module is idle.
  assign qe_o = reg2hw_ctrl_i.operation.qe & reg2hw_ctrl_i.mode.qe &
      reg2hw_ctrl_i.key_len.qe & reg2hw_ctrl_i.sideload.qe &
      reg2hw_ctrl_i.prng_reseed_rate.qe & reg2hw_ctrl_i.manual_operation.qe;

  // Get and resolve values from register interface.
  assign op = aes_op_e'(reg2hw_ctrl_i.operation.q);
  always_comb begin : operation_get
    unique case (op)
      AES_ENC: ctrl_wd.operation = AES_ENC;
      AES_DEC: ctrl_wd.operation = AES_DEC;
      default: ctrl_wd.operation = AES_ENC; // unsupported values are mapped to AES_ENC
    endcase
  end

  assign mode = aes_mode_e'(reg2hw_ctrl_i.mode.q);
  always_comb begin : mode_get
    unique case (mode)
      AES_ECB: ctrl_wd.mode = AES_ECB;
      AES_CBC: ctrl_wd.mode = AES_CBC;
      AES_CFB: ctrl_wd.mode = AES_CFB;
      AES_OFB: ctrl_wd.mode = AES_OFB;
      AES_CTR: ctrl_wd.mode = AES_CTR;
      default: ctrl_wd.mode = AES_NONE; // unsupported values are mapped to AES_NONE
    endcase
  end

  assign key_len = key_len_e'(reg2hw_ctrl_i.key_len.q);
  always_comb begin : key_len_get
    unique case (key_len)
      AES_128: ctrl_wd.key_len = AES_128;
      AES_256: ctrl_wd.key_len = AES_256;
      AES_192: ctrl_wd.key_len = AES192Enable ? AES_192 : AES_256;
      default: ctrl_wd.key_len = AES_256; // unsupported values are mapped to AES_256
    endcase
  end

  assign ctrl_wd.sideload = reg2hw_ctrl_i.sideload.q;

  assign prng_reseed_rate = prs_rate_e'(reg2hw_ctrl_i.prng_reseed_rate.q);
  always_comb begin : prng_reseed_rate_get
    unique case (prng_reseed_rate)
      PER_1:   ctrl_wd.prng_reseed_rate = PER_1;
      PER_64:  ctrl_wd.prng_reseed_rate = PER_64;
      PER_8K:  ctrl_wd.prng_reseed_rate = PER_8K;
      default: ctrl_wd.prng_reseed_rate = PER_1; // unsupported values are mapped to PER_1.
    endcase
  end

  assign ctrl_wd.manual_operation = reg2hw_ctrl_i.manual_operation.q;

  // SEC_CM: MAIN.CONFIG.SHADOW
  // Instantiate one shadowed register primitive per field. An update error in a field should
  // only prevent the update of the affected field.
  prim_subreg_shadow #(
    .DW      ($bits(aes_op_e)),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (AES_CTRL_SHADOWED_OPERATION_RESVAL)
  ) u_ctrl_reg_shadowed_operation (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .re         (reg2hw_ctrl_i.operation.re),
    .we         (we_i),
    .wd         ({ctrl_wd.operation}),
    .de         (1'b0),
    .d          ('0),
    .qe         (),
    .q          (hw2reg_ctrl_o.operation.d),
    .qs         (),
    .ds         (),
    .phase      (phase_operation),
    .err_update (err_update_operation),
    .err_storage(err_storage_operation)
  );

  prim_subreg_shadow #(
    .DW      ($bits(aes_mode_e)),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (AES_CTRL_SHADOWED_MODE_RESVAL)
  ) u_ctrl_reg_shadowed_mode (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .re         (reg2hw_ctrl_i.mode.re),
    .we         (we_i),
    .wd         ({ctrl_wd.mode}),
    .de         (1'b0),
    .d          ('0),
    .qe         (),
    .q          (hw2reg_ctrl_o.mode.d),
    .qs         (),
    .ds         (),
    .phase      (phase_mode),
    .err_update (err_update_mode),
    .err_storage(err_storage_mode)
  );

  prim_subreg_shadow #(
    .DW      ($bits(key_len_e)),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (AES_CTRL_SHADOWED_KEY_LEN_RESVAL)
  ) u_ctrl_reg_shadowed_key_len (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .re         (reg2hw_ctrl_i.key_len.re),
    .we         (we_i),
    .wd         ({ctrl_wd.key_len}),
    .de         (1'b0),
    .d          ('0),
    .qe         (),
    .q          (hw2reg_ctrl_o.key_len.d),
    .qs         (),
    .ds         (),
    .phase      (phase_key_len),
    .err_update (err_update_key_len),
    .err_storage(err_storage_key_len)
  );

  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (AES_CTRL_SHADOWED_SIDELOAD_RESVAL)
  ) u_ctrl_reg_shadowed_sideload (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .re         (reg2hw_ctrl_i.sideload.re),
    .we         (we_i),
    .wd         (ctrl_wd.sideload),
    .de         (1'b0),
    .d          ('0),
    .qe         (),
    .q          (hw2reg_ctrl_o.sideload.d),
    .qs         (),
    .ds         (),
    .phase      (phase_key_sideload),
    .err_update (err_update_sideload),
    .err_storage(err_storage_sideload)
  );

  prim_subreg_shadow #(
    .DW      ($bits(prs_rate_e)),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (AES_CTRL_SHADOWED_PRNG_RESEED_RATE_RESVAL)
  ) u_ctrl_reg_shadowed_prng_reseed_rate (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .re         (reg2hw_ctrl_i.prng_reseed_rate.re),
    .we         (we_i),
    .wd         ({ctrl_wd.prng_reseed_rate}),
    .de         (1'b0),
    .d          ('0),
    .qe         (),
    .q          (hw2reg_ctrl_o.prng_reseed_rate.d),
    .qs         (),
    .ds         (),
    .phase      (phase_prng_reseed_rate),
    .err_update (err_update_prng_reseed_rate),
    .err_storage(err_storage_prng_reseed_rate)
  );

  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (AES_CTRL_SHADOWED_MANUAL_OPERATION_RESVAL)
  ) u_ctrl_reg_shadowed_manual_operation (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .re         (reg2hw_ctrl_i.manual_operation.re),
    .we         (we_i),
    .wd         (ctrl_wd.manual_operation),
    .de         (1'b0),
    .d          ('0),
    .qe         (),
    .q          (hw2reg_ctrl_o.manual_operation.d),
    .qs         (),
    .ds         (),
    .phase      (phase_manual_operation),
    .err_update (err_update_manual_operation),
    .err_storage(err_storage_manual_operation)
  );

  // Collect phase signals.
  assign phase_o = phase_operation | phase_mode | phase_key_len | phase_key_sideload |
      phase_prng_reseed_rate | phase_manual_operation;

  // Collect alerts.
  assign err_update_o = err_update_operation | err_update_mode | err_update_key_len |
      err_update_sideload | err_update_prng_reseed_rate | err_update_manual_operation;
  assign err_storage_o = err_storage_operation | err_storage_mode | err_storage_key_len |
      err_storage_sideload | err_storage_prng_reseed_rate | err_storage_manual_operation;

  // Generate shorter references.
  // Doing that here as opposed to in aes_core avoids several Verilator lint errors.
  assign operation_o        = aes_op_e'(hw2reg_ctrl_o.operation.d);
  assign mode_o             = aes_mode_e'(hw2reg_ctrl_o.mode.d);
  assign key_len_o          = key_len_e'(hw2reg_ctrl_o.key_len.d);
  assign sideload_o         = hw2reg_ctrl_o.sideload.d;
  assign prng_reseed_rate_o = prs_rate_e'(hw2reg_ctrl_o.prng_reseed_rate.d);
  assign manual_operation_o = hw2reg_ctrl_o.manual_operation.d;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES core implementation

`include "prim_assert.sv"

module aes_core
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          AES192Enable         = 1,
  parameter bit          SecMasking           = 1,
  parameter sbox_impl_e  SecSBoxImpl          = SBoxImplDom,
  parameter int unsigned SecStartTriggerDelay = 0,
  parameter bit          SecAllowForcingMasks = 0,
  parameter bit          SecSkipPRNGReseeding = 0,
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,

  localparam int         NumShares            = SecMasking ? 2 : 1, // derived parameter

  parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingSharePerm = RndCnstClearingSharePermDefault,
  parameter masking_lfsr_seed_t  RndCnstMaskingLfsrSeed   = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t  RndCnstMaskingLfsrPerm   = RndCnstMaskingLfsrPermDefault
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  input  logic                        rst_shadowed_ni,

  // Entropy request interfaces for clearing and masking PRNGs
  output logic                        entropy_clearing_req_o,
  input  logic                        entropy_clearing_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_clearing_i,
  output logic                        entropy_masking_req_o,
  input  logic                        entropy_masking_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_masking_i,

  // Key manager (keymgr) key sideload interface
  input  keymgr_pkg::hw_key_req_t     keymgr_key_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t         lc_escalate_en_i,

  // Alerts
  input  logic                        shadowed_storage_err_i,
  input  logic                        shadowed_update_err_i,
  input  logic                        intg_err_alert_i,
  output logic                        alert_recov_o,
  output logic                        alert_fatal_o,

  // Bus Interface
  input  aes_reg2hw_t                 reg2hw,
  output aes_hw2reg_t                 hw2reg
);

  // Signals
  logic                                       ctrl_qe;
  logic                                       ctrl_we;
  logic                                       ctrl_phase;
  aes_op_e                                    aes_op_q;
  aes_mode_e                                  aes_mode_q;
  ciph_op_e                                   cipher_op;
  ciph_op_e                                   cipher_op_buf;
  key_len_e                                   key_len_q;
  logic                                       sideload_q;
  prs_rate_e                                  prng_reseed_rate_q;
  logic                                       manual_operation_q;
  logic                                       ctrl_reg_err_update;
  logic                                       ctrl_reg_err_storage;
  logic                                       ctrl_err_update;
  logic                                       ctrl_err_storage;
  logic                                       ctrl_err_storage_d;
  logic                                       ctrl_err_storage_q;
  logic                                       ctrl_alert;
  logic                                       key_touch_forces_reseed;
  logic                                       force_masks;
  logic                                       mux_sel_err;
  logic                                       sp_enc_err_d, sp_enc_err_q;
  logic                                       clear_on_fatal;

  logic                       [3:0][3:0][7:0] state_in;
  logic                      [SISelWidth-1:0] state_in_sel_raw;
  si_sel_e                                    state_in_sel_ctrl;
  si_sel_e                                    state_in_sel;
  logic                                       state_in_sel_err;
  logic                       [3:0][3:0][7:0] add_state_in;
  logic                   [AddSISelWidth-1:0] add_state_in_sel_raw;
  add_si_sel_e                                add_state_in_sel_ctrl;
  add_si_sel_e                                add_state_in_sel;
  logic                                       add_state_in_sel_err;

  logic                       [3:0][3:0][7:0] state_mask;
  logic                       [3:0][3:0][7:0] state_init [NumShares];
  logic                       [3:0][3:0][7:0] state_done [NumShares];
  logic                       [3:0][3:0][7:0] state_out;

  logic                [NumRegsKey-1:0][31:0] key_init [NumSharesKey];
  logic                [NumRegsKey-1:0]       key_init_qe [NumSharesKey];
  logic                [NumRegsKey-1:0]       key_init_qe_buf [NumSharesKey];
  logic                [NumRegsKey-1:0][31:0] key_init_d [NumSharesKey];
  logic                [NumRegsKey-1:0][31:0] key_init_q [NumSharesKey];
  logic                [NumRegsKey-1:0][31:0] key_init_cipher [NumShares];
  sp2v_e               [NumRegsKey-1:0]       key_init_we_ctrl [NumSharesKey];
  sp2v_e               [NumRegsKey-1:0]       key_init_we [NumSharesKey];
  logic                 [KeyInitSelWidth-1:0] key_init_sel_raw;
  key_init_sel_e                              key_init_sel_ctrl;
  key_init_sel_e                              key_init_sel;
  logic                                       key_init_sel_err;
  logic                [NumRegsKey-1:0][31:0] key_sideload [NumSharesKey];

  logic                 [NumRegsIv-1:0][31:0] iv;
  logic                 [NumRegsIv-1:0]       iv_qe;
  logic                 [NumRegsIv-1:0]       iv_qe_buf;
  logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] iv_d;
  logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] iv_q;
  sp2v_e [NumSlicesCtr-1:0]                   iv_we_ctrl;
  sp2v_e [NumSlicesCtr-1:0]                   iv_we;
  logic                      [IVSelWidth-1:0] iv_sel_raw;
  iv_sel_e                                    iv_sel_ctrl;
  iv_sel_e                                    iv_sel;
  logic                                       iv_sel_err;

  logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] ctr;
  sp2v_e [NumSlicesCtr-1:0]                   ctr_we;
  sp2v_e                                      ctr_incr;
  sp2v_e                                      ctr_ready;
  logic                                       ctr_alert;

  logic               [NumRegsData-1:0][31:0] data_in_prev_d;
  logic               [NumRegsData-1:0][31:0] data_in_prev_q;
  sp2v_e                                      data_in_prev_we_ctrl;
  sp2v_e                                      data_in_prev_we;
  logic                     [DIPSelWidth-1:0] data_in_prev_sel_raw;
  dip_sel_e                                   data_in_prev_sel_ctrl;
  dip_sel_e                                   data_in_prev_sel;
  logic                                       data_in_prev_sel_err;

  logic               [NumRegsData-1:0][31:0] data_in;
  logic               [NumRegsData-1:0]       data_in_qe;
  logic               [NumRegsData-1:0]       data_in_qe_buf;
  logic                                       data_in_we;

  logic                       [3:0][3:0][7:0] add_state_out;
  logic                   [AddSOSelWidth-1:0] add_state_out_sel_raw;
  add_so_sel_e                                add_state_out_sel_ctrl;
  add_so_sel_e                                add_state_out_sel;
  logic                                       add_state_out_sel_err;

  logic               [NumRegsData-1:0][31:0] data_out_d;
  logic               [NumRegsData-1:0][31:0] data_out_q;
  sp2v_e                                      data_out_we_ctrl;
  sp2v_e                                      data_out_we;
  logic               [NumRegsData-1:0]       data_out_re;
  logic               [NumRegsData-1:0]       data_out_re_buf;

  sp2v_e                                      cipher_in_valid;
  sp2v_e                                      cipher_in_ready;
  sp2v_e                                      cipher_out_valid;
  sp2v_e                                      cipher_out_ready;
  sp2v_e                                      cipher_crypt;
  sp2v_e                                      cipher_crypt_busy;
  sp2v_e                                      cipher_dec_key_gen;
  sp2v_e                                      cipher_dec_key_gen_busy;
  logic                                       cipher_prng_reseed;
  logic                                       cipher_prng_reseed_busy;
  logic                                       cipher_key_clear;
  logic                                       cipher_key_clear_busy;
  logic                                       cipher_data_out_clear;
  logic                                       cipher_data_out_clear_busy;
  logic                                       cipher_alert;

  // Pseudo-random data for clearing purposes
  logic                [WidthPRDClearing-1:0] cipher_prd_clearing [NumShares];
  logic                [WidthPRDClearing-1:0] prd_clearing [NumSharesKey];
  logic                                       prd_clearing_upd_req;
  logic                                       prd_clearing_upd_ack;
  logic                                       prd_clearing_rsd_req;
  logic                                       prd_clearing_rsd_ack;
  logic                               [127:0] prd_clearing_128 [NumShares];
  logic                               [255:0] prd_clearing_256 [NumSharesKey];

  // Unused signals
  logic               [NumRegsData-1:0][31:0] unused_data_out_q;

  // The clearing PRNG provides pseudo-random data for register clearing purposes.
  aes_prng_clearing #(
    .Width                ( WidthPRDClearing         ),
    .EntropyWidth         ( EntropyWidth             ),
    .SecSkipPRNGReseeding ( SecSkipPRNGReseeding     ),
    .RndCnstLfsrSeed      ( RndCnstClearingLfsrSeed  ),
    .RndCnstLfsrPerm      ( RndCnstClearingLfsrPerm  ),
    .RndCnstSharePerm     ( RndCnstClearingSharePerm )
  ) u_aes_prng_clearing (
    .clk_i         ( clk_i                  ),
    .rst_ni        ( rst_ni                 ),

    .data_req_i    ( prd_clearing_upd_req   ),
    .data_ack_o    ( prd_clearing_upd_ack   ),
    .data_o        ( prd_clearing           ),
    .reseed_req_i  ( prd_clearing_rsd_req   ),
    .reseed_ack_o  ( prd_clearing_rsd_ack   ),

    .entropy_req_o ( entropy_clearing_req_o ),
    .entropy_ack_i ( entropy_clearing_ack_i ),
    .entropy_i     ( entropy_clearing_i     )
  );

  // Generate clearing signals of appropriate widths.
  // Different shares need to be cleared with different pseudo-random data.
  for (genvar s = 0; s < NumShares; s++) begin : gen_prd_clearing_128_shares
    for (genvar c = 0; c < NumChunksPRDClearing128; c++) begin : gen_prd_clearing_128
      assign prd_clearing_128[s][c * WidthPRDClearing +: WidthPRDClearing] = prd_clearing[s];
    end
  end
  // The initial key is always provided in two shares. The two shares of the initial key register
  // need to be cleared with different pseudo-random data.
  for (genvar s = 0; s < NumSharesKey; s++) begin : gen_prd_clearing_256_shares
    for (genvar c = 0; c < NumChunksPRDClearing256; c++) begin : gen_prd_clearing_256
      assign prd_clearing_256[s][c * WidthPRDClearing +: WidthPRDClearing] = prd_clearing[s];
    end
  end

  ////////////
  // Inputs //
  ////////////

  always_comb begin : key_init_get
    for (int i = 0; i < NumRegsKey; i++) begin
      key_init[0][i]    = reg2hw.key_share0[i].q;
      key_init_qe[0][i] = reg2hw.key_share0[i].qe;
      key_init[1][i]    = reg2hw.key_share1[i].q;
      key_init_qe[1][i] = reg2hw.key_share1[i].qe;
    end
  end

  prim_sec_anchor_buf #(
    .Width ( NumSharesKey * NumRegsKey )
  ) u_prim_buf_key_init_qe (
    .in_i  ( {key_init_qe[1],     key_init_qe[0]}     ),
    .out_o ( {key_init_qe_buf[1], key_init_qe_buf[0]} )
  );

  always_comb begin : key_sideload_get
    for (int s = 0; s < NumSharesKey; s++) begin
      for (int i = 0; i < NumRegsKey; i++) begin
        key_sideload[s][i] = keymgr_key_i.key[s][i * 32 +: 32];
      end
    end
  end

  always_comb begin : iv_get
    for (int i = 0; i < NumRegsIv; i++) begin
      iv[i]    = reg2hw.iv[i].q;
      iv_qe[i] = reg2hw.iv[i].qe;
    end
  end

  prim_sec_anchor_buf #(
    .Width ( NumRegsIv )
  ) u_prim_buf_iv_qe (
    .in_i  ( iv_qe     ),
    .out_o ( iv_qe_buf )
  );

  always_comb begin : data_in_get
    for (int i = 0; i < NumRegsData; i++) begin
      data_in[i]    = reg2hw.data_in[i].q;
      data_in_qe[i] = reg2hw.data_in[i].qe;
    end
  end

  prim_sec_anchor_buf #(
    .Width ( NumRegsData )
  ) u_prim_buf_data_in_qe (
    .in_i  ( data_in_qe     ),
    .out_o ( data_in_qe_buf )
  );

  always_comb begin : data_out_get
    for (int i = 0; i < NumRegsData; i++) begin
      // data_out is actually hwo, but we need hrw for hwre
      unused_data_out_q[i] = reg2hw.data_out[i].q;
      data_out_re[i]       = reg2hw.data_out[i].re;
    end
  end

  prim_sec_anchor_buf #(
    .Width ( NumRegsData )
  ) u_prim_buf_data_out_re (
    .in_i  ( data_out_re     ),
    .out_o ( data_out_re_buf )
  );

  //////////////////////
  // Key, IV and Data //
  //////////////////////

  // SEC_CM: KEY.SEC_WIPE
  // SEC_CM: KEY.SIDELOAD
  // Initial Key registers
  always_comb begin : key_init_mux
    unique case (key_init_sel)
      KEY_INIT_INPUT:  key_init_d = key_init;
      KEY_INIT_KEYMGR: key_init_d = key_sideload;
      KEY_INIT_CLEAR:  key_init_d = prd_clearing_256;
      default:         key_init_d = prd_clearing_256;
    endcase
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : key_init_reg
    if (!rst_ni) begin
      key_init_q <= '{default: '0};
    end else begin
      for (int s = 0; s < NumSharesKey; s++) begin
        for (int i = 0; i < NumRegsKey; i++) begin
          if (key_init_we[s][i] == SP2V_HIGH) begin
            key_init_q[s][i] <= key_init_d[s][i];
          end
        end
      end
    end
  end

  // SEC_CM: IV.CONFIG.SEC_WIPE
  // IV registers
  always_comb begin : iv_mux
    unique case (iv_sel)
      IV_INPUT:        iv_d = iv;
      IV_DATA_OUT:     iv_d = data_out_d;
      IV_DATA_OUT_RAW: iv_d = aes_transpose(state_out);
      IV_DATA_IN_PREV: iv_d = data_in_prev_q;
      IV_CTR:          iv_d = ctr;
      IV_CLEAR:        iv_d = prd_clearing_128[0];
      default:         iv_d = prd_clearing_128[0];
    endcase
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : iv_reg
    if (!rst_ni) begin
      iv_q <= '0;
    end else begin
      for (int i = 0; i < NumSlicesCtr; i++) begin
        if (iv_we[i] == SP2V_HIGH) begin
          iv_q[i] <= iv_d[i];
        end
      end
    end
  end

  // SEC_CM: DATA_REG.SEC_WIPE
  // Previous input data register
  always_comb begin : data_in_prev_mux
    unique case (data_in_prev_sel)
      DIP_DATA_IN: data_in_prev_d = data_in;
      DIP_CLEAR:   data_in_prev_d = prd_clearing_128[0];
      default:     data_in_prev_d = prd_clearing_128[0];
    endcase
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : data_in_prev_reg
    if (!rst_ni) begin
      data_in_prev_q <= '0;
    end else if (data_in_prev_we == SP2V_HIGH) begin
      data_in_prev_q <= data_in_prev_d;
    end
  end

  /////////////
  // Counter //
  /////////////

  aes_ctr u_aes_ctr (
    .clk_i    ( clk_i     ),
    .rst_ni   ( rst_ni    ),

    .incr_i   ( ctr_incr  ),
    .ready_o  ( ctr_ready ),
    .alert_o  ( ctr_alert ),

    .ctr_i    ( iv_q      ),
    .ctr_o    ( ctr       ),
    .ctr_we_o ( ctr_we    )
  );

  /////////////////
  // Cipher Core //
  /////////////////

  // Cipher core operation
  assign cipher_op = (aes_mode_q == AES_ECB && aes_op_q == AES_ENC) ? CIPH_FWD :
                     (aes_mode_q == AES_ECB && aes_op_q == AES_DEC) ? CIPH_INV :
                     (aes_mode_q == AES_CBC && aes_op_q == AES_ENC) ? CIPH_FWD :
                     (aes_mode_q == AES_CBC && aes_op_q == AES_DEC) ? CIPH_INV :
                     (aes_mode_q == AES_CFB)                        ? CIPH_FWD :
                     (aes_mode_q == AES_OFB)                        ? CIPH_FWD :
                     (aes_mode_q == AES_CTR)                        ? CIPH_FWD : CIPH_FWD;

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  logic [$bits(ciph_op_e)-1:0] cipher_op_raw;
  prim_buf #(
    .Width($bits(ciph_op_e))
  ) u_prim_buf_op (
    .in_i(cipher_op),
    .out_o(cipher_op_raw)
  );
  assign cipher_op_buf = ciph_op_e'(cipher_op_raw);

  for (genvar s = 0; s < NumShares; s++) begin : gen_cipher_prd_clearing
    assign cipher_prd_clearing[s] = prd_clearing[s];
  end

  // Convert input data/IV to state format (every word corresponds to one state column).
  // Mux for state input
  always_comb begin : state_in_mux
    unique case (state_in_sel)
      SI_ZERO: state_in = '0;
      SI_DATA: state_in = aes_transpose(data_in);
      default: state_in = '0;
    endcase
  end

  // Mux for addition to state input
  always_comb begin : add_state_in_mux
    unique case (add_state_in_sel)
      ADD_SI_ZERO: add_state_in = '0;
      ADD_SI_IV:   add_state_in = aes_transpose(iv_q);
      default:     add_state_in = '0;
    endcase
  end

  if (!SecMasking) begin : gen_state_init_unmasked
    assign state_init[0] = state_in ^ add_state_in;

    logic [3:0][3:0][7:0] unused_state_mask;
    assign unused_state_mask = state_mask;

  end else begin : gen_state_init_masked
    assign state_init[0] = (state_in ^ add_state_in) ^ state_mask; // Masked data share
    assign state_init[1] = state_mask;                             // Mask share
  end

  if (!SecMasking) begin : gen_key_init_unmasked
    // Combine the two key shares for the unmasked cipher core. This causes SCA leakage of the key
    // and thus should be avoided.
    assign key_init_cipher[0] = key_init_q[0] ^ key_init_q[1];

  end else begin : gen_key_init_masked
    // Forward the masked key share and the mask share to the masked cipher core.
    assign key_init_cipher    = key_init_q;
  end

  // SEC_CM: KEY.MASKING
  // Cipher core
  aes_cipher_core #(
    .AES192Enable           ( AES192Enable           ),
    .SecMasking             ( SecMasking             ),
    .SecSBoxImpl            ( SecSBoxImpl            ),
    .SecAllowForcingMasks   ( SecAllowForcingMasks   ),
    .SecSkipPRNGReseeding   ( SecSkipPRNGReseeding   ),
    .RndCnstMaskingLfsrSeed ( RndCnstMaskingLfsrSeed ),
    .RndCnstMaskingLfsrPerm ( RndCnstMaskingLfsrPerm )
  ) u_aes_cipher_core (
    .clk_i            ( clk_i                      ),
    .rst_ni           ( rst_ni                     ),

    .in_valid_i       ( cipher_in_valid            ),
    .in_ready_o       ( cipher_in_ready            ),

    .out_valid_o      ( cipher_out_valid           ),
    .out_ready_i      ( cipher_out_ready           ),

    .cfg_valid_i      ( ~ctrl_err_storage          ), // Used for gating assertions only.
    .op_i             ( cipher_op_buf              ),
    .key_len_i        ( key_len_q                  ),
    .crypt_i          ( cipher_crypt               ),
    .crypt_o          ( cipher_crypt_busy          ),
    .dec_key_gen_i    ( cipher_dec_key_gen         ),
    .dec_key_gen_o    ( cipher_dec_key_gen_busy    ),
    .prng_reseed_i    ( cipher_prng_reseed         ),
    .prng_reseed_o    ( cipher_prng_reseed_busy    ),
    .key_clear_i      ( cipher_key_clear           ),
    .key_clear_o      ( cipher_key_clear_busy      ),
    .data_out_clear_i ( cipher_data_out_clear      ),
    .data_out_clear_o ( cipher_data_out_clear_busy ),
    .alert_fatal_i    ( alert_fatal_o              ),
    .alert_o          ( cipher_alert               ),

    .prd_clearing_i   ( cipher_prd_clearing        ),

    .force_masks_i    ( force_masks                ),
    .data_in_mask_o   ( state_mask                 ),
    .entropy_req_o    ( entropy_masking_req_o      ),
    .entropy_ack_i    ( entropy_masking_ack_i      ),
    .entropy_i        ( entropy_masking_i          ),

    .state_init_i     ( state_init                 ),
    .key_init_i       ( key_init_cipher            ),
    .state_o          ( state_done                 )
  );

  if (!SecMasking) begin : gen_state_out_unmasked
    assign state_out = state_done[0];
  end else begin : gen_state_out_masked
    // Unmask the cipher core output. This might get reworked in the future when masking the
    // counter and feedback path through the IV regs.

    // Only unmask the final cipher core output. Unmasking intermediate output data causes
    // additional SCA leakage and thus has to be avoided. Forward PRD instead of a determinsitic
    // value to avoid leaking the cipher core output when it becomes valid.
    logic [3:0][3:0][7:0] state_done_muxed [NumShares];
    for (genvar s = 0; s < NumShares; s++) begin : gen_state_done_muxed
      assign state_done_muxed[s] =
          (cipher_out_valid == SP2V_HIGH) ? state_done[s] : prd_clearing_128[s];
    end

    // Avoid aggressive synthesis optimizations.
    logic [3:0][3:0][7:0] state_done_buf [NumShares];
    prim_buf #(
      .Width ( 128 * NumShares )
    ) u_prim_state_done_muxed (
      .in_i  ( {state_done_muxed[1], state_done_muxed[0]} ),
      .out_o ( {state_done_buf[1],   state_done_buf[0]}   )
    );

    // Unmask the cipher core output.
    assign state_out = state_done_buf[0] ^ state_done_buf[1];
  end

  // Mux for addition to state output
  always_comb begin : add_state_out_mux
    unique case (add_state_out_sel)
      ADD_SO_ZERO: add_state_out = '0;
      ADD_SO_IV:   add_state_out = aes_transpose(iv_q);
      ADD_SO_DIP:  add_state_out = aes_transpose(data_in_prev_q);
      default:     add_state_out = '0;
    endcase
  end

  // Convert output state to output data format (every column corresponds to one output word).
  assign data_out_d = aes_transpose(state_out ^ add_state_out);

  //////////////////////
  // Control Register //
  //////////////////////

  // Shadowed register primitve
  aes_ctrl_reg_shadowed #(
    .AES192Enable ( AES192Enable )
  ) u_ctrl_reg_shadowed (
    .clk_i              ( clk_i                ),
    .rst_ni             ( rst_ni               ),
    .rst_shadowed_ni    ( rst_shadowed_ni      ),
    .qe_o               ( ctrl_qe              ),
    .we_i               ( ctrl_we              ),
    .phase_o            ( ctrl_phase           ),
    .operation_o        ( aes_op_q             ),
    .mode_o             ( aes_mode_q           ),
    .key_len_o          ( key_len_q            ),
    .sideload_o         ( sideload_q           ),
    .prng_reseed_rate_o ( prng_reseed_rate_q   ),
    .manual_operation_o ( manual_operation_q   ),
    .err_update_o       ( ctrl_reg_err_update  ),
    .err_storage_o      ( ctrl_reg_err_storage ),
    .reg2hw_ctrl_i      ( reg2hw.ctrl_shadowed ),
    .hw2reg_ctrl_o      ( hw2reg.ctrl_shadowed )
  );

  // Auxiliary control register signals
  assign key_touch_forces_reseed = reg2hw.ctrl_aux_shadowed.key_touch_forces_reseed.q;
  assign force_masks             = reg2hw.ctrl_aux_shadowed.force_masks.q;

  /////////////
  // Control //
  /////////////

  // Control
  aes_control #(
    .SecMasking           ( SecMasking           ),
    .SecStartTriggerDelay ( SecStartTriggerDelay )
  ) u_aes_control (
    .clk_i                     ( clk_i                                  ),
    .rst_ni                    ( rst_ni                                 ),

    .ctrl_qe_i                 ( ctrl_qe                                ),
    .ctrl_we_o                 ( ctrl_we                                ),
    .ctrl_phase_i              ( ctrl_phase                             ),
    .ctrl_err_storage_i        ( ctrl_err_storage                       ),
    .op_i                      ( aes_op_q                               ),
    .mode_i                    ( aes_mode_q                             ),
    .cipher_op_i               ( cipher_op_buf                          ),
    .sideload_i                ( sideload_q                             ),
    .prng_reseed_rate_i        ( prng_reseed_rate_q                     ),
    .manual_operation_i        ( manual_operation_q                     ),
    .key_touch_forces_reseed_i ( key_touch_forces_reseed                ),
    .start_i                   ( reg2hw.trigger.start.q                 ),
    .key_iv_data_in_clear_i    ( reg2hw.trigger.key_iv_data_in_clear.q  ),
    .data_out_clear_i          ( reg2hw.trigger.data_out_clear.q        ),
    .prng_reseed_i             ( reg2hw.trigger.prng_reseed.q           ),
    .mux_sel_err_i             ( mux_sel_err                            ),
    .sp_enc_err_i              ( sp_enc_err_q                           ),
    .lc_escalate_en_i          ( lc_escalate_en_i                       ),
    .alert_fatal_i             ( alert_fatal_o                          ),
    .alert_o                   ( ctrl_alert                             ),

    .key_sideload_valid_i      ( keymgr_key_i.valid                     ),
    .key_init_qe_i             ( key_init_qe_buf                        ),
    .iv_qe_i                   ( iv_qe_buf                              ),
    .data_in_qe_i              ( data_in_qe_buf                         ),
    .data_out_re_i             ( data_out_re_buf                        ),
    .data_in_we_o              ( data_in_we                             ),
    .data_out_we_o             ( data_out_we_ctrl                       ),

    .data_in_prev_sel_o        ( data_in_prev_sel_ctrl                  ),
    .data_in_prev_we_o         ( data_in_prev_we_ctrl                   ),

    .state_in_sel_o            ( state_in_sel_ctrl                      ),
    .add_state_in_sel_o        ( add_state_in_sel_ctrl                  ),
    .add_state_out_sel_o       ( add_state_out_sel_ctrl                 ),

    .ctr_incr_o                ( ctr_incr                               ),
    .ctr_ready_i               ( ctr_ready                              ),
    .ctr_we_i                  ( ctr_we                                 ),

    .cipher_in_valid_o         ( cipher_in_valid                        ),
    .cipher_in_ready_i         ( cipher_in_ready                        ),
    .cipher_out_valid_i        ( cipher_out_valid                       ),
    .cipher_out_ready_o        ( cipher_out_ready                       ),
    .cipher_crypt_o            ( cipher_crypt                           ),
    .cipher_crypt_i            ( cipher_crypt_busy                      ),
    .cipher_dec_key_gen_o      ( cipher_dec_key_gen                     ),
    .cipher_dec_key_gen_i      ( cipher_dec_key_gen_busy                ),
    .cipher_prng_reseed_o      ( cipher_prng_reseed                     ),
    .cipher_prng_reseed_i      ( cipher_prng_reseed_busy                ),
    .cipher_key_clear_o        ( cipher_key_clear                       ),
    .cipher_key_clear_i        ( cipher_key_clear_busy                  ),
    .cipher_data_out_clear_o   ( cipher_data_out_clear                  ),
    .cipher_data_out_clear_i   ( cipher_data_out_clear_busy             ),

    .key_init_sel_o            ( key_init_sel_ctrl                      ),
    .key_init_we_o             ( key_init_we_ctrl                       ),
    .iv_sel_o                  ( iv_sel_ctrl                            ),
    .iv_we_o                   ( iv_we_ctrl                             ),

    .prng_data_req_o           ( prd_clearing_upd_req                   ),
    .prng_data_ack_i           ( prd_clearing_upd_ack                   ),
    .prng_reseed_req_o         ( prd_clearing_rsd_req                   ),
    .prng_reseed_ack_i         ( prd_clearing_rsd_ack                   ),

    .start_o                   ( hw2reg.trigger.start.d                 ),
    .start_we_o                ( hw2reg.trigger.start.de                ),
    .key_iv_data_in_clear_o    ( hw2reg.trigger.key_iv_data_in_clear.d  ),
    .key_iv_data_in_clear_we_o ( hw2reg.trigger.key_iv_data_in_clear.de ),
    .data_out_clear_o          ( hw2reg.trigger.data_out_clear.d        ),
    .data_out_clear_we_o       ( hw2reg.trigger.data_out_clear.de       ),
    .prng_reseed_o             ( hw2reg.trigger.prng_reseed.d           ),
    .prng_reseed_we_o          ( hw2reg.trigger.prng_reseed.de          ),

    .idle_o                    ( hw2reg.status.idle.d                   ),
    .idle_we_o                 ( hw2reg.status.idle.de                  ),
    .stall_o                   ( hw2reg.status.stall.d                  ),
    .stall_we_o                ( hw2reg.status.stall.de                 ),
    .output_lost_i             ( reg2hw.status.output_lost.q            ),
    .output_lost_o             ( hw2reg.status.output_lost.d            ),
    .output_lost_we_o          ( hw2reg.status.output_lost.de           ),
    .output_valid_o            ( hw2reg.status.output_valid.d           ),
    .output_valid_we_o         ( hw2reg.status.output_valid.de          ),
    .input_ready_o             ( hw2reg.status.input_ready.d            ),
    .input_ready_we_o          ( hw2reg.status.input_ready.de           )
  );

  // SEC_CM: DATA_REG.SEC_WIPE
  // Input data register clear
  always_comb begin : data_in_reg_clear
    for (int i = 0; i < NumRegsData; i++) begin
      hw2reg.data_in[i].d  = prd_clearing_128[0][i * 32 +: 32];
      hw2reg.data_in[i].de = data_in_we;
    end
  end

  ///////////////
  // Selectors //
  ///////////////

  // We use sparse encodings for these mux selector signals and must ensure that:
  // 1. The synthesis tool doesn't optimize away the sparse encoding.
  // 2. The selector signal is always valid. More precisely, an alert or SVA is triggered if a
  //    selector signal takes on an invalid value.
  // 3. The alert signal remains asserted until reset even if the selector signal becomes valid
  //    again. This is achieved by driving the control FSM into the terminal error state whenever
  //    any mux selector signal becomes invalid.
  //
  // If any mux selector signal becomes invalid, the control FSM further prevents any data from
  // being released from the cipher core by de-asserting the write enable of the output data
  // registers.

  aes_sel_buf_chk #(
    .Num      ( DIPSelNum   ),
    .Width    ( DIPSelWidth ),
    .EnSecBuf ( 1'b1        )
  ) u_aes_data_in_prev_sel_buf_chk (
    .clk_i  ( clk_i                 ),
    .rst_ni ( rst_ni                ),
    .sel_i  ( data_in_prev_sel_ctrl ),
    .sel_o  ( data_in_prev_sel_raw  ),
    .err_o  ( data_in_prev_sel_err  )
  );
  assign data_in_prev_sel = dip_sel_e'(data_in_prev_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( SISelNum   ),
    .Width    ( SISelWidth ),
    .EnSecBuf ( 1'b1       )
  ) u_aes_state_in_sel_buf_chk (
    .clk_i  ( clk_i             ),
    .rst_ni ( rst_ni            ),
    .sel_i  ( state_in_sel_ctrl ),
    .sel_o  ( state_in_sel_raw  ),
    .err_o  ( state_in_sel_err  )
  );
  assign state_in_sel = si_sel_e'(state_in_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( AddSISelNum   ),
    .Width    ( AddSISelWidth ),
    .EnSecBuf ( 1'b1          )
  ) u_aes_add_state_in_sel_buf_chk (
    .clk_i  ( clk_i                 ),
    .rst_ni ( rst_ni                ),
    .sel_i  ( add_state_in_sel_ctrl ),
    .sel_o  ( add_state_in_sel_raw  ),
    .err_o  ( add_state_in_sel_err  )
  );
  assign add_state_in_sel = add_si_sel_e'(add_state_in_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( AddSOSelNum   ),
    .Width    ( AddSOSelWidth ),
    .EnSecBuf ( 1'b1          )
  ) u_aes_add_state_out_sel_buf_chk (
    .clk_i  ( clk_i                  ),
    .rst_ni ( rst_ni                 ),
    .sel_i  ( add_state_out_sel_ctrl ),
    .sel_o  ( add_state_out_sel_raw  ),
    .err_o  ( add_state_out_sel_err  )
  );
  assign add_state_out_sel = add_so_sel_e'(add_state_out_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( KeyInitSelNum   ),
    .Width    ( KeyInitSelWidth ),
    .EnSecBuf ( 1'b1            )
  ) u_aes_key_init_sel_buf_chk (
    .clk_i  ( clk_i             ),
    .rst_ni ( rst_ni            ),
    .sel_i  ( key_init_sel_ctrl ),
    .sel_o  ( key_init_sel_raw  ),
    .err_o  ( key_init_sel_err  )
  );
  assign key_init_sel = key_init_sel_e'(key_init_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( IVSelNum   ),
    .Width    ( IVSelWidth ),
    .EnSecBuf ( 1'b1       )
  ) u_aes_iv_sel_buf_chk (
    .clk_i  ( clk_i       ),
    .rst_ni ( rst_ni      ),
    .sel_i  ( iv_sel_ctrl ),
    .sel_o  ( iv_sel_raw  ),
    .err_o  ( iv_sel_err  )
  );
  assign iv_sel = iv_sel_e'(iv_sel_raw);

  // Signal invalid mux selector signals to control FSM which will lock up and trigger an alert.
  assign mux_sel_err = data_in_prev_sel_err | state_in_sel_err | add_state_in_sel_err |
      add_state_out_sel_err | key_init_sel_err | iv_sel_err;

  //////////////////////////////
  // Sparsely Encoded Signals //
  //////////////////////////////

  // We use sparse encodings for various critical signals and must ensure that:
  // 1. The synthesis tool doesn't optimize away the sparse encoding.
  // 2. The sparsely encoded signal is always valid. More precisely, an alert or SVA is triggered
  //    if a sparse signal takes on an invalid value.
  // 3. The alert signal remains asserted until reset even if the sparse signal becomes valid again
  //    This is achieved by driving the control FSM into the terminal error state whenever any
  //    sparsely encoded signal becomes invalid.
  //
  // If any sparsely encoded signal becomes invalid, the core controller further immediately
  // de-asserts the data_out_we_o signal to prevent any data from being released.

  // We use vectors of sparsely encoded signals to reduce code duplication.
  localparam int unsigned NumSp2VSig = NumSharesKey * NumRegsKey + NumSlicesCtr + 2;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig_chk;
  logic  [NumSp2VSig-1:0][Sp2VWidth-1:0] sp2v_sig_chk_raw;
  logic  [NumSp2VSig-1:0]                sp2v_sig_err;

  for (genvar s = 0; s < NumSharesKey; s++) begin : gen_use_key_init_we_ctrl_shares
    for (genvar i = 0; i < NumRegsKey; i++) begin : gen_use_key_init_we_ctrl
      assign sp2v_sig[s * NumRegsKey + i] = key_init_we_ctrl[s][i];
    end
  end
  for (genvar i = 0; i < NumSlicesCtr; i++) begin : gen_use_iv_we_ctrl
    assign sp2v_sig[NumSharesKey * NumRegsKey + i] = iv_we_ctrl[i];
  end
  assign sp2v_sig[NumSharesKey * NumRegsKey + NumSlicesCtr + 0] = data_in_prev_we_ctrl;
  assign sp2v_sig[NumSharesKey * NumRegsKey + NumSlicesCtr + 1] = data_out_we_ctrl;

  // All signals inside sp2v_sig are eventually converted to single-rail signals.
  localparam bit [NumSp2VSig-1:0] Sp2VEnSecBuf = {NumSp2VSig{1'b1}};

  // Individually check sparsely encoded signals.
  for (genvar i = 0; i < NumSp2VSig; i++) begin : gen_sel_buf_chk
    aes_sel_buf_chk #(
      .Num      ( Sp2VNum         ),
      .Width    ( Sp2VWidth       ),
      .EnSecBuf ( Sp2VEnSecBuf[i] )
    ) u_aes_sp2v_sig_buf_chk_i (
      .clk_i  ( clk_i               ),
      .rst_ni ( rst_ni              ),
      .sel_i  ( sp2v_sig[i]         ),
      .sel_o  ( sp2v_sig_chk_raw[i] ),
      .err_o  ( sp2v_sig_err[i]     )
    );
    assign sp2v_sig_chk[i] = sp2v_e'(sp2v_sig_chk_raw[i]);
  end

  for (genvar s = 0; s < NumSharesKey; s++) begin : gen_key_init_we_shares
    for (genvar i = 0; i < NumRegsKey; i++) begin : gen_key_init_we
      assign key_init_we[s][i] = sp2v_sig_chk[s * NumRegsKey + i];
    end
  end
  for (genvar i = 0; i < NumSlicesCtr; i++) begin : gen_iv_we
    assign iv_we[i]      = sp2v_sig_chk[NumSharesKey * NumRegsKey + i];
  end
  assign data_in_prev_we = sp2v_sig_chk[NumSharesKey * NumRegsKey + NumSlicesCtr + 0];
  assign data_out_we     = sp2v_sig_chk[NumSharesKey * NumRegsKey + NumSlicesCtr + 1];

  // Collect encoding errors.
  // We instantiate the checker modules as close as possible to where the sparsely encoded signals
  // are used. Here, we collect also encoding errors detected in other places of the core.
  assign sp_enc_err_d = |sp2v_sig_err;

  // We need to register the collected error signal to avoid circular loops in the core controller
  // related to iv_we and data_out_we.
  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_sp_enc_err
    if (!rst_ni) begin
      sp_enc_err_q <= 1'b0;
    end else if (sp_enc_err_d) begin
      sp_enc_err_q <= 1'b1;
    end
  end

  /////////////
  // Outputs //
  /////////////

  always_ff @(posedge clk_i or negedge rst_ni) begin : data_out_reg
    if (!rst_ni) begin
      data_out_q <= '0;
    end else if (data_out_we == SP2V_HIGH) begin
      data_out_q <= data_out_d;
    end
  end

  always_comb begin : key_reg_put
    for (int i = 0; i < NumRegsKey; i++) begin
      hw2reg.key_share0[i].d = key_init_q[0][i];
      hw2reg.key_share1[i].d = key_init_q[1][i];
    end
  end

  always_comb begin : iv_reg_put
    for (int i = 0; i < NumRegsIv; i++) begin
      // Software updates IV in chunks of 32 bits. Internally, the counter updates SliceSizeCtr
      // bits at a time.
      hw2reg.iv[i].d  = {iv_q[2 * i + 1], iv_q[2 * i]};
    end
  end

  always_comb begin : data_out_put
    for (int i = 0; i < NumRegsData; i++) begin
      hw2reg.data_out[i].d = data_out_q[i];
    end
  end

  ////////////
  // Alerts //
  ////////////

  // Should fatal alerts clear the status register?
  assign clear_on_fatal = ClearStatusOnFatalAlert ? alert_fatal_o : 1'b0;

  // Recoverable alert conditions are signaled as a single alert event.
  assign ctrl_err_update = ctrl_reg_err_update | shadowed_update_err_i;
  assign alert_recov_o = ctrl_err_update;

  // The recoverable alert is observable via status register until the AES operation is restarted
  // by re-writing the Control Register. Fatal alerts clear all other bits in the status register.
  assign hw2reg.status.alert_recov_ctrl_update_err.d  = ctrl_err_update & ~clear_on_fatal;
  assign hw2reg.status.alert_recov_ctrl_update_err.de = ctrl_err_update | ctrl_we | clear_on_fatal;

  // Fatal alert conditions need to remain asserted until reset.
  assign ctrl_err_storage_d = ctrl_reg_err_storage | shadowed_storage_err_i;
  always_ff @(posedge clk_i or negedge rst_ni) begin : ctrl_err_storage_reg
    if (!rst_ni) begin
      ctrl_err_storage_q <= 1'b0;
    end else if (ctrl_err_storage_d) begin
      ctrl_err_storage_q <= 1'b1;
    end
  end
  assign ctrl_err_storage = ctrl_err_storage_d | ctrl_err_storage_q;

  // Collect fatal alert signals.
  assign alert_fatal_o = ctrl_err_storage |
                         ctr_alert        |
                         cipher_alert     |
                         ctrl_alert       |
                         intg_err_alert_i;

  // Make the fatal alert observable via status register.
  assign hw2reg.status.alert_fatal_fault.d  = alert_fatal_o;
  assign hw2reg.status.alert_fatal_fault.de = alert_fatal_o;

  // Unused alert signals
  logic unused_alert_signals;
  assign unused_alert_signals = ^reg2hw.alert_test;

  // Unused inputs
  logic unused_idle;
  assign unused_idle = reg2hw.status.idle.q;

  ////////////////
  // Assertions //
  ////////////////

  // Create a lint error to reduce the risk of accidentally disabling the masking.
  `ASSERT_STATIC_LINT_ERROR(AesCoreSecMaskingNonDefault, SecMasking == 1)

  // Selectors must be known/valid
  `ASSERT(AesModeValid, !ctrl_err_storage |-> aes_mode_q inside {
      AES_ECB,
      AES_CBC,
      AES_CFB,
      AES_OFB,
      AES_CTR,
      AES_NONE
      })
  `ASSERT(AesOpValid, !ctrl_err_storage |-> aes_op_q inside {
      AES_ENC,
      AES_DEC
      })

  // Check parameters
  `ASSERT_INIT(AesNumSlicesCtr, NumSlicesCtr == 8)

  // Signals used for assertions only.
  logic [3:0][31:0] state_done_transposed, unused_state_done_transposed;
  if (!SecMasking) begin : gen_state_done_transposed_unmasked
    assign state_done_transposed = aes_transpose(state_done[0]);
  end else begin : gen_state_done_transposed_masked
    assign state_done_transposed = aes_transpose(state_done[0] ^ state_done[1]);
  end
  assign unused_state_done_transposed = state_done_transposed;

  // Ensure that upon local escalation of any of the FSMs, no intermediate state is released from
  // the cipher core into the software readable output data or IV registers.
  `ASSERT(AesSecCmDataRegLocalEscDataOut, $changed(data_out_q) && alert_fatal_o &&
      ($past(cipher_crypt, 2) == SP2V_HIGH || $past(cipher_crypt_busy, 2) == SP2V_HIGH) |=>
      ($past(data_out_q) != $past(state_done_transposed, 2)) &&
      ($past(data_out_q) != $past(state_done_transposed, 2) ^ $past(iv_q, 2)) &&
      ($past(data_out_q) != $past(state_done_transposed, 2) ^ $past(data_in_prev_q, 2)))

  `ASSERT(AesSecCmDataRegLocalEscIv, $changed(iv_q) && alert_fatal_o &&
      ($past(cipher_crypt, 2) == SP2V_HIGH || $past(cipher_crypt_busy, 2) == SP2V_HIGH) |=>
      ($past(iv_q) != $past(state_done_transposed, 2)) &&
      ($past(iv_q) != $past(state_done_transposed, 2) ^ $past(iv_q, 2)) &&
      ($past(iv_q) != $past(state_done_transposed, 2) ^ $past(data_in_prev_q, 2)))

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES counter for CTR mode
//
// This module uses one counter with a width of SliceSizeCtr to iteratively increment the 128-bit
// counter value.

module aes_ctr import aes_pkg::*;
(
  input  logic                                       clk_i,
  input  logic                                       rst_ni,

  input  sp2v_e                                      incr_i,
  output sp2v_e                                      ready_o,
  output logic                                       alert_o,

  input  logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] ctr_i,
  output logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] ctr_o,
  output sp2v_e [NumSlicesCtr-1:0]                   ctr_we_o
);

  // Reverse byte order - unrelated to NumSlicesCtr and SliceSizeCtr
  function automatic logic [15:0][7:0] aes_rev_order_byte(logic [15:0][7:0] in);
    logic [15:0][7:0] out;
    for (int i = 0; i < 16; i++) begin
      out[i] = in[15-i];
    end
    return out;
  endfunction

  // Reverse sp2v order
  function automatic sp2v_e [NumSlicesCtr-1:0] aes_rev_order_sp2v(sp2v_e [NumSlicesCtr-1:0] in);
    sp2v_e [NumSlicesCtr-1:0] out;
    for (int i = 0; i < NumSlicesCtr; i++) begin
      out[i] = in[NumSlicesCtr - 1 - i];
    end
    return out;
  endfunction

  // Signals
  logic                   [SliceIdxWidth-1:0] ctr_slice_idx;

  logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] ctr_i_rev; // 8 times 2 bytes
  logic  [NumSlicesCtr-1:0][SliceSizeCtr-1:0] ctr_o_rev; // 8 times 2 bytes
  sp2v_e [NumSlicesCtr-1:0]                   ctr_we_o_rev;
  sp2v_e                                      ctr_we;

  logic                    [SliceSizeCtr-1:0] ctr_i_slice;
  logic                    [SliceSizeCtr-1:0] ctr_o_slice;

  sp2v_e                                      incr;
  logic                                       incr_err;
  logic                                       mr_err;

  // Sparsified FSM signals. These are needed for connecting the individual bits of the Sp2V
  // signals to the single-rail FSMs.
  logic    [Sp2VWidth-1:0]                    sp_incr;
  logic    [Sp2VWidth-1:0]                    sp_ready;
  logic    [Sp2VWidth-1:0]                    sp_ctr_we;

  // Multi-rail signals. These are outputs of the single-rail FSMs and need combining.
  logic    [Sp2VWidth-1:0]                    mr_alert;
  logic    [Sp2VWidth-1:0][SliceIdxWidth-1:0] mr_ctr_slice_idx;
  logic    [Sp2VWidth-1:0] [SliceSizeCtr-1:0] mr_ctr_o_slice;

  ////////////
  // Inputs //
  ////////////

  // Reverse byte order
  assign ctr_i_rev = aes_rev_order_byte(ctr_i);

  // SEC_CM: CTRL.SPARSE
  // Check sparsely encoded incr signal.
  logic [Sp2VWidth-1:0] incr_raw;
  aes_sel_buf_chk #(
    .Num      ( Sp2VNum   ),
    .Width    ( Sp2VWidth ),
    .EnSecBuf ( 1'b0      )
  ) u_aes_sb_en_buf_chk (
    .clk_i  ( clk_i    ),
    .rst_ni ( rst_ni   ),
    .sel_i  ( incr_i   ),
    .sel_o  ( incr_raw ),
    .err_o  ( incr_err )
  );
  assign incr = sp2v_e'(incr_raw);

  /////////////
  // Counter //
  /////////////

  // We do SliceSizeCtr bits at a time.
  assign ctr_i_slice = ctr_i_rev[ctr_slice_idx];

  /////////
  // FSM //
  /////////

  // Convert sp2v_e signals to sparsified inputs.
  assign sp_incr = {incr};

  // SEC_CM: CTR.FSM.REDUN
  // For every bit in the Sp2V signals, one separate rail is instantiated. The inputs and outputs
  // of every rail are buffered to prevent aggressive synthesis optimizations.
  for (genvar i = 0; i < Sp2VWidth; i++) begin : gen_fsm
    if (SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_fsm_p
      aes_ctr_fsm_p u_aes_ctr_fsm_i (
        .clk_i           ( clk_i               ),
        .rst_ni          ( rst_ni              ),

        .incr_i          ( sp_incr[i]          ), // Sparsified
        .ready_o         ( sp_ready[i]         ), // Sparsified
        .incr_err_i      ( incr_err            ),
        .mr_err_i        ( mr_err              ),
        .alert_o         ( mr_alert[i]         ), // OR-combine

        .ctr_slice_idx_o ( mr_ctr_slice_idx[i] ), // OR-combine
        .ctr_slice_i     ( ctr_i_slice         ),
        .ctr_slice_o     ( mr_ctr_o_slice[i]   ), // OR-combine
        .ctr_we_o        ( sp_ctr_we[i]        )  // Sparsified
      );
    end else begin : gen_fsm_n
      aes_ctr_fsm_n u_aes_ctr_fsm_i (
        .clk_i           ( clk_i               ),
        .rst_ni          ( rst_ni              ),

        .incr_ni         ( sp_incr[i]          ), // Sparsified
        .ready_no        ( sp_ready[i]         ), // Sparsified
        .incr_err_i      ( incr_err            ),
        .mr_err_i        ( mr_err              ),
        .alert_o         ( mr_alert[i]         ), // OR-combine

        .ctr_slice_idx_o ( mr_ctr_slice_idx[i] ), // OR-combine
        .ctr_slice_i     ( ctr_i_slice         ),
        .ctr_slice_o     ( mr_ctr_o_slice[i]   ), // OR-combine
        .ctr_we_no       ( sp_ctr_we[i]        )  // Sparsified
      );
    end
  end

  // Convert sparsified outputs to sp2v_e type.
  assign ready_o = sp2v_e'(sp_ready);
  assign ctr_we  = sp2v_e'(sp_ctr_we);

  // Combine single-bit FSM outputs.
  // OR: One bit is sufficient to drive the corresponding output bit high.
  assign alert_o = |mr_alert;

  // Combine multi-bit FSM outputs. We simply OR them together and compare the values
  // to detect errors.
  always_comb begin : combine_sparse_signals
    ctr_slice_idx = '0;
    ctr_o_slice   = '0;
    mr_err        = 1'b0;

    for (int i = 0; i < Sp2VWidth; i++) begin
      ctr_slice_idx |= mr_ctr_slice_idx[i];
      ctr_o_slice   |= mr_ctr_o_slice[i];
    end

    for (int i = 0; i < Sp2VWidth; i++) begin
      if (ctr_slice_idx != mr_ctr_slice_idx[i] ||
          ctr_o_slice   != mr_ctr_o_slice[i]) begin
        mr_err = 1'b1;
      end
    end
  end

  /////////////
  // Outputs //
  /////////////

  // Combine input and counter output.
  always_comb begin
    ctr_o_rev                = ctr_i_rev;
    ctr_o_rev[ctr_slice_idx] = ctr_o_slice;
  end

  // Generate the sliced write enable.
  always_comb begin
    ctr_we_o_rev                = {NumSlicesCtr{SP2V_LOW}};
    ctr_we_o_rev[ctr_slice_idx] = ctr_we;
  end

  // Reverse byte and bit order.
  assign ctr_o    = aes_rev_order_byte(ctr_o_rev);
  assign ctr_we_o = aes_rev_order_sp2v(ctr_we_o_rev);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES counter FSM for CTR mode

`include "prim_assert.sv"

module aes_ctr_fsm import aes_pkg::*;
(
  input  logic                     clk_i,
  input  logic                     rst_ni,

  input  logic                     incr_i,     // Sparsify using multi-rail.
  output logic                     ready_o,    // Sparsify using multi-rail.
  input  logic                     incr_err_i,
  input  logic                     mr_err_i,
  output logic                     alert_o,

  output logic [SliceIdxWidth-1:0] ctr_slice_idx_o,
  input  logic  [SliceSizeCtr-1:0] ctr_slice_i,
  output logic  [SliceSizeCtr-1:0] ctr_slice_o,
  output logic                     ctr_we_o    // Sparsify using multi-rail.
);

  // Signals
  aes_ctr_e                 aes_ctr_ns, aes_ctr_cs;
  logic [SliceIdxWidth-1:0] ctr_slice_idx_d, ctr_slice_idx_q;
  logic                     ctr_carry_d, ctr_carry_q;

  logic    [SliceSizeCtr:0] ctr_value;

  /////////////
  // Counter //
  /////////////

  // We do SliceSizeCtr bits at a time.
  assign ctr_value   = ctr_slice_i + {{(SliceSizeCtr-1){1'b0}}, ctr_carry_q};
  assign ctr_slice_o = ctr_value[SliceSizeCtr-1:0];

  /////////////
  // Control //
  /////////////

  // FSM
  always_comb begin : aes_ctr_fsm_comb

    // Outputs
    ready_o         = 1'b0;
    ctr_we_o        = 1'b0;
    alert_o         = 1'b0;

    // FSM
    aes_ctr_ns      = aes_ctr_cs;
    ctr_slice_idx_d = ctr_slice_idx_q;
    ctr_carry_d     = ctr_carry_q;

    unique case (aes_ctr_cs)
      CTR_IDLE: begin
        ready_o = 1'b1;
        if (incr_i == 1'b1) begin
          // Initialize slice index and carry bit.
          ctr_slice_idx_d = '0;
          ctr_carry_d     = 1'b1;
          aes_ctr_ns      = CTR_INCR;
        end
      end

      CTR_INCR: begin
        // Increment slice index.
        ctr_slice_idx_d = ctr_slice_idx_q + SliceIdxWidth'(1);
        ctr_carry_d     = ctr_value[SliceSizeCtr];
        ctr_we_o        = 1'b1;

        if (ctr_slice_idx_q == {SliceIdxWidth{1'b1}}) begin
          aes_ctr_ns = CTR_IDLE;
        end
      end

      CTR_ERROR: begin
        // SEC_CM: CTR.FSM.LOCAL_ESC
        // Terminal error state
        alert_o = 1'b1;
      end

      // We should never get here. If we do (e.g. via a malicious
      // glitch), error out immediately.
      default: begin
        aes_ctr_ns = CTR_ERROR;
        alert_o = 1'b1;
      end
    endcase

    // Unconditionally jump into the terminal error state in case an error is detected.
    if (incr_err_i || mr_err_i) begin
      aes_ctr_ns = CTR_ERROR;
    end
  end

  // Registers
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      ctr_slice_idx_q <= '0;
      ctr_carry_q     <= '0;
    end else begin
      ctr_slice_idx_q <= ctr_slice_idx_d;
      ctr_carry_q     <= ctr_carry_d;
    end
  end

  // SEC_CM: CTR.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, aes_ctr_ns, aes_ctr_cs, aes_ctr_e, CTR_IDLE)

  // Forward slice index.
  assign ctr_slice_idx_o = ctr_slice_idx_q;

  ////////////////
  // Assertions //
  ////////////////
  `ASSERT(AesCtrStateValid, !alert_o |-> aes_ctr_cs inside {
      CTR_IDLE,
      CTR_INCR
      })

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES counter FSM for CTR mode
//
// This module contains the AES counter FSM operating on and producing the positive values of
// important control signals.

module aes_ctr_fsm_p import aes_pkg::*;
(
  input  logic                     clk_i,
  input  logic                     rst_ni,

  input  logic                     incr_i,          // Sparsify
  output logic                     ready_o,         // Sparsify
  input  logic                     incr_err_i,
  input  logic                     mr_err_i,
  output logic                     alert_o,

  output logic [SliceIdxWidth-1:0] ctr_slice_idx_o,
  input  logic  [SliceSizeCtr-1:0] ctr_slice_i,
  output logic  [SliceSizeCtr-1:0] ctr_slice_o,
  output logic                     ctr_we_o         // Sparsify
);

  /////////////////////
  // Input Buffering //
  /////////////////////

  localparam int NumInBufBits = $bits({
    incr_i,
    incr_err_i,
    mr_err_i,
    ctr_slice_i
  });

  logic [NumInBufBits-1:0] in, in_buf;

  assign in = {
    incr_i,
    incr_err_i,
    mr_err_i,
    ctr_slice_i
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumInBufBits)
  ) u_prim_buf_in (
    .in_i(in),
    .out_o(in_buf)
  );

  logic                    incr;
  logic                    incr_err;
  logic                    mr_err;
  logic [SliceSizeCtr-1:0] ctr_i_slice;

  assign {incr,
          incr_err,
          mr_err,
          ctr_i_slice} = in_buf;

  // Intermediate output signals
  logic                     ready;
  logic                     alert;
  logic [SliceIdxWidth-1:0] ctr_slice_idx;
  logic  [SliceSizeCtr-1:0] ctr_o_slice;
  logic                     ctr_we;

  /////////////////
  // Regular FSM //
  /////////////////

  aes_ctr_fsm u_aes_ctr_fsm (
    .clk_i           ( clk_i         ),
    .rst_ni          ( rst_ni        ),

    .incr_i          ( incr          ),
    .ready_o         ( ready         ),
    .incr_err_i      ( incr_err      ),
    .mr_err_i        ( mr_err        ),
    .alert_o         ( alert         ),

    .ctr_slice_idx_o ( ctr_slice_idx ),
    .ctr_slice_i     ( ctr_i_slice   ),
    .ctr_slice_o     ( ctr_o_slice   ),
    .ctr_we_o        ( ctr_we        )
  );

  //////////////////////
  // Output Buffering //
  //////////////////////

  localparam int NumOutBufBits = $bits({
    ready_o,
    alert_o,
    ctr_slice_idx_o,
    ctr_slice_o,
    ctr_we_o
  });

  logic [NumOutBufBits-1:0] out, out_buf;

  assign out = {
    ready,
    alert,
    ctr_slice_idx,
    ctr_o_slice,
    ctr_we
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumOutBufBits)
  ) u_prim_buf_out (
    .in_i(out),
    .out_o(out_buf)
  );

  assign {ready_o,
          alert_o,
          ctr_slice_idx_o,
          ctr_slice_o,
          ctr_we_o} = out_buf;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES counter FSM for CTR mode
//
// This module contains the AES counter FSM operating on and producing the negated values of
// important control signals. This is achieved by:
// - instantiating the regular AES counter FSM operating on and producing the positive values of
//   these signals, and
// - inverting these signals between the regular FSM and the prim_buf synthesis barriers.
// Synthesis tools will then push the inverters into the actual FSM.

module aes_ctr_fsm_n import aes_pkg::*;
(
  input  logic                     clk_i,
  input  logic                     rst_ni,

  input  logic                     incr_ni,         // Sparsify using multi-rail.
  output logic                     ready_no,        // Sparsify using multi-rail.
  input  logic                     incr_err_i,
  input  logic                     mr_err_i,
  output logic                     alert_o,

  output logic [SliceIdxWidth-1:0] ctr_slice_idx_o,
  input  logic  [SliceSizeCtr-1:0] ctr_slice_i,
  output logic  [SliceSizeCtr-1:0] ctr_slice_o,
  output logic                     ctr_we_no        // Sparsify using multi-rail.
);

  /////////////////////
  // Input Buffering //
  /////////////////////

  localparam int NumInBufBits = $bits({
    incr_ni,
    incr_err_i,
    mr_err_i,
    ctr_slice_i
  });

  logic [NumInBufBits-1:0] in, in_buf;

  assign in = {
    incr_ni,
    incr_err_i,
    mr_err_i,
    ctr_slice_i
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumInBufBits)
  ) u_prim_buf_in (
    .in_i(in),
    .out_o(in_buf)
  );

  logic                    incr_n;
  logic                    incr_err;
  logic                    mr_err;
  logic [SliceSizeCtr-1:0] ctr_i_slice;

  assign {incr_n,
          incr_err,
          mr_err,
          ctr_i_slice} = in_buf;

  // Intermediate output signals
  logic                     ready;
  logic                     alert;
  logic [SliceIdxWidth-1:0] ctr_slice_idx;
  logic  [SliceSizeCtr-1:0] ctr_o_slice;
  logic                     ctr_we;

  /////////////////
  // Regular FSM //
  /////////////////

  // The regular FSM operates on and produces the positive values of important control signals.
  // Invert *_n input signals here to get the positive values for the regular FSM. To obtain the
  // negated outputs, important output signals are inverted further below. Thanks to the prim_buf
  // synthesis optimization barriers, tools will push the inverters into the regular FSM.
  aes_ctr_fsm u_aes_ctr_fsm (
    .clk_i           ( clk_i         ),
    .rst_ni          ( rst_ni        ),

    .incr_i          ( ~incr_n       ), // Invert for regular FSM.
    .ready_o         ( ready         ), // Invert below for negated output.
    .incr_err_i      ( incr_err      ),
    .mr_err_i        ( mr_err        ),
    .alert_o         ( alert         ),

    .ctr_slice_idx_o ( ctr_slice_idx ),
    .ctr_slice_i     ( ctr_i_slice   ),
    .ctr_slice_o     ( ctr_o_slice   ),
    .ctr_we_o        ( ctr_we        )  // Invert below for negated output.
  );

  //////////////////////
  // Output Buffering //
  //////////////////////

  localparam int NumOutBufBits = $bits({
    ready_no,
    alert_o,
    ctr_slice_idx_o,
    ctr_slice_o,
    ctr_we_no
  });

  logic [NumOutBufBits-1:0] out, out_buf;

  // Important output control signals need to be inverted here. Synthesis tools will push the
  // inverters back into the regular FSM.
  assign out = {
    ~ready,
    alert,
    ctr_slice_idx,
    ctr_o_slice,
    ~ctr_we
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumOutBufBits)
  ) u_prim_buf_out (
    .in_i(out),
    .out_o(out_buf)
  );

  assign {ready_no,
          alert_o,
          ctr_slice_idx_o,
          ctr_slice_o,
          ctr_we_no} = out_buf;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES main control
//
// This module controls the interplay of input/output registers and the AES cipher core.

`include "prim_assert.sv"

module aes_control
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          SecMasking           = 0,
  parameter int unsigned SecStartTriggerDelay = 0
) (
  input  logic                      clk_i,
  input  logic                      rst_ni,

  // Main control signals
  input  logic                      ctrl_qe_i,
  output logic                      ctrl_we_o,
  input  logic                      ctrl_phase_i,
  input  logic                      ctrl_err_storage_i,
  input  aes_op_e                   op_i,
  input  aes_mode_e                 mode_i,
  input  ciph_op_e                  cipher_op_i,
  input  logic                      sideload_i,
  input  prs_rate_e                 prng_reseed_rate_i,
  input  logic                      manual_operation_i,
  input  logic                      key_touch_forces_reseed_i,
  input  logic                      start_i,
  input  logic                      key_iv_data_in_clear_i,
  input  logic                      data_out_clear_i,
  input  logic                      prng_reseed_i,
  input  logic                      mux_sel_err_i,
  input  logic                      sp_enc_err_i,
  input  lc_ctrl_pkg::lc_tx_t       lc_escalate_en_i,
  input  logic                      alert_fatal_i,
  output logic                      alert_o,

  // I/O register read/write enables
  input  logic                      key_sideload_valid_i,
  input  logic     [NumRegsKey-1:0] key_init_qe_i [NumSharesKey],
  input  logic      [NumRegsIv-1:0] iv_qe_i,
  input  logic    [NumRegsData-1:0] data_in_qe_i,
  input  logic    [NumRegsData-1:0] data_out_re_i,
  output logic                      data_in_we_o,
  output sp2v_e                     data_out_we_o,

  // Previous input data register
  output dip_sel_e                  data_in_prev_sel_o,
  output sp2v_e                     data_in_prev_we_o,

  // Cipher I/O muxes
  output si_sel_e                   state_in_sel_o,
  output add_si_sel_e               add_state_in_sel_o,
  output add_so_sel_e               add_state_out_sel_o,

  // Counter
  output sp2v_e                     ctr_incr_o,
  input  sp2v_e                     ctr_ready_i,
  input  sp2v_e  [NumSlicesCtr-1:0] ctr_we_i,

  // Cipher core control and sync
  output sp2v_e                     cipher_in_valid_o,
  input  sp2v_e                     cipher_in_ready_i,
  input  sp2v_e                     cipher_out_valid_i,
  output sp2v_e                     cipher_out_ready_o,
  output sp2v_e                     cipher_crypt_o,
  input  sp2v_e                     cipher_crypt_i,
  output sp2v_e                     cipher_dec_key_gen_o,
  input  sp2v_e                     cipher_dec_key_gen_i,
  output logic                      cipher_prng_reseed_o,
  input  logic                      cipher_prng_reseed_i,
  output logic                      cipher_key_clear_o,
  input  logic                      cipher_key_clear_i,
  output logic                      cipher_data_out_clear_o,
  input  logic                      cipher_data_out_clear_i,

  // Initial key registers
  output key_init_sel_e             key_init_sel_o,
  output sp2v_e    [NumRegsKey-1:0] key_init_we_o [NumSharesKey],

  // IV registers
  output iv_sel_e                   iv_sel_o,
  output sp2v_e  [NumSlicesCtr-1:0] iv_we_o,

  // Pseudo-random number generator interface
  output logic                      prng_data_req_o,
  input  logic                      prng_data_ack_i,
  output logic                      prng_reseed_req_o,
  input  logic                      prng_reseed_ack_i,

  // Trigger register
  output logic                      start_o,
  output logic                      start_we_o,
  output logic                      key_iv_data_in_clear_o,
  output logic                      key_iv_data_in_clear_we_o,
  output logic                      data_out_clear_o,
  output logic                      data_out_clear_we_o,
  output logic                      prng_reseed_o,
  output logic                      prng_reseed_we_o,

  // Status register
  output logic                      idle_o,
  output logic                      idle_we_o,
  output logic                      stall_o,
  output logic                      stall_we_o,
  input  logic                      output_lost_i,
  output logic                      output_lost_o,
  output logic                      output_lost_we_o,
  output logic                      output_valid_o,
  output logic                      output_valid_we_o,
  output logic                      input_ready_o,
  output logic                      input_ready_we_o
);

  // Optional delay of manual start trigger
  logic start_trigger;

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(AesSecStartTriggerDelayNonDefault, SecStartTriggerDelay == 0)

  if (SecStartTriggerDelay > 0) begin : gen_start_delay
    // Delay the manual start trigger input for SCA measurements.
    localparam int unsigned WidthCounter = $clog2(SecStartTriggerDelay+1);
    logic [WidthCounter-1:0] count_d, count_q;

    // Clear counter when input goes low. Keep value if the specified delay is reached.
    assign count_d = !start_i       ? '0      :
                      start_trigger ? count_q : count_q + 1'b1;
    assign start_trigger = (count_q == SecStartTriggerDelay[WidthCounter-1:0]) ? 1'b1 : 1'b0;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        count_q <= '0;
      end else begin
        count_q <= count_d;
      end
    end

  end else begin : gen_no_start_delay
    // Directly forward the manual start trigger input.
    assign start_trigger = start_i;
  end

  // Signals
  sp2v_e                         ctr_ready;
  sp2v_e      [NumSlicesCtr-1:0] ctr_we;
  sp2v_e                         cipher_in_ready;
  sp2v_e                         cipher_out_valid;
  sp2v_e                         cipher_crypt;
  sp2v_e                         cipher_dec_key_gen;
  logic                          mux_sel_err;
  logic                          mr_err;
  logic                          sp_enc_err;

  // Sparsified FSM signals. These are needed for connecting the individual bits of the Sp2V
  // signals to the single-rail FSMs.
  logic          [Sp2VWidth-1:0] sp_data_out_we;
  logic          [Sp2VWidth-1:0] sp_data_in_prev_we;
  logic          [Sp2VWidth-1:0] sp_ctr_incr;
  logic          [Sp2VWidth-1:0] sp_ctr_ready;
  logic          [Sp2VWidth-1:0] sp_cipher_in_valid;
  logic          [Sp2VWidth-1:0] sp_cipher_in_ready;
  logic          [Sp2VWidth-1:0] sp_cipher_out_valid;
  logic          [Sp2VWidth-1:0] sp_cipher_out_ready;
  logic          [Sp2VWidth-1:0] sp_in_cipher_crypt;
  logic          [Sp2VWidth-1:0] sp_out_cipher_crypt;
  logic          [Sp2VWidth-1:0] sp_in_cipher_dec_key_gen;
  logic          [Sp2VWidth-1:0] sp_out_cipher_dec_key_gen;

  // Multi-rail signals. These are outputs of the single-rail FSMs and need combining.
  logic          [Sp2VWidth-1:0] mr_ctrl_we;
  logic          [Sp2VWidth-1:0] mr_alert;
  logic          [Sp2VWidth-1:0] mr_data_in_we;
  dip_sel_e      [Sp2VWidth-1:0] mr_data_in_prev_sel;
  si_sel_e       [Sp2VWidth-1:0] mr_state_in_sel;
  add_si_sel_e   [Sp2VWidth-1:0] mr_add_state_in_sel;
  add_so_sel_e   [Sp2VWidth-1:0] mr_add_state_out_sel;
  logic          [Sp2VWidth-1:0] mr_cipher_prng_reseed;
  logic          [Sp2VWidth-1:0] mr_cipher_key_clear;
  logic          [Sp2VWidth-1:0] mr_cipher_data_out_clear;
  key_init_sel_e [Sp2VWidth-1:0] mr_key_init_sel;
  iv_sel_e       [Sp2VWidth-1:0] mr_iv_sel;
  logic          [Sp2VWidth-1:0] mr_prng_data_req;
  logic          [Sp2VWidth-1:0] mr_prng_reseed_req;
  logic          [Sp2VWidth-1:0] mr_start_we;
  logic          [Sp2VWidth-1:0] mr_key_iv_data_in_clear_we;
  logic          [Sp2VWidth-1:0] mr_data_out_clear_we;
  logic          [Sp2VWidth-1:0] mr_prng_reseed;
  logic          [Sp2VWidth-1:0] mr_prng_reseed_we;
  logic          [Sp2VWidth-1:0] mr_idle;
  logic          [Sp2VWidth-1:0] mr_idle_we;
  logic          [Sp2VWidth-1:0] mr_stall;
  logic          [Sp2VWidth-1:0] mr_stall_we;
  logic          [Sp2VWidth-1:0] mr_output_lost;
  logic          [Sp2VWidth-1:0] mr_output_lost_we;
  logic          [Sp2VWidth-1:0] mr_output_valid;
  logic          [Sp2VWidth-1:0] mr_output_valid_we;
  logic          [Sp2VWidth-1:0] mr_input_ready;
  logic          [Sp2VWidth-1:0] mr_input_ready_we;

  // To ease interfacing with the individual FSM rails, some signals need to be converted to packed
  // arrays.
  logic [Sp2VWidth-1:0][NumSharesKey-1:0][NumRegsKey-1:0]                int_key_init_we;
  logic                [NumSharesKey-1:0][NumRegsKey-1:0][Sp2VWidth-1:0] log_key_init_we;
  logic                [NumSharesKey-1:0][NumRegsKey-1:0]                int_key_init_qe;
  for (genvar s = 0; s < NumSharesKey; s++) begin : gen_conv_key_init_wqe_shares
    for (genvar i = 0; i < NumRegsKey; i++) begin : gen_conv_key_init_wqe_regs
      assign int_key_init_qe[s][i] = key_init_qe_i[s][i];
      for (genvar j = 0; j < Sp2VWidth; j++) begin : gen_conv_key_init_wqe_log
        assign log_key_init_we[s][i][j] = int_key_init_we[j][s][i];
      end
      assign key_init_we_o[s][i] = sp2v_e'(log_key_init_we[s][i]);
    end
  end
  logic [Sp2VWidth-1:0][NumSlicesCtr-1:0]                int_ctr_we;
  logic                [NumSlicesCtr-1:0][Sp2VWidth-1:0] log_ctr_we;
  logic [Sp2VWidth-1:0][NumSlicesCtr-1:0]                int_iv_we;
  logic                [NumSlicesCtr-1:0][Sp2VWidth-1:0] log_iv_we;
  for (genvar i = 0; i < NumSlicesCtr; i++) begin : gen_conv_ctr_iv_we_slices
    assign log_ctr_we[i] = {ctr_we[i]};
    for (genvar j = 0; j < Sp2VWidth; j++) begin : gen_conv_ctr_iv_we_log
      assign int_ctr_we[j][i] = log_ctr_we[i][j];
      assign log_iv_we[i][j]  = int_iv_we[j][i];
    end
    assign iv_we_o[i] = sp2v_e'(log_iv_we[i]);
  end

  /////////
  // FSM //
  /////////

  // Convert sp2v_e signals to sparsified inputs.
  assign sp_ctr_ready             = {ctr_ready};
  assign sp_cipher_in_ready       = {cipher_in_ready};
  assign sp_cipher_out_valid      = {cipher_out_valid};
  assign sp_in_cipher_crypt       = {cipher_crypt};
  assign sp_in_cipher_dec_key_gen = {cipher_dec_key_gen};

  // SEC_CM: MAIN.FSM.REDUN
  // For every bit in the Sp2V signals, one separate rail is instantiated. The inputs and outputs
  // of every rail are buffered to prevent aggressive synthesis optimizations.
  for (genvar i = 0; i < Sp2VWidth; i++) begin : gen_fsm
    if (SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_fsm_p
      aes_control_fsm_p #(
        .SecMasking ( SecMasking )
      ) u_aes_control_fsm_i (
        .clk_i                     ( clk_i                         ),
        .rst_ni                    ( rst_ni                        ),

        .ctrl_qe_i                 ( ctrl_qe_i                     ),
        .ctrl_we_o                 ( mr_ctrl_we[i]                 ), // AND-combine
        .ctrl_phase_i              ( ctrl_phase_i                  ),
        .ctrl_err_storage_i        ( ctrl_err_storage_i            ),
        .op_i                      ( op_i                          ),
        .mode_i                    ( mode_i                        ),
        .cipher_op_i               ( cipher_op_i                   ),
        .sideload_i                ( sideload_i                    ),
        .prng_reseed_rate_i        ( prng_reseed_rate_i            ),
        .manual_operation_i        ( manual_operation_i            ),
        .key_touch_forces_reseed_i ( key_touch_forces_reseed_i     ),
        .start_i                   ( start_trigger                 ),
        .key_iv_data_in_clear_i    ( key_iv_data_in_clear_i        ),
        .data_out_clear_i          ( data_out_clear_i              ),
        .prng_reseed_i             ( prng_reseed_i                 ),
        .mux_sel_err_i             ( mux_sel_err                   ),
        .sp_enc_err_i              ( sp_enc_err                    ),
        .lc_escalate_en_i          ( lc_escalate_en_i              ),
        .alert_fatal_i             ( alert_fatal_i                 ),
        .alert_o                   ( mr_alert[i]                   ), // OR-combine

        .key_sideload_valid_i      ( key_sideload_valid_i          ),
        .key_init_qe_i             ( int_key_init_qe               ),
        .iv_qe_i                   ( iv_qe_i                       ),
        .data_in_qe_i              ( data_in_qe_i                  ),
        .data_out_re_i             ( data_out_re_i                 ),
        .data_in_we_o              ( mr_data_in_we[i]              ), // AND-combine
        .data_out_we_o             ( sp_data_out_we[i]             ), // Sparsified

        .data_in_prev_sel_o        ( mr_data_in_prev_sel[i]        ), // OR-combine
        .data_in_prev_we_o         ( sp_data_in_prev_we[i]         ), // Sparsified

        .state_in_sel_o            ( mr_state_in_sel[i]            ), // OR-combine
        .add_state_in_sel_o        ( mr_add_state_in_sel[i]        ), // OR-combine
        .add_state_out_sel_o       ( mr_add_state_out_sel[i]       ), // OR-combine

        .ctr_incr_o                ( sp_ctr_incr[i]                ), // Sparsified
        .ctr_ready_i               ( sp_ctr_ready[i]               ), // Sparsified
        .ctr_we_i                  ( int_ctr_we[i]                 ), // Sparsified

        .cipher_in_valid_o         ( sp_cipher_in_valid[i]         ), // Sparsified
        .cipher_in_ready_i         ( sp_cipher_in_ready[i]         ), // Sparsified
        .cipher_out_valid_i        ( sp_cipher_out_valid[i]        ), // Sparsified
        .cipher_out_ready_o        ( sp_cipher_out_ready[i]        ), // Sparsified
        .cipher_crypt_o            ( sp_out_cipher_crypt[i]        ), // Sparsified
        .cipher_crypt_i            ( sp_in_cipher_crypt[i]         ), // Sparsified
        .cipher_dec_key_gen_o      ( sp_out_cipher_dec_key_gen[i]  ), // Sparsified
        .cipher_dec_key_gen_i      ( sp_in_cipher_dec_key_gen[i]   ), // Sparsified
        .cipher_prng_reseed_o      ( mr_cipher_prng_reseed[i]      ), // OR-combine
        .cipher_prng_reseed_i      ( cipher_prng_reseed_i          ),
        .cipher_key_clear_o        ( mr_cipher_key_clear[i]        ), // OR-combine
        .cipher_key_clear_i        ( cipher_key_clear_i            ),
        .cipher_data_out_clear_o   ( mr_cipher_data_out_clear[i]   ), // OR-combine
        .cipher_data_out_clear_i   ( cipher_data_out_clear_i       ),

        .key_init_sel_o            ( mr_key_init_sel[i]            ), // OR-combine
        .key_init_we_o             ( int_key_init_we[i]            ), // Sparsified

        .iv_sel_o                  ( mr_iv_sel[i]                  ), // OR-combine
        .iv_we_o                   ( int_iv_we[i]                  ), // Sparsified

        .prng_data_req_o           ( mr_prng_data_req[i]           ), // OR-combine
        .prng_data_ack_i           ( prng_data_ack_i               ),
        .prng_reseed_req_o         ( mr_prng_reseed_req[i]         ), // OR-combine
        .prng_reseed_ack_i         ( prng_reseed_ack_i             ),

        .start_we_o                ( mr_start_we[i]                ), // OR-combine
        .key_iv_data_in_clear_we_o ( mr_key_iv_data_in_clear_we[i] ), // AND-combine
        .data_out_clear_we_o       ( mr_data_out_clear_we[i]       ), // AND-combine
        .prng_reseed_o             ( mr_prng_reseed[i]             ), // OR-combine
        .prng_reseed_we_o          ( mr_prng_reseed_we[i]          ), // OR-combine

        .idle_o                    ( mr_idle[i]                    ), // AND-combine
        .idle_we_o                 ( mr_idle_we[i]                 ), // AND-combine
        .stall_o                   ( mr_stall[i]                   ), // AND-combine
        .stall_we_o                ( mr_stall_we[i]                ), // AND-combine
        .output_lost_i             ( output_lost_i                 ), // AND-combine
        .output_lost_o             ( mr_output_lost[i]             ), // AND-combine
        .output_lost_we_o          ( mr_output_lost_we[i]          ), // AND-combine
        .output_valid_o            ( mr_output_valid[i]            ), // AND-combine
        .output_valid_we_o         ( mr_output_valid_we[i]         ), // AND-combine
        .input_ready_o             ( mr_input_ready[i]             ), // AND-combine
        .input_ready_we_o          ( mr_input_ready_we[i]          )  // AND-combine
      );
    end else begin : gen_fsm_n
      aes_control_fsm_n #(
        .SecMasking ( SecMasking )
      ) u_aes_control_fsm_i (
        .clk_i                     ( clk_i                         ),
        .rst_ni                    ( rst_ni                        ),

        .ctrl_qe_i                 ( ctrl_qe_i                     ),
        .ctrl_we_o                 ( mr_ctrl_we[i]                 ), // AND-combine
        .ctrl_phase_i              ( ctrl_phase_i                  ),
        .ctrl_err_storage_i        ( ctrl_err_storage_i            ),
        .op_i                      ( op_i                          ),
        .mode_i                    ( mode_i                        ),
        .cipher_op_i               ( cipher_op_i                   ),
        .sideload_i                ( sideload_i                    ),
        .prng_reseed_rate_i        ( prng_reseed_rate_i            ),
        .manual_operation_i        ( manual_operation_i            ),
        .key_touch_forces_reseed_i ( key_touch_forces_reseed_i     ),
        .start_i                   ( start_trigger                 ),
        .key_iv_data_in_clear_i    ( key_iv_data_in_clear_i        ),
        .data_out_clear_i          ( data_out_clear_i              ),
        .prng_reseed_i             ( prng_reseed_i                 ),
        .mux_sel_err_i             ( mux_sel_err                   ),
        .sp_enc_err_i              ( sp_enc_err                    ),
        .lc_escalate_en_i          ( lc_escalate_en_i              ),
        .alert_fatal_i             ( alert_fatal_i                 ),
        .alert_o                   ( mr_alert[i]                   ), // OR-combine

        .key_sideload_valid_i      ( key_sideload_valid_i          ),
        .key_init_qe_i             ( int_key_init_qe               ),
        .iv_qe_i                   ( iv_qe_i                       ),
        .data_in_qe_i              ( data_in_qe_i                  ),
        .data_out_re_i             ( data_out_re_i                 ),
        .data_in_we_o              ( mr_data_in_we[i]              ), // AND-combine
        .data_out_we_no            ( sp_data_out_we[i]             ), // Sparsified

        .data_in_prev_sel_o        ( mr_data_in_prev_sel[i]        ), // OR-combine
        .data_in_prev_we_no        ( sp_data_in_prev_we[i]         ), // Sparsified

        .state_in_sel_o            ( mr_state_in_sel[i]            ), // OR-combine
        .add_state_in_sel_o        ( mr_add_state_in_sel[i]        ), // OR-combine
        .add_state_out_sel_o       ( mr_add_state_out_sel[i]       ), // OR-combine

        .ctr_incr_no               ( sp_ctr_incr[i]                ), // Sparsified
        .ctr_ready_ni              ( sp_ctr_ready[i]               ), // Sparsified
        .ctr_we_ni                 ( int_ctr_we[i]                 ), // Sparsified

        .cipher_in_valid_no        ( sp_cipher_in_valid[i]         ), // Sparsified
        .cipher_in_ready_ni        ( sp_cipher_in_ready[i]         ), // Sparsified
        .cipher_out_valid_ni       ( sp_cipher_out_valid[i]        ), // Sparsified
        .cipher_out_ready_no       ( sp_cipher_out_ready[i]        ), // Sparsified
        .cipher_crypt_no           ( sp_out_cipher_crypt[i]        ), // Sparsified
        .cipher_crypt_ni           ( sp_in_cipher_crypt[i]         ), // Sparsified
        .cipher_dec_key_gen_no     ( sp_out_cipher_dec_key_gen[i]  ), // Sparsified
        .cipher_dec_key_gen_ni     ( sp_in_cipher_dec_key_gen[i]   ), // Sparsified
        .cipher_prng_reseed_o      ( mr_cipher_prng_reseed[i]      ), // OR-combine
        .cipher_prng_reseed_i      ( cipher_prng_reseed_i          ),
        .cipher_key_clear_o        ( mr_cipher_key_clear[i]        ), // OR-combine
        .cipher_key_clear_i        ( cipher_key_clear_i            ),
        .cipher_data_out_clear_o   ( mr_cipher_data_out_clear[i]   ), // OR-combine
        .cipher_data_out_clear_i   ( cipher_data_out_clear_i       ),

        .key_init_sel_o            ( mr_key_init_sel[i]            ), // OR-combine
        .key_init_we_no            ( int_key_init_we[i]            ), // Sparsified

        .iv_sel_o                  ( mr_iv_sel[i]                  ), // OR-combine
        .iv_we_no                  ( int_iv_we[i]                  ), // Sparsified

        .prng_data_req_o           ( mr_prng_data_req[i]           ), // OR-combine
        .prng_data_ack_i           ( prng_data_ack_i               ),
        .prng_reseed_req_o         ( mr_prng_reseed_req[i]         ), // OR-combine
        .prng_reseed_ack_i         ( prng_reseed_ack_i             ),

        .start_we_o                ( mr_start_we[i]                ), // OR-combine
        .key_iv_data_in_clear_we_o ( mr_key_iv_data_in_clear_we[i] ), // AND-combine
        .data_out_clear_we_o       ( mr_data_out_clear_we[i]       ), // AND-combine
        .prng_reseed_o             ( mr_prng_reseed[i]             ), // OR-combine
        .prng_reseed_we_o          ( mr_prng_reseed_we[i]          ), // OR-combine

        .idle_o                    ( mr_idle[i]                    ), // AND-combine
        .idle_we_o                 ( mr_idle_we[i]                 ), // AND-combine
        .stall_o                   ( mr_stall[i]                   ), // AND-combine
        .stall_we_o                ( mr_stall_we[i]                ), // AND-combine
        .output_lost_i             ( output_lost_i                 ), // AND-combine
        .output_lost_o             ( mr_output_lost[i]             ), // AND-combine
        .output_lost_we_o          ( mr_output_lost_we[i]          ), // AND-combine
        .output_valid_o            ( mr_output_valid[i]            ), // AND-combine
        .output_valid_we_o         ( mr_output_valid_we[i]         ), // AND-combine
        .input_ready_o             ( mr_input_ready[i]             ), // AND-combine
        .input_ready_we_o          ( mr_input_ready_we[i]          )  // AND-combine
      );
    end
  end

  // Convert sparsified outputs to sp2v_e type.
  assign data_out_we_o        = sp2v_e'(sp_data_out_we);
  assign data_in_prev_we_o    = sp2v_e'(sp_data_in_prev_we);
  assign ctr_incr_o           = sp2v_e'(sp_ctr_incr);
  assign cipher_in_valid_o    = sp2v_e'(sp_cipher_in_valid);
  assign cipher_out_ready_o   = sp2v_e'(sp_cipher_out_ready);
  assign cipher_crypt_o       = sp2v_e'(sp_out_cipher_crypt);
  assign cipher_dec_key_gen_o = sp2v_e'(sp_out_cipher_dec_key_gen);

  // Combine single-bit FSM outputs.
  // OR: One bit is sufficient to drive the corresponding output bit high.
  assign alert_o                   = |mr_alert;
  assign cipher_prng_reseed_o      = |mr_cipher_prng_reseed;
  assign cipher_key_clear_o        = |mr_cipher_key_clear;
  assign cipher_data_out_clear_o   = |mr_cipher_data_out_clear;
  assign prng_data_req_o           = |mr_prng_data_req;
  assign prng_reseed_req_o         = |mr_prng_reseed_req;
  assign start_we_o                = |mr_start_we;
  assign prng_reseed_o             = |mr_prng_reseed;
  assign prng_reseed_we_o          = |mr_prng_reseed_we;

  // AND: Only if all bits are high, the corresponding action should be triggered.
  assign ctrl_we_o                 = &mr_ctrl_we;
  assign data_in_we_o              = &mr_data_in_we;
  assign key_iv_data_in_clear_we_o = &mr_key_iv_data_in_clear_we;
  assign data_out_clear_we_o       = &mr_data_out_clear_we;
  assign idle_o                    = &mr_idle;
  assign idle_we_o                 = &mr_idle_we;
  assign stall_o                   = &mr_stall;
  assign stall_we_o                = &mr_stall_we;
  assign output_lost_o             = &mr_output_lost;
  assign output_lost_we_o          = &mr_output_lost_we;
  assign output_valid_o            = &mr_output_valid;
  assign output_valid_we_o         = &mr_output_valid_we;
  assign input_ready_o             = &mr_input_ready;
  assign input_ready_we_o          = &mr_input_ready_we;

  // Combine multi-bit, sparse FSM outputs. We simply OR them together. If the FSMs don't provide
  // the same outputs, two cases are possible:
  // - An invalid encoding results: A downstream checker will fire, see mux_sel_err_i.
  // - A valid encoding results: The outputs are compared below to cover this case, see mr_err;
  always_comb begin : combine_sparse_signals
    data_in_prev_sel_o  = dip_sel_e'({DIPSelWidth{1'b0}});
    state_in_sel_o      = si_sel_e'({SISelWidth{1'b0}});
    add_state_in_sel_o  = add_si_sel_e'({AddSISelWidth{1'b0}});
    add_state_out_sel_o = add_so_sel_e'({AddSOSelWidth{1'b0}});
    key_init_sel_o      = key_init_sel_e'({KeyInitSelWidth{1'b0}});
    iv_sel_o            = iv_sel_e'({IVSelWidth{1'b0}});
    mr_err              = 1'b0;

    for (int i = 0; i < Sp2VWidth; i++) begin
      data_in_prev_sel_o  = dip_sel_e'({data_in_prev_sel_o}     | {mr_data_in_prev_sel[i]});
      state_in_sel_o      = si_sel_e'({state_in_sel_o}          | {mr_state_in_sel[i]});
      add_state_in_sel_o  = add_si_sel_e'({add_state_in_sel_o}  | {mr_add_state_in_sel[i]});
      add_state_out_sel_o = add_so_sel_e'({add_state_out_sel_o} | {mr_add_state_out_sel[i]});
      key_init_sel_o      = key_init_sel_e'({key_init_sel_o}    | {mr_key_init_sel[i]});
      iv_sel_o            = iv_sel_e'({iv_sel_o}                | {mr_iv_sel[i]});
    end

    for (int i = 0; i < Sp2VWidth; i++) begin
      if (data_in_prev_sel_o  != mr_data_in_prev_sel[i]  ||
          state_in_sel_o      != mr_state_in_sel[i]      ||
          add_state_in_sel_o  != mr_add_state_in_sel[i]  ||
          add_state_out_sel_o != mr_add_state_out_sel[i] ||
          key_init_sel_o      != mr_key_init_sel[i]      ||
          iv_sel_o            != mr_iv_sel[i]) begin
        mr_err = 1'b1;
      end
    end
  end

  // Collect errors in mux selector signals.
  assign mux_sel_err = mux_sel_err_i | mr_err;

  //////////////////////////////
  // Sparsely Encoded Signals //
  //////////////////////////////

  // SEC_CM: CTRL.SPARSE
  // We use sparse encodings for various critical signals and must ensure that:
  // 1. The synthesis tool doesn't optimize away the sparse encoding.
  // 2. The sparsely encoded signal is always valid. More precisely, an alert or SVA is triggered
  //    if a sparse signal takes on an invalid value.
  // 3. The alert signal remains asserted until reset even if the sparse signal becomes valid again
  //    This is achieved by driving the control FSM into the terminal error state whenever any
  //    sparsely encoded signal becomes invalid.
  //
  // If any sparsely encoded signal becomes invalid, the controller further immediately de-asserts
  // data_out_we_o and other write-enable signals to prevent any data from being released.

  // We use vectors of sparsely encoded signals to reduce code duplication.
  localparam int unsigned NumSp2VSig = 5 + NumSlicesCtr;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig_chk;
  logic  [NumSp2VSig-1:0][Sp2VWidth-1:0] sp2v_sig_chk_raw;
  logic  [NumSp2VSig-1:0]                sp2v_sig_err;

  assign sp2v_sig[0] = cipher_in_ready_i;
  assign sp2v_sig[1] = cipher_out_valid_i;
  assign sp2v_sig[2] = cipher_crypt_i;
  assign sp2v_sig[3] = cipher_dec_key_gen_i;
  assign sp2v_sig[4] = ctr_ready_i;
  for (genvar i = 0; i < NumSlicesCtr; i++) begin : gen_use_ctr_we_i
    assign sp2v_sig[5+i] = ctr_we_i[i];
  end

  // All signals inside sp2v_sig are driven and consumed by multi-rail FSMs.
  localparam bit [NumSp2VSig-1:0] Sp2VEnSecBuf = '0;

  // Individually check sparsely encoded signals.
  for (genvar i = 0; i < NumSp2VSig; i++) begin : gen_sel_buf_chk
    aes_sel_buf_chk #(
      .Num      ( Sp2VNum         ),
      .Width    ( Sp2VWidth       ),
      .EnSecBuf ( Sp2VEnSecBuf[i] )
    ) u_aes_sp2v_sig_buf_chk_i (
      .clk_i  ( clk_i               ),
      .rst_ni ( rst_ni              ),
      .sel_i  ( sp2v_sig[i]         ),
      .sel_o  ( sp2v_sig_chk_raw[i] ),
      .err_o  ( sp2v_sig_err[i]     )
    );
    assign sp2v_sig_chk[i] = sp2v_e'(sp2v_sig_chk_raw[i]);
  end

  assign cipher_in_ready    = sp2v_sig_chk[0];
  assign cipher_out_valid   = sp2v_sig_chk[1];
  assign cipher_crypt       = sp2v_sig_chk[2];
  assign cipher_dec_key_gen = sp2v_sig_chk[3];
  assign ctr_ready          = sp2v_sig_chk[4];
  for (genvar i = 0; i < NumSlicesCtr; i++) begin : gen_ctr_we
    assign ctr_we[i]        = sp2v_sig_chk[5+i];
  end

  // Collect encoding errors.
  // We instantiate the checker modules as close as possible to where the sparsely encoded signals
  // are used. Here, we collect also encoding errors detected in other places of the core.
  assign sp_enc_err = |sp2v_sig_err | sp_enc_err_i;

  //////////////////////
  // Trigger Register //
  //////////////////////
  // Most triggers are only ever cleared by control.
  assign start_o                   = 1'b0;
  assign key_iv_data_in_clear_o    = 1'b0;
  assign data_out_clear_o          = 1'b0;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES main control FSM
//
// This module contains the main control FSM handling the interplay of input/output registers and
// the AES cipher core.

`include "prim_assert.sv"

module aes_control_fsm
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit SecMasking = 0
) (
  input  logic                                    clk_i,
  input  logic                                    rst_ni,

  // Main control signals
  input  logic                                    ctrl_qe_i,
  output logic                                    ctrl_we_o,
  input  logic                                    ctrl_phase_i,
  input  logic                                    ctrl_err_storage_i,
  input  aes_op_e                                 op_i,
  input  aes_mode_e                               mode_i,
  input  ciph_op_e                                cipher_op_i,
  input  logic                                    sideload_i,
  input  prs_rate_e                               prng_reseed_rate_i,
  input  logic                                    manual_operation_i,
  input  logic                                    key_touch_forces_reseed_i,
  input  logic                                    start_i,
  input  logic                                    key_iv_data_in_clear_i,
  input  logic                                    data_out_clear_i,
  input  logic                                    prng_reseed_i,
  input  logic                                    mux_sel_err_i,
  input  logic                                    sp_enc_err_i,
  input  lc_ctrl_pkg::lc_tx_t                     lc_escalate_en_i,
  input  logic                                    alert_fatal_i,
  output logic                                    alert_o,

  // I/O register read/write enables
  input  logic                                    key_sideload_valid_i,
  input  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_qe_i,
  input  logic                    [NumRegsIv-1:0] iv_qe_i,
  input  logic                  [NumRegsData-1:0] data_in_qe_i,
  input  logic                  [NumRegsData-1:0] data_out_re_i,
  output logic                                    data_in_we_o,
  output logic                                    data_out_we_o,           // Sparsify

  // Previous input data register
  output dip_sel_e                                data_in_prev_sel_o,
  output logic                                    data_in_prev_we_o,       // Sparsify

  // Cipher I/O muxes
  output si_sel_e                                 state_in_sel_o,
  output add_si_sel_e                             add_state_in_sel_o,
  output add_so_sel_e                             add_state_out_sel_o,

  // Counter
  output logic                                    ctr_incr_o,              // Sparsify
  input  logic                                    ctr_ready_i,             // Sparsify
  input  logic                 [NumSlicesCtr-1:0] ctr_we_i,                // Sparsify

  // Cipher core control and sync
  output logic                                    cipher_in_valid_o,       // Sparsify
  input  logic                                    cipher_in_ready_i,       // Sparsify
  input  logic                                    cipher_out_valid_i,      // Sparsify
  output logic                                    cipher_out_ready_o,      // Sparsify
  output logic                                    cipher_crypt_o,          // Sparsify
  input  logic                                    cipher_crypt_i,          // Sparsify
  output logic                                    cipher_dec_key_gen_o,    // Sparsify
  input  logic                                    cipher_dec_key_gen_i,    // Sparsify
  output logic                                    cipher_prng_reseed_o,
  input  logic                                    cipher_prng_reseed_i,
  output logic                                    cipher_key_clear_o,
  input  logic                                    cipher_key_clear_i,
  output logic                                    cipher_data_out_clear_o,
  input  logic                                    cipher_data_out_clear_i,

  // Initial key registers
  output key_init_sel_e                           key_init_sel_o,
  output logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_we_o,           // Sparsify

  // IV registers
  output iv_sel_e                                 iv_sel_o,
  output logic                 [NumSlicesCtr-1:0] iv_we_o,                 // Sparsify

  // Pseudo-random number generator interface
  output logic                                    prng_data_req_o,
  input  logic                                    prng_data_ack_i,
  output logic                                    prng_reseed_req_o,
  input  logic                                    prng_reseed_ack_i,

  // Trigger register
  output logic                                    start_we_o,
  output logic                                    key_iv_data_in_clear_we_o,
  output logic                                    data_out_clear_we_o,
  output logic                                    prng_reseed_o,
  output logic                                    prng_reseed_we_o,

  // Status register
  output logic                                    idle_o,
  output logic                                    idle_we_o,
  output logic                                    stall_o,
  output logic                                    stall_we_o,
  input  logic                                    output_lost_i,
  output logic                                    output_lost_o,
  output logic                                    output_lost_we_o,
  output logic                                    output_valid_o,
  output logic                                    output_valid_we_o,
  output logic                                    input_ready_o,
  output logic                                    input_ready_we_o
);

  // Signals
  aes_ctrl_e                aes_ctrl_ns, aes_ctrl_cs;
  logic                     prng_reseed_done_d, prng_reseed_done_q;

  logic                     key_init_clear;
  logic                     key_init_new;
  logic                     key_init_new_pulse;
  logic                     key_init_load;
  logic                     key_init_arm;
  logic                     key_init_ready;
  logic                     key_sideload;

  logic  [NumSlicesCtr-1:0] iv_qe;
  logic                     iv_clear;
  logic                     iv_load;
  logic                     iv_arm;
  logic                     iv_ready;

  logic   [NumRegsData-1:0] data_in_new_d, data_in_new_q;
  logic                     data_in_new;
  logic                     data_in_load;

  logic   [NumRegsData-1:0] data_out_read_d, data_out_read_q;
  logic                     data_out_read;
  logic                     output_valid_q;

  logic                     cfg_valid;
  logic                     no_alert;
  logic                     cipher_op_err;
  logic                     start_common, start_ecb, start_cbc, start_cfb, start_ofb, start_ctr;
  logic                     start;
  logic                     start_core;
  logic                     finish;
  logic                     crypt;
  logic                     cipher_out_done;
  logic                     doing_cbc_enc, doing_cbc_dec;
  logic                     doing_cfb_enc, doing_cfb_dec;
  logic                     doing_ofb;
  logic                     doing_ctr;
  logic                     ctrl_we_q;
  logic                     clear_in_out_status;
  logic                     clear_on_fatal;

  logic                     start_we;
  logic                     key_iv_data_in_clear_we;
  logic                     data_out_clear_we;
  logic                     prng_reseed_we;

  logic                     idle;
  logic                     idle_we;
  logic                     stall;
  logic                     stall_we;
  logic                     output_lost;
  logic                     output_lost_we;
  logic                     output_valid;
  logic                     output_valid_we;
  logic                     input_ready;
  logic                     input_ready_we;

  logic                     block_ctr_expr;
  logic                     block_ctr_decr;

  // Software updates IV in chunks of 32 bits, the counter updates SliceSizeCtr bits at a time.
  // Convert word write enable to internal half-word write enable.
  assign iv_qe = {iv_qe_i[3], iv_qe_i[3], iv_qe_i[2], iv_qe_i[2],
                  iv_qe_i[1], iv_qe_i[1], iv_qe_i[0], iv_qe_i[0]};

  // The cipher core is only ever allowed to start or finish if the control register holds a valid
  // configuration and if no fatal alert condition occured.
  assign cfg_valid = ~((mode_i == AES_NONE) | ctrl_err_storage_i);
  assign no_alert  = ~alert_fatal_i;

  // cipher_op_i is obtained from the configuration of the control register with additional logic.
  assign cipher_op_err = ~(cipher_op_i == CIPH_FWD || cipher_op_i == CIPH_INV);

  // Check common start conditions. These are needed for any mode, unless we are running in
  // manual mode.
  assign start_common = key_init_ready & data_in_new &
      // If key sideload is enabled, we only start if the key is valid.
      (sideload_i ? key_sideload_valid_i : 1'b1);

  // Check mode-specific start conditions. If the IV (and counter) is needed, we only start if
  // also the IV (and counter) is ready.
  assign start_ecb = (mode_i == AES_ECB);
  assign start_cbc = (mode_i == AES_CBC) & iv_ready;
  assign start_cfb = (mode_i == AES_CFB) & iv_ready;
  assign start_ofb = (mode_i == AES_OFB) & iv_ready;
  assign start_ctr = (mode_i == AES_CTR) & iv_ready & ctr_ready_i;

  // If set to start manually, we just wait for the trigger. Otherwise, check common as well as
  // mode-specific start conditions.
  assign start = cfg_valid & no_alert &
      // Manual operation has priority.
      (manual_operation_i ? start_i  :
          // Check start conditions for automatic operation.
          ((start_ecb |
            start_cbc |
            start_cfb |
            start_ofb |
            start_ctr) & start_common));

  // If not set to overwrite data, we wait for any previous output data to be read. data_out_read
  // synchronously clears output_valid_q, unless new output data is written in the exact same
  // clock cycle.
  assign finish = cfg_valid & no_alert &
      // Manual operation has priority.
      (manual_operation_i ? 1'b1 :
          // Make sure previous output data has been read.
          (~output_valid_q | data_out_read));

  // Helper signals for FSM
  assign crypt = cipher_crypt_o | cipher_crypt_i;

  assign doing_cbc_enc = (mode_i == AES_CBC && op_i == AES_ENC) & crypt;
  assign doing_cbc_dec = (mode_i == AES_CBC && op_i == AES_DEC) & crypt;
  assign doing_cfb_enc = (mode_i == AES_CFB && op_i == AES_ENC) & crypt;
  assign doing_cfb_dec = (mode_i == AES_CFB && op_i == AES_DEC) & crypt;
  assign doing_ofb     = (mode_i == AES_OFB)                    & crypt;
  assign doing_ctr     = (mode_i == AES_CTR)                    & crypt;

  // FSM
  always_comb begin : aes_ctrl_fsm

    // Previous input data register control
    data_in_prev_sel_o = DIP_CLEAR;
    data_in_prev_we_o  = 1'b0;

    // Cipher I/O mux control
    state_in_sel_o      = SI_DATA;
    add_state_in_sel_o  = ADD_SI_ZERO;
    add_state_out_sel_o = ADD_SO_ZERO;

    // Counter control
    ctr_incr_o = 1'b0;

    // Cipher core control
    cipher_in_valid_o       = 1'b0;
    cipher_out_ready_o      = 1'b0;
    cipher_out_done         = 1'b0;
    cipher_crypt_o          = 1'b0;
    cipher_dec_key_gen_o    = 1'b0;
    cipher_prng_reseed_o    = 1'b0;
    cipher_key_clear_o      = 1'b0;
    cipher_data_out_clear_o = 1'b0;

    // Initial key registers
    key_init_sel_o = sideload_i ? KEY_INIT_KEYMGR : KEY_INIT_INPUT;
    key_init_we_o = {NumSharesKey * NumRegsKey{1'b0}};

    // IV registers
    iv_sel_o = IV_INPUT;
    iv_we_o  = {NumSlicesCtr{1'b0}};

    // Control register
    ctrl_we_o = 1'b0;

    // Alert
    alert_o = 1'b0;

    // Pseudo-random number generator control
    prng_data_req_o   = 1'b0;
    prng_reseed_req_o = 1'b0;

    // Trigger register control
    start_we                = 1'b0;
    key_iv_data_in_clear_we = 1'b0;
    data_out_clear_we       = 1'b0;
    prng_reseed_we          = 1'b0;

    // Status register
    idle     = 1'b0;
    idle_we  = 1'b0;
    stall    = 1'b0;
    stall_we = 1'b0;

    // Key, data I/O register control
    data_in_load  = 1'b0;
    data_in_we_o  = 1'b0;
    data_out_we_o = 1'b0;

    // Register status tracker control
    key_init_clear = 1'b0;
    key_init_load  = 1'b0;
    key_init_arm   = 1'b0;
    iv_clear       = 1'b0;
    iv_load        = 1'b0;
    iv_arm         = 1'b0;

    // Block counter
    block_ctr_decr = 1'b0;

    // FSM
    aes_ctrl_ns        = aes_ctrl_cs;
    start_core         = 1'b0;
    prng_reseed_done_d = prng_reseed_done_q | prng_reseed_ack_i;

    unique case (aes_ctrl_cs)

      CTRL_IDLE: begin
        // The core is about to start encryption/decryption or another action.
        start_core = start | key_iv_data_in_clear_i | data_out_clear_i | prng_reseed_i;

        // Update status register. A write to the main control register (if sideload is enabled)
        // or writing the last key register can initiate a PRNG reseed operation via trigger
        // register. To avoid that subsequent writes to the main control, key or IV registers
        // collide with the start of the reseed operation, de-assert the idle bit.
        idle    = ~(start_core | (prng_reseed_o & prng_reseed_we_o));
        idle_we = 1'b1;

        // Clear the start trigger when seeing invalid configurations or performing automatic
        // operation.
        start_we = start_i & ((mode_i == AES_NONE) | ~manual_operation_i);

        if (!start_core) begin
          // Initial key and IV updates are ignored if the core is about to start. If key sideload
          // is enabled, software writes to the initial key registers are ignored.
          key_init_we_o = sideload_i ? {NumSharesKey * NumRegsKey{key_sideload}} : key_init_qe_i;
          iv_we_o       = iv_qe;

          // Updates to the control register are only allowed if the core is not about to start and
          // there isn't a storage error. A storage error is unrecoverable and requires a reset.
          ctrl_we_o      = !ctrl_err_storage_i ? ctrl_qe_i : 1'b0;

          // Control register updates clear all register status trackers.
          key_init_clear = ctrl_we_o;
          iv_clear       = ctrl_we_o;
        end

        if (prng_reseed_i) begin
          // PRNG reseeding has highest priority.
          if (!SecMasking) begin
            prng_reseed_done_d = 1'b0;
            aes_ctrl_ns        = CTRL_PRNG_RESEED;
          end else begin
            // In case masking is enabled, also the masking PRNG inside the cipher core needs to
            // be reseeded.
            cipher_prng_reseed_o = 1'b1;

            // Perform handshake.
            cipher_in_valid_o = 1'b1;
            if (cipher_in_ready_i) begin
              prng_reseed_done_d = 1'b0;
              aes_ctrl_ns        = CTRL_PRNG_RESEED;
            end
          end

        end else if (key_iv_data_in_clear_i || data_out_clear_i) begin
          // To clear registers, we must first request fresh pseudo-random data.
          aes_ctrl_ns = CTRL_PRNG_UPDATE;

        end else if (start) begin
          // Signal that we want to start encryption/decryption.
          cipher_crypt_o = 1'b1;

          // Signal if the cipher core shall reseed the masking PRNG.
          cipher_prng_reseed_o = block_ctr_expr;

          // We got a new initial key, but want to do decryption. The cipher core must first
          // generate the start key for decryption.
          cipher_dec_key_gen_o = (cipher_op_i == CIPH_INV) ? key_init_new : 1'b0;

          // Previous input data register control
          data_in_prev_sel_o = doing_cbc_dec ? DIP_DATA_IN :
                               doing_cfb_enc ? DIP_DATA_IN :
                               doing_cfb_dec ? DIP_DATA_IN :
                               doing_ofb     ? DIP_DATA_IN :
                               doing_ctr     ? DIP_DATA_IN : DIP_CLEAR;
          data_in_prev_we_o  = doing_cbc_dec |
                               doing_cfb_enc |
                               doing_cfb_dec |
                               doing_ofb     |
                               doing_ctr;

          // State input mux control
          state_in_sel_o     = doing_cfb_enc ? SI_ZERO :
                               doing_cfb_dec ? SI_ZERO :
                               doing_ofb     ? SI_ZERO :
                               doing_ctr     ? SI_ZERO : SI_DATA;

          // State input additon mux control
          add_state_in_sel_o = doing_cbc_enc ? ADD_SI_IV :
                               doing_cfb_enc ? ADD_SI_IV :
                               doing_cfb_dec ? ADD_SI_IV :
                               doing_ofb     ? ADD_SI_IV :
                               doing_ctr     ? ADD_SI_IV : ADD_SI_ZERO;

          // We have work for the cipher core, perform handshake.
          cipher_in_valid_o = 1'b1;
          if (cipher_in_ready_i) begin
            // Do not yet clear a possible start trigger if we are just starting the generation of
            // the start key for decryption.
            start_we    = ~cipher_dec_key_gen_o;
            aes_ctrl_ns = CTRL_LOAD;
          end
        end
      end

      CTRL_LOAD: begin
        // Signal that we have used the current key, IV, data input to register status tracking.
        key_init_load =  cipher_dec_key_gen_i; // This key is no longer "new", but still clean.
        key_init_arm  = ~cipher_dec_key_gen_i; // The key is still "new", prevent partial updates.
        iv_load       = ~cipher_dec_key_gen_i & (doing_cbc_enc |
                                                 doing_cbc_dec |
                                                 doing_cfb_enc |
                                                 doing_cfb_dec |
                                                 doing_ofb     |
                                                 doing_ctr);
        data_in_load  = ~cipher_dec_key_gen_i;

        // Trigger counter increment.
        ctr_incr_o   = doing_ctr;

        // Unless we are just generating the start key for decryption, we must update the PRNG.
        aes_ctrl_ns  = !cipher_dec_key_gen_i ? CTRL_PRNG_UPDATE : CTRL_FINISH;
      end

      CTRL_PRNG_UPDATE: begin
        // Fresh pseudo-random data is used to:
        // - clear the state in the final cipher round,
        // - clear any other registers in the CLEAR_I/CO states.

        // IV control in case of ongoing encryption/decryption
        // - CTR: IV registers are updated by counter during cipher operation
        iv_sel_o = doing_ctr ? IV_CTR   : IV_INPUT;
        iv_we_o  = doing_ctr ? ctr_we_i : {NumSlicesCtr{1'b0}};

        // Request fresh pseudo-random data, perform handshake.
        prng_data_req_o = 1'b1;
        if (prng_data_ack_i) begin

          // Ongoing encryption/decryption operations have the highest priority. The clear triggers
          // might have become asserted after the handshake with the cipher core.
          if (cipher_crypt_i) begin
            aes_ctrl_ns = CTRL_FINISH;

          end else if (key_iv_data_in_clear_i || data_out_clear_i) begin
            // To clear the output data registers, we re-use the muxing resources of the cipher
            // core. To clear all key material, some key registers inside the cipher core need to
            // be cleared.
            cipher_key_clear_o      = key_iv_data_in_clear_i;
            cipher_data_out_clear_o = data_out_clear_i;

            // We have work for the cipher core, perform handshake.
            cipher_in_valid_o = 1'b1;
            if (cipher_in_ready_i) begin
              aes_ctrl_ns = CTRL_CLEAR_I;
            end
          end else begin
            // Another write to the trigger register must have overwritten the trigger bits that
            // actually caused us to enter this state. Just return.
            aes_ctrl_ns = CTRL_IDLE;
          end // cipher_crypt_i
        end // prng_data_ack_i
      end

      CTRL_PRNG_RESEED: begin
        // Request a reseed of the clearing PRNG.
        prng_reseed_req_o = ~prng_reseed_done_q;

        if (!SecMasking) begin
          if (prng_reseed_done_q) begin
            // Clear the trigger and return.
            prng_reseed_we     = 1'b1;
            prng_reseed_done_d = 1'b0;
            aes_ctrl_ns        = CTRL_IDLE;
          end

        end else begin
          // In case masking is used, we must also wait for the cipher core to reseed the internal
          // masking PRNG. Perform handshake.
          cipher_out_ready_o = prng_reseed_done_q;
          if (cipher_out_ready_o && cipher_out_valid_i) begin
            // Clear the trigger and return.
            prng_reseed_we     = 1'b1;
            prng_reseed_done_d = 1'b0;
            aes_ctrl_ns        = CTRL_IDLE;
          end
        end
      end

      CTRL_FINISH: begin
        // Wait for cipher core to finish.

        if (cipher_dec_key_gen_i) begin
          // We are ready.
          cipher_out_ready_o = 1'b1;
          if (cipher_out_valid_i) begin
            block_ctr_decr = 1'b1;
            aes_ctrl_ns    = CTRL_IDLE;
          end
        end else begin
          // Handshake signals: We are ready once the output data registers can be written. Don't
          // let data propagate in case of mux selector or sparsely encoded signals taking on
          // invalid values.
          cipher_out_ready_o = finish;
          cipher_out_done    = finish & cipher_out_valid_i &
              ~mux_sel_err_i & ~sp_enc_err_i & ~cipher_op_err;

          // Signal if the cipher core is stalled (because previous output has not yet been read).
          stall    = ~finish & cipher_out_valid_i;
          stall_we = 1'b1;

          // State out addition mux control
          add_state_out_sel_o = doing_cbc_dec ? ADD_SO_IV  :
                                doing_cfb_enc ? ADD_SO_DIP :
                                doing_cfb_dec ? ADD_SO_DIP :
                                doing_ofb     ? ADD_SO_DIP :
                                doing_ctr     ? ADD_SO_DIP : ADD_SO_ZERO;

          // IV control
          // - CBC/CFB/OFB: IV registers are only updated when cipher finishes.
          // - CTR: IV registers are updated by counter during cipher operation.
          iv_sel_o = doing_cbc_enc ? IV_DATA_OUT     :
                     doing_cbc_dec ? IV_DATA_IN_PREV :
                     doing_cfb_enc ? IV_DATA_OUT     :
                     doing_cfb_dec ? IV_DATA_IN_PREV :
                     doing_ofb     ? IV_DATA_OUT_RAW :
                     doing_ctr     ? IV_CTR          : IV_INPUT;
          iv_we_o  = doing_cbc_enc ||
                     doing_cbc_dec ||
                     doing_cfb_enc ||
                     doing_cfb_dec ||
                     doing_ofb     ? {NumSlicesCtr{cipher_out_done}} :
                     doing_ctr     ? ctr_we_i                        : {NumSlicesCtr{1'b0}};

          // Arm the IV status tracker: After finishing, the IV registers can be written again
          // by software. We need to make sure software does not partially update the IV.
          iv_arm = (doing_cbc_enc |
                    doing_cbc_dec |
                    doing_cfb_enc |
                    doing_cfb_dec |
                    doing_ofb     |
                    doing_ctr) & cipher_out_done;

          // Proceed upon successful handshake.
          if (cipher_out_done) begin
            block_ctr_decr = 1'b1;
            data_out_we_o  = 1'b1;
            aes_ctrl_ns    = CTRL_IDLE;
          end
        end
      end

      CTRL_CLEAR_I: begin
        // Clear input registers such as Initial Key, IV and input data registers.
        if (key_iv_data_in_clear_i) begin
          // Initial Key
          key_init_sel_o = KEY_INIT_CLEAR;
          key_init_we_o  = {NumSharesKey * NumRegsKey{1'b1}};
          key_init_clear = 1'b1;

          // IV
          iv_sel_o = IV_CLEAR;
          iv_we_o  = {NumSlicesCtr{1'b1}};
          iv_clear = 1'b1;

          // Input data
          data_in_we_o       = 1'b1;
          data_in_prev_sel_o = DIP_CLEAR;
          data_in_prev_we_o  = 1'b1;
        end
        aes_ctrl_ns = CTRL_CLEAR_CO;
      end

      CTRL_CLEAR_CO: begin
        // Wait for cipher core to clear internal Full Key and Decryption Key registers and/or
        // the state register and clear output data registers afterwards.

        // Perform handshake with cipher core.
        cipher_out_ready_o = 1'b1;
        if (cipher_out_valid_i) begin

          // Full Key and Decryption Key registers are cleared by the cipher core.
          // key_iv_data_in_clear_i is acknowledged by the cipher core with cipher_key_clear_i.
          if (cipher_key_clear_i) begin
            // Clear the trigger bit.
            key_iv_data_in_clear_we = 1'b1;
          end

          // To clear the output data registers, we re-use the muxing resources of the cipher core.
          // data_out_clear_i is acknowledged by the cipher core with cipher_data_out_clear_i.
          if (cipher_data_out_clear_i) begin
            // Clear output data and the trigger bit. Don't release data from cipher core in case
            // of mux selector or sparsely encoded signals taking on invalid values.
            data_out_we_o     = ~mux_sel_err_i & ~sp_enc_err_i & ~cipher_op_err;
            data_out_clear_we = 1'b1;
          end

          aes_ctrl_ns = CTRL_IDLE;
        end
      end

      CTRL_ERROR: begin
        // SEC_CM: MAIN.FSM.GLOBAL_ESC
        // SEC_CM: MAIN.FSM.LOCAL_ESC
        // Terminal error state
        alert_o = 1'b1;
      end

      // We should never get here. If we do (e.g. via a malicious glitch), error out immediately.
      default: begin
        aes_ctrl_ns = CTRL_ERROR;
        alert_o = 1'b1;
      end
    endcase

    // Unconditionally jump into the terminal error state in case a mux selector or a sparsely
    // encoded signal becomes invalid, or if the life cycle controller triggers an escalation.
    if (mux_sel_err_i || sp_enc_err_i || cipher_op_err ||
            lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      aes_ctrl_ns = CTRL_ERROR;
    end
  end

  // SEC_CM: MAIN.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, aes_ctrl_ns, aes_ctrl_cs, aes_ctrl_e, CTRL_IDLE)

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_fsm
    if (!rst_ni) begin
      prng_reseed_done_q <= 1'b0;
    end else begin
      prng_reseed_done_q <= prng_reseed_done_d;
    end
  end

  /////////////////////
  // Status Tracking //
  /////////////////////

  // We only take a new sideload key if sideload is enabled, if the provided sideload key is marked
  // as valid, and after the control register has been written for the second time. After that
  // point we don't update the key anymore, as we don't have a notion of when it actually changes.
  // This would be required to trigger decryption key generation for ECB/CBC decryption.
  // To update the sideload key, software has to:
  // 1) wait unitl AES is idle,
  // 2) wait for the key manager to provide the new key,
  // 3) start a new message by writing the control register and providing the IV (if needed).
  assign key_sideload = sideload_i & key_sideload_valid_i & ctrl_we_q & ~ctrl_phase_i;

  // We only use clean initial keys. Either software/counter has updated
  // - all initial key registers, or
  // - none of the initial key registers but the registers were updated in the past.
  aes_reg_status #(
    .Width ( $bits(key_init_we_o) )
  ) u_reg_status_key_init (
    .clk_i       ( clk_i              ),
    .rst_ni      ( rst_ni             ),
    .we_i        ( key_init_we_o      ),
    .use_i       ( key_init_load      ),
    .clear_i     ( key_init_clear     ),
    .arm_i       ( key_init_arm       ),
    .new_o       ( key_init_new       ),
    .new_pulse_o ( key_init_new_pulse ),
    .clean_o     ( key_init_ready     )
  );

  // We only use clean and unused IVs. Either software/counter has updated
  // - all IV registers, or
  // - none of the IV registers but the registers were updated in the past
  // and this particular IV has not yet been used.
  aes_reg_status #(
    .Width ( $bits(iv_we_o) )
  ) u_reg_status_iv (
    .clk_i       ( clk_i    ),
    .rst_ni      ( rst_ni   ),
    .we_i        ( iv_we_o  ),
    .use_i       ( iv_load  ),
    .clear_i     ( iv_clear ),
    .arm_i       ( iv_arm   ),
    .new_o       ( iv_ready ),
    .new_pulse_o (          ),
    .clean_o     (          )
  );

  // Input and output data register status tracking detects if:
  // - A complete new data input block is available, and
  // - An output data block has been read completely.
  // The status tracking needs to be cleared upon writes to the control register. The clearing is
  // applied one cycle later here to avoid zero-latency loops. This additional delay is not
  // relevant as if we are about to start encryption/decryption, we anyway don't allow writes
  // to the control register.
  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_ctrl_we
    if (!rst_ni) begin
      ctrl_we_q <= 1'b0;
    end else begin
      ctrl_we_q <= ctrl_we_o;
    end
  end
  assign clear_in_out_status = ctrl_we_q;

  // Collect writes to data input registers. Cleared if:
  // - data is loaded into cipher core,
  // - clearing data input registers with random data (all data_in_qe_i bits high in next cycle),
  // - clearing the status tracking.
  assign data_in_new_d = data_in_load || &data_in_qe_i || clear_in_out_status ? '0 :
      data_in_new_q | data_in_qe_i;
  assign data_in_new   = &data_in_new_d;

  // Collect reads of data output registers. data_out_read is high for one clock cycle only and
  // clears output_valid_q unless new output is written in the exact same cycle. Cleared if:
  // - clearing data ouput registers with random data,
  // - clearing the status tracking.
  assign data_out_read_d = &data_out_read_q || clear_in_out_status ? '0 :
      data_out_read_q | data_out_re_i;
  assign data_out_read   = &data_out_read_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_edge_detection
    if (!rst_ni) begin
      data_in_new_q   <= '0;
      data_out_read_q <= '0;
    end else begin
      data_in_new_q   <= data_in_new_d;
      data_out_read_q <= data_out_read_d;
    end
  end

  // Status register bits for data input and output
  // Cleared to 1 if:
  // - data is loaded into cipher core,
  // - clearing data input registers with random data,
  // - clearing the status tracking.
  assign input_ready    = ~data_in_new;
  assign input_ready_we =  data_in_new | data_in_load | data_in_we_o | clear_in_out_status;

  // Cleared if:
  // - all data output registers have been read (unless new output is written in the same cycle),
  // - clearing data ouput registers with random data,
  // - clearing the status tracking.
  assign output_valid    = data_out_we_o & ~data_out_clear_we;
  assign output_valid_we = data_out_we_o | data_out_read | data_out_clear_we |
      clear_in_out_status;

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_output_valid
    if (!rst_ni) begin
      output_valid_q <= '0;
    end else if (output_valid_we) begin
      output_valid_q <= output_valid;
    end
  end

  // Output lost status register bit
  // Cleared when updating the Control Register. Set when overwriting previous output data that has
  // not yet been read.
  assign output_lost    = ctrl_we_o     ? 1'b0 :
                          output_lost_i ? 1'b1 : output_valid_q & ~data_out_read;
  assign output_lost_we = ctrl_we_o | data_out_we_o;

  // Should fatal alerts clear the status and trigger register?
  assign clear_on_fatal = ClearStatusOnFatalAlert ? alert_fatal_i : 1'b0;

  /////////////////////
  // Status Register //
  /////////////////////
  assign idle_o            = clear_on_fatal ? 1'b0 : idle;
  assign idle_we_o         = clear_on_fatal ? 1'b1 : idle_we;
  assign stall_o           = clear_on_fatal ? 1'b0 : stall;
  assign stall_we_o        = clear_on_fatal ? 1'b1 : stall_we;
  assign output_lost_o     = clear_on_fatal ? 1'b0 : output_lost;
  assign output_lost_we_o  = clear_on_fatal ? 1'b1 : output_lost_we;
  assign output_valid_o    = clear_on_fatal ? 1'b0 : output_valid;
  assign output_valid_we_o = clear_on_fatal ? 1'b1 : output_valid_we;
  assign input_ready_o     = clear_on_fatal ? 1'b0 : input_ready;
  assign input_ready_we_o  = clear_on_fatal ? 1'b1 : input_ready_we;

  //////////////////////
  // Trigger Register //
  //////////////////////
  // Most triggers are only ever cleared by control. Fatal alerts clear all bits in the trigger
  // register.
  assign start_we_o                = clear_on_fatal ? 1'b1 : start_we;
  assign key_iv_data_in_clear_we_o = clear_on_fatal ? 1'b1 : key_iv_data_in_clear_we;
  assign data_out_clear_we_o       = clear_on_fatal ? 1'b1 : data_out_clear_we;

  // If configured, trigger the reseeding of the PRNGs used for clearing and masking purposes after
  // the key has been updated.
  assign prng_reseed_o    = clear_on_fatal     ? 1'b0 :
                            key_init_new_pulse ? 1'b1 : 1'b0;
  assign prng_reseed_we_o = clear_on_fatal     ? 1'b1                      :
                            key_init_new_pulse ? key_touch_forces_reseed_i : prng_reseed_we;

  ////////////////////////////
  // PRNG Reseeding Counter //
  ////////////////////////////
  // Count the number of blocks since the start of the message to determine when the masking PRNG
  // inside the cipher core needs to be reseeded.
  if (SecMasking) begin : gen_block_ctr
    logic                     block_ctr_set;
    logic [BlockCtrWidth-1:0] block_ctr_d, block_ctr_q;
    logic [BlockCtrWidth-1:0] block_ctr_set_val, block_ctr_decr_val;

    assign block_ctr_expr = block_ctr_q == '0;
    assign block_ctr_set  = ctrl_we_q | (block_ctr_decr & (block_ctr_expr | cipher_prng_reseed_i));

    assign block_ctr_set_val  = prng_reseed_rate_i == PER_1  ? '0                   :
                                prng_reseed_rate_i == PER_64 ? BlockCtrWidth'(63)   :
                                prng_reseed_rate_i == PER_8K ? BlockCtrWidth'(8191) : '0;

    assign block_ctr_decr_val = block_ctr_q - BlockCtrWidth'(1);

    assign block_ctr_d = block_ctr_set  ? block_ctr_set_val  :
                         block_ctr_decr ? block_ctr_decr_val : block_ctr_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin : reg_block_ctr
      if (!rst_ni) begin
        block_ctr_q <= '0;
      end else begin
        block_ctr_q <= block_ctr_d;
      end
    end

  end else begin : gen_no_block_ctr
    assign block_ctr_expr = 1'b0;

    // Tie off unused signals.
    logic      unused_block_ctr_decr;
    prs_rate_e unused_prng_reseed_rate;
    logic      unused_cipher_prng_reseed;
    assign unused_block_ctr_decr     = block_ctr_decr;
    assign unused_prng_reseed_rate   = prng_reseed_rate_i;
    assign unused_cipher_prng_reseed = cipher_prng_reseed_i;
  end

  ////////////////
  // Assertions //
  ////////////////

  // Create a lint error to reduce the risk of accidentally disabling the masking.
  `ASSERT_STATIC_LINT_ERROR(AesControlFsmSecMaskingNonDefault, SecMasking == 1)

  // Selectors must be known/valid
  `ASSERT(AesModeValid, !ctrl_err_storage_i |-> mode_i inside {
      AES_ECB,
      AES_CBC,
      AES_CFB,
      AES_OFB,
      AES_CTR,
      AES_NONE
      })
  `ASSERT(AesOpValid, !ctrl_err_storage_i |-> op_i inside {
      AES_ENC,
      AES_DEC
      })
  `ASSERT(AesCiphOpValid, !cipher_op_err |-> cipher_op_i inside {
      CIPH_FWD,
      CIPH_INV
      })
  `ASSERT(AesControlStateValid, !alert_o |-> aes_ctrl_cs inside {
      CTRL_IDLE,
      CTRL_LOAD,
      CTRL_PRNG_UPDATE,
      CTRL_PRNG_RESEED,
      CTRL_FINISH,
      CTRL_CLEAR_I,
      CTRL_CLEAR_CO
      })

  // Check parameters
  `ASSERT_INIT(AesNumSlicesCtr, NumSlicesCtr == 8)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES main control FSM
//
// This module contains the main control FSM handling the interplay of input/output registers and
// the AES cipher core. This version operates on and produces the positive values of important
// control signals.

`include "prim_assert.sv"

module aes_control_fsm_p
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit SecMasking = 0
) (
  input  logic                                    clk_i,
  input  logic                                    rst_ni,

  // Main control signals
  input  logic                                    ctrl_qe_i,
  output logic                                    ctrl_we_o,
  input  logic                                    ctrl_phase_i,
  input  logic                                    ctrl_err_storage_i,
  input  aes_op_e                                 op_i,
  input  aes_mode_e                               mode_i,
  input  ciph_op_e                                cipher_op_i,
  input  logic                                    sideload_i,
  input  prs_rate_e                               prng_reseed_rate_i,
  input  logic                                    manual_operation_i,
  input  logic                                    key_touch_forces_reseed_i,
  input  logic                                    start_i,
  input  logic                                    key_iv_data_in_clear_i,
  input  logic                                    data_out_clear_i,
  input  logic                                    prng_reseed_i,
  input  logic                                    mux_sel_err_i,
  input  logic                                    sp_enc_err_i,
  input  lc_ctrl_pkg::lc_tx_t                     lc_escalate_en_i,
  input  logic                                    alert_fatal_i,
  output logic                                    alert_o,

  // I/O register read/write enables
  input  logic                                    key_sideload_valid_i,
  input  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_qe_i,
  input  logic                    [NumRegsIv-1:0] iv_qe_i,
  input  logic                  [NumRegsData-1:0] data_in_qe_i,
  input  logic                  [NumRegsData-1:0] data_out_re_i,
  output logic                                    data_in_we_o,
  output logic                                    data_out_we_o,           // Sparsify

  // Previous input data register
  output dip_sel_e                                data_in_prev_sel_o,
  output logic                                    data_in_prev_we_o,       // Sparsify

  // Cipher I/O muxes
  output si_sel_e                                 state_in_sel_o,
  output add_si_sel_e                             add_state_in_sel_o,
  output add_so_sel_e                             add_state_out_sel_o,

  // Counter
  output logic                                    ctr_incr_o,              // Sparsify
  input  logic                                    ctr_ready_i,             // Sparsify
  input  logic                 [NumSlicesCtr-1:0] ctr_we_i,                // Sparsify

  // Cipher core control and sync
  output logic                                    cipher_in_valid_o,       // Sparsify
  input  logic                                    cipher_in_ready_i,       // Sparsify
  input  logic                                    cipher_out_valid_i,      // Sparsify
  output logic                                    cipher_out_ready_o,      // Sparsify
  output logic                                    cipher_crypt_o,          // Sparsify
  input  logic                                    cipher_crypt_i,          // Sparsify
  output logic                                    cipher_dec_key_gen_o,    // Sparsify
  input  logic                                    cipher_dec_key_gen_i,    // Sparsify
  output logic                                    cipher_prng_reseed_o,
  input  logic                                    cipher_prng_reseed_i,
  output logic                                    cipher_key_clear_o,
  input  logic                                    cipher_key_clear_i,
  output logic                                    cipher_data_out_clear_o,
  input  logic                                    cipher_data_out_clear_i,

  // Initial key registers
  output key_init_sel_e                           key_init_sel_o,
  output logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_we_o,           // Sparsify

  // IV registers
  output iv_sel_e                                 iv_sel_o,
  output logic                 [NumSlicesCtr-1:0] iv_we_o,                 // Sparsify

  // Pseudo-random number generator interface
  output logic                                    prng_data_req_o,
  input  logic                                    prng_data_ack_i,
  output logic                                    prng_reseed_req_o,
  input  logic                                    prng_reseed_ack_i,

  // Trigger register
  output logic                                    start_we_o,
  output logic                                    key_iv_data_in_clear_we_o,
  output logic                                    data_out_clear_we_o,
  output logic                                    prng_reseed_o,
  output logic                                    prng_reseed_we_o,

  // Status register
  output logic                                    idle_o,
  output logic                                    idle_we_o,
  output logic                                    stall_o,
  output logic                                    stall_we_o,
  input  logic                                    output_lost_i,
  output logic                                    output_lost_o,
  output logic                                    output_lost_we_o,
  output logic                                    output_valid_o,
  output logic                                    output_valid_we_o,
  output logic                                    input_ready_o,
  output logic                                    input_ready_we_o
);

  /////////////////////
  // Input Buffering //
  /////////////////////

  localparam int NumInBufBits = $bits({
    ctrl_qe_i,
    ctrl_phase_i,
    ctrl_err_storage_i,
    op_i,
    mode_i,
    cipher_op_i,
    sideload_i,
    prng_reseed_rate_i,
    manual_operation_i,
    key_touch_forces_reseed_i,
    start_i,
    key_iv_data_in_clear_i,
    data_out_clear_i,
    prng_reseed_i,
    mux_sel_err_i,
    sp_enc_err_i,
    lc_escalate_en_i,
    alert_fatal_i,
    key_sideload_valid_i,
    key_init_qe_i,
    iv_qe_i,
    data_in_qe_i,
    data_out_re_i,
    ctr_ready_i,
    ctr_we_i,
    cipher_in_ready_i,
    cipher_out_valid_i,
    cipher_crypt_i,
    cipher_dec_key_gen_i,
    cipher_prng_reseed_i,
    cipher_key_clear_i,
    cipher_data_out_clear_i,
    prng_data_ack_i,
    prng_reseed_ack_i,
    output_lost_i
  });

  logic [NumInBufBits-1:0] in, in_buf;

  assign in = {
    ctrl_qe_i,
    ctrl_phase_i,
    ctrl_err_storage_i,
    op_i,
    mode_i,
    cipher_op_i,
    sideload_i,
    prng_reseed_rate_i,
    manual_operation_i,
    key_touch_forces_reseed_i,
    start_i,
    key_iv_data_in_clear_i,
    data_out_clear_i,
    prng_reseed_i,
    mux_sel_err_i,
    sp_enc_err_i,
    lc_escalate_en_i,
    alert_fatal_i,
    key_sideload_valid_i,
    key_init_qe_i,
    iv_qe_i,
    data_in_qe_i,
    data_out_re_i,
    ctr_ready_i,
    ctr_we_i,
    cipher_in_ready_i,
    cipher_out_valid_i,
    cipher_crypt_i,
    cipher_dec_key_gen_i,
    cipher_prng_reseed_i,
    cipher_key_clear_i,
    cipher_data_out_clear_i,
    prng_data_ack_i,
    prng_reseed_ack_i,
    output_lost_i
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumInBufBits)
  ) u_prim_buf_in (
    .in_i(in),
    .out_o(in_buf)
  );

  logic                                    ctrl_qe;
  logic                                    ctrl_phase;
  logic                                    ctrl_err_storage;
  aes_op_e                                 op;
  aes_mode_e                               mode;
  ciph_op_e                                cipher_op;
  logic             [$bits(cipher_op)-1:0] cipher_op_raw;
  logic                                    sideload;
  prs_rate_e                               prng_reseed_rate;
  logic                                    manual_operation;
  logic                                    key_touch_forces_reseed;
  logic                                    start;
  logic                                    key_iv_data_in_clear;
  logic                                    data_out_clear;
  logic                                    prng_reseed_in_buf;
  logic                                    mux_sel_err;
  logic                                    sp_enc_err;
  lc_ctrl_pkg::lc_tx_t                     lc_escalate_en;
  logic                                    alert_fatal;
  logic                                    key_sideload_valid;
  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_qe;
  logic                    [NumRegsIv-1:0] iv_qe;
  logic                  [NumRegsData-1:0] data_in_qe;
  logic                  [NumRegsData-1:0] data_out_re;
  logic                                    ctr_ready;
  logic                 [NumSlicesCtr-1:0] ctr_we;
  logic                                    cipher_in_ready;
  logic                                    cipher_out_valid;
  logic                                    cipher_crypt_in_buf;
  logic                                    cipher_dec_key_gen_in_buf;
  logic                                    cipher_prng_reseed_in_buf;
  logic                                    cipher_key_clear_in_buf;
  logic                                    cipher_data_out_clear_in_buf;
  logic                                    prng_data_ack;
  logic                                    prng_reseed_ack;
  logic                                    output_lost_in_buf;

  assign {ctrl_qe,
          ctrl_phase,
          ctrl_err_storage,
          op,
          mode,
          cipher_op_raw,
          sideload,
          prng_reseed_rate,
          manual_operation,
          key_touch_forces_reseed,
          start,
          key_iv_data_in_clear,
          data_out_clear,
          prng_reseed_in_buf,
          mux_sel_err,
          sp_enc_err,
          lc_escalate_en,
          alert_fatal,
          key_sideload_valid,
          key_init_qe,
          iv_qe,
          data_in_qe,
          data_out_re,
          ctr_ready,
          ctr_we,
          cipher_in_ready,
          cipher_out_valid,
          cipher_crypt_in_buf,
          cipher_dec_key_gen_in_buf,
          cipher_prng_reseed_in_buf,
          cipher_key_clear_in_buf,
          cipher_data_out_clear_in_buf,
          prng_data_ack,
          prng_reseed_ack,
          output_lost_in_buf} = in_buf;

  assign cipher_op = ciph_op_e'(cipher_op_raw);

  // Intermediate output signals
  logic                                    ctrl_we;
  logic                                    alert;
  logic                                    data_in_we;
  logic                                    data_out_we;
  dip_sel_e                                data_in_prev_sel;
  logic                                    data_in_prev_we;
  si_sel_e                                 state_in_sel;
  add_si_sel_e                             add_state_in_sel;
  add_so_sel_e                             add_state_out_sel;
  logic                                    ctr_incr;
  logic                                    cipher_in_valid;
  logic                                    cipher_out_ready;
  logic                                    cipher_crypt_out_buf;
  logic                                    cipher_dec_key_gen_out_buf;
  logic                                    cipher_prng_reseed_out_buf;
  logic                                    cipher_key_clear_out_buf;
  logic                                    cipher_data_out_clear_out_buf;
  key_init_sel_e                           key_init_sel;
  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_we;
  iv_sel_e                                 iv_sel;
  logic                 [NumSlicesCtr-1:0] iv_we;
  logic                                    prng_data_req;
  logic                                    prng_reseed_req;
  logic                                    start_we;
  logic                                    key_iv_data_in_clear_we;
  logic                                    data_out_clear_we;
  logic                                    prng_reseed_out_buf;
  logic                                    prng_reseed_we;
  logic                                    idle;
  logic                                    idle_we;
  logic                                    stall;
  logic                                    stall_we;
  logic                                    output_lost_out_buf;
  logic                                    output_lost_we;
  logic                                    output_valid;
  logic                                    output_valid_we;
  logic                                    input_ready;
  logic                                    input_ready_we;

  /////////////////
  // Regular FSM //
  /////////////////

  aes_control_fsm #(
    .SecMasking ( SecMasking )
  ) u_aes_control_fsm (
    .clk_i                     ( clk_i                         ),
    .rst_ni                    ( rst_ni                        ),

    .ctrl_qe_i                 ( ctrl_qe                       ),
    .ctrl_we_o                 ( ctrl_we                       ),
    .ctrl_phase_i              ( ctrl_phase                    ),
    .ctrl_err_storage_i        ( ctrl_err_storage              ),
    .op_i                      ( op                            ),
    .mode_i                    ( mode                          ),
    .cipher_op_i               ( cipher_op                     ),
    .sideload_i                ( sideload                      ),
    .prng_reseed_rate_i        ( prng_reseed_rate              ),
    .manual_operation_i        ( manual_operation              ),
    .key_touch_forces_reseed_i ( key_touch_forces_reseed       ),
    .start_i                   ( start                         ),
    .key_iv_data_in_clear_i    ( key_iv_data_in_clear          ),
    .data_out_clear_i          ( data_out_clear                ),
    .prng_reseed_i             ( prng_reseed_in_buf            ),
    .mux_sel_err_i             ( mux_sel_err                   ),
    .sp_enc_err_i              ( sp_enc_err                    ),
    .lc_escalate_en_i          ( lc_escalate_en                ),
    .alert_fatal_i             ( alert_fatal                   ),
    .alert_o                   ( alert                         ),

    .key_sideload_valid_i      ( key_sideload_valid            ),
    .key_init_qe_i             ( key_init_qe                   ),
    .iv_qe_i                   ( iv_qe                         ),
    .data_in_qe_i              ( data_in_qe                    ),
    .data_out_re_i             ( data_out_re                   ),
    .data_in_we_o              ( data_in_we                    ),
    .data_out_we_o             ( data_out_we                   ),

    .data_in_prev_sel_o        ( data_in_prev_sel              ),
    .data_in_prev_we_o         ( data_in_prev_we               ),

    .state_in_sel_o            ( state_in_sel                  ),
    .add_state_in_sel_o        ( add_state_in_sel              ),
    .add_state_out_sel_o       ( add_state_out_sel             ),

    .ctr_incr_o                ( ctr_incr                      ),
    .ctr_ready_i               ( ctr_ready                     ),
    .ctr_we_i                  ( ctr_we                        ),

    .cipher_in_valid_o         ( cipher_in_valid               ),
    .cipher_in_ready_i         ( cipher_in_ready               ),
    .cipher_out_valid_i        ( cipher_out_valid              ),
    .cipher_out_ready_o        ( cipher_out_ready              ),
    .cipher_crypt_o            ( cipher_crypt_out_buf          ),
    .cipher_crypt_i            ( cipher_crypt_in_buf           ),
    .cipher_dec_key_gen_o      ( cipher_dec_key_gen_out_buf    ),
    .cipher_dec_key_gen_i      ( cipher_dec_key_gen_in_buf     ),
    .cipher_prng_reseed_o      ( cipher_prng_reseed_out_buf    ),
    .cipher_prng_reseed_i      ( cipher_prng_reseed_in_buf     ),
    .cipher_key_clear_o        ( cipher_key_clear_out_buf      ),
    .cipher_key_clear_i        ( cipher_key_clear_in_buf       ),
    .cipher_data_out_clear_o   ( cipher_data_out_clear_out_buf ),
    .cipher_data_out_clear_i   ( cipher_data_out_clear_in_buf  ),

    .key_init_sel_o            ( key_init_sel                  ),
    .key_init_we_o             ( key_init_we                   ),

    .iv_sel_o                  ( iv_sel                        ),
    .iv_we_o                   ( iv_we                         ),

    .prng_data_req_o           ( prng_data_req                 ),
    .prng_data_ack_i           ( prng_data_ack                 ),
    .prng_reseed_req_o         ( prng_reseed_req               ),
    .prng_reseed_ack_i         ( prng_reseed_ack               ),

    .start_we_o                ( start_we                      ),
    .key_iv_data_in_clear_we_o ( key_iv_data_in_clear_we       ),
    .data_out_clear_we_o       ( data_out_clear_we             ),
    .prng_reseed_o             ( prng_reseed_out_buf           ),
    .prng_reseed_we_o          ( prng_reseed_we                ),

    .idle_o                    ( idle                          ),
    .idle_we_o                 ( idle_we                       ),
    .stall_o                   ( stall                         ),
    .stall_we_o                ( stall_we                      ),
    .output_lost_i             ( output_lost_in_buf            ),
    .output_lost_o             ( output_lost_out_buf           ),
    .output_lost_we_o          ( output_lost_we                ),
    .output_valid_o            ( output_valid                  ),
    .output_valid_we_o         ( output_valid_we               ),
    .input_ready_o             ( input_ready                   ),
    .input_ready_we_o          ( input_ready_we                )
  );

  //////////////////////
  // Output Buffering //
  //////////////////////

  localparam int NumOutBufBits = $bits({
    ctrl_we_o,
    alert_o,
    data_in_we_o,
    data_out_we_o,
    data_in_prev_sel_o,
    data_in_prev_we_o,
    state_in_sel_o,
    add_state_in_sel_o,
    add_state_out_sel_o,
    ctr_incr_o,
    cipher_in_valid_o,
    cipher_out_ready_o,
    cipher_crypt_o,
    cipher_dec_key_gen_o,
    cipher_prng_reseed_o,
    cipher_key_clear_o,
    cipher_data_out_clear_o,
    key_init_sel_o,
    key_init_we_o,
    iv_sel_o,
    iv_we_o,
    prng_data_req_o,
    prng_reseed_req_o,
    start_we_o,
    key_iv_data_in_clear_we_o,
    data_out_clear_we_o,
    prng_reseed_o,
    prng_reseed_we_o,
    idle_o,
    idle_we_o,
    stall_o,
    stall_we_o,
    output_lost_o,
    output_lost_we_o,
    output_valid_o,
    output_valid_we_o,
    input_ready_o,
    input_ready_we_o
  });

  logic [NumOutBufBits-1:0] out, out_buf;

  assign out = {
    ctrl_we,
    alert,
    data_in_we,
    data_out_we,
    data_in_prev_sel,
    data_in_prev_we,
    state_in_sel,
    add_state_in_sel,
    add_state_out_sel,
    ctr_incr,
    cipher_in_valid,
    cipher_out_ready,
    cipher_crypt_out_buf,
    cipher_dec_key_gen_out_buf,
    cipher_prng_reseed_out_buf,
    cipher_key_clear_out_buf,
    cipher_data_out_clear_out_buf,
    key_init_sel,
    key_init_we,
    iv_sel,
    iv_we,
    prng_data_req,
    prng_reseed_req,
    start_we,
    key_iv_data_in_clear_we,
    data_out_clear_we,
    prng_reseed_out_buf,
    prng_reseed_we,
    idle,
    idle_we,
    stall,
    stall_we,
    output_lost_out_buf,
    output_lost_we,
    output_valid,
    output_valid_we,
    input_ready,
    input_ready_we
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumOutBufBits)
  ) u_prim_buf_out (
    .in_i(out),
    .out_o(out_buf)
  );

  assign {ctrl_we_o,
          alert_o,
          data_in_we_o,
          data_out_we_o,
          data_in_prev_sel_o,
          data_in_prev_we_o,
          state_in_sel_o,
          add_state_in_sel_o,
          add_state_out_sel_o,
          ctr_incr_o,
          cipher_in_valid_o,
          cipher_out_ready_o,
          cipher_crypt_o,
          cipher_dec_key_gen_o,
          cipher_prng_reseed_o,
          cipher_key_clear_o,
          cipher_data_out_clear_o,
          key_init_sel_o,
          key_init_we_o,
          iv_sel_o,
          iv_we_o,
          prng_data_req_o,
          prng_reseed_req_o,
          start_we_o,
          key_iv_data_in_clear_we_o,
          data_out_clear_we_o,
          prng_reseed_o,
          prng_reseed_we_o,
          idle_o,
          idle_we_o,
          stall_o,
          stall_we_o,
          output_lost_o,
          output_lost_we_o,
          output_valid_o,
          output_valid_we_o,
          input_ready_o,
          input_ready_we_o} = out_buf;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES main control FSM
//
// This module contains the main control FSM handling the interplay of input/output registers and
// the AES cipher core. This version operates on and produces the negated values of important
// control signals. This is achieved by:
// - instantiating the regular main control FSM operating on and producing the positive values of
//   these signals, and
// - inverting these signals between the regular FSM and the prim_buf synthesis barriers.
// Synthesis tools will then push the inverters into the actual FSM.

`include "prim_assert.sv"

module aes_control_fsm_n
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit SecMasking = 0
) (
  input  logic                                    clk_i,
  input  logic                                    rst_ni,

  // Main control signals
  input  logic                                    ctrl_qe_i,
  output logic                                    ctrl_we_o,
  input  logic                                    ctrl_phase_i,
  input  logic                                    ctrl_err_storage_i,
  input  aes_op_e                                 op_i,
  input  aes_mode_e                               mode_i,
  input  ciph_op_e                                cipher_op_i,
  input  logic                                    sideload_i,
  input  prs_rate_e                               prng_reseed_rate_i,
  input  logic                                    manual_operation_i,
  input  logic                                    key_touch_forces_reseed_i,
  input  logic                                    start_i,
  input  logic                                    key_iv_data_in_clear_i,
  input  logic                                    data_out_clear_i,
  input  logic                                    prng_reseed_i,
  input  logic                                    mux_sel_err_i,
  input  logic                                    sp_enc_err_i,
  input  lc_ctrl_pkg::lc_tx_t                     lc_escalate_en_i,
  input  logic                                    alert_fatal_i,
  output logic                                    alert_o,

  // I/O register read/write enables
  input  logic                                    key_sideload_valid_i,
  input  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_qe_i,
  input  logic                    [NumRegsIv-1:0] iv_qe_i,
  input  logic                  [NumRegsData-1:0] data_in_qe_i,
  input  logic                  [NumRegsData-1:0] data_out_re_i,
  output logic                                    data_in_we_o,
  output logic                                    data_out_we_no,          // Sparsify

  // Previous input data register
  output dip_sel_e                                data_in_prev_sel_o,
  output logic                                    data_in_prev_we_no,      // Sparsify

  // Cipher I/O muxes
  output si_sel_e                                 state_in_sel_o,
  output add_si_sel_e                             add_state_in_sel_o,
  output add_so_sel_e                             add_state_out_sel_o,

  // Counter
  output logic                                    ctr_incr_no,             // Sparsify
  input  logic                                    ctr_ready_ni,            // Sparsify
  input  logic                 [NumSlicesCtr-1:0] ctr_we_ni,               // Sparsify

  // Cipher core control and sync
  output logic                                    cipher_in_valid_no,      // Sparsify
  input  logic                                    cipher_in_ready_ni,      // Sparsify
  input  logic                                    cipher_out_valid_ni,     // Sparsify
  output logic                                    cipher_out_ready_no,     // Sparsify
  output logic                                    cipher_crypt_no,         // Sparsify
  input  logic                                    cipher_crypt_ni,         // Sparsify
  output logic                                    cipher_dec_key_gen_no,   // Sparsify
  input  logic                                    cipher_dec_key_gen_ni,   // Sparsify
  output logic                                    cipher_prng_reseed_o,
  input  logic                                    cipher_prng_reseed_i,
  output logic                                    cipher_key_clear_o,
  input  logic                                    cipher_key_clear_i,
  output logic                                    cipher_data_out_clear_o,
  input  logic                                    cipher_data_out_clear_i,

  // Initial key registers
  output key_init_sel_e                           key_init_sel_o,
  output logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_we_no,          // Sparsify

  // IV registers
  output iv_sel_e                                 iv_sel_o,
  output logic                 [NumSlicesCtr-1:0] iv_we_no,                // Sparsify

  // Pseudo-random number generator interface
  output logic                                    prng_data_req_o,
  input  logic                                    prng_data_ack_i,
  output logic                                    prng_reseed_req_o,
  input  logic                                    prng_reseed_ack_i,

  // Trigger register
  output logic                                    start_we_o,
  output logic                                    key_iv_data_in_clear_we_o,
  output logic                                    data_out_clear_we_o,
  output logic                                    prng_reseed_o,
  output logic                                    prng_reseed_we_o,

  // Status register
  output logic                                    idle_o,
  output logic                                    idle_we_o,
  output logic                                    stall_o,
  output logic                                    stall_we_o,
  input  logic                                    output_lost_i,
  output logic                                    output_lost_o,
  output logic                                    output_lost_we_o,
  output logic                                    output_valid_o,
  output logic                                    output_valid_we_o,
  output logic                                    input_ready_o,
  output logic                                    input_ready_we_o
);

  /////////////////////
  // Input Buffering //
  /////////////////////

  localparam int NumInBufBits = $bits({
    ctrl_qe_i,
    ctrl_phase_i,
    ctrl_err_storage_i,
    op_i,
    mode_i,
    cipher_op_i,
    sideload_i,
    prng_reseed_rate_i,
    manual_operation_i,
    key_touch_forces_reseed_i,
    start_i,
    key_iv_data_in_clear_i,
    data_out_clear_i,
    prng_reseed_i,
    mux_sel_err_i,
    sp_enc_err_i,
    lc_escalate_en_i,
    alert_fatal_i,
    key_sideload_valid_i,
    key_init_qe_i,
    iv_qe_i,
    data_in_qe_i,
    data_out_re_i,
    ctr_ready_ni,
    ctr_we_ni,
    cipher_in_ready_ni,
    cipher_out_valid_ni,
    cipher_crypt_ni,
    cipher_dec_key_gen_ni,
    cipher_prng_reseed_i,
    cipher_key_clear_i,
    cipher_data_out_clear_i,
    prng_data_ack_i,
    prng_reseed_ack_i,
    output_lost_i
  });

  logic [NumInBufBits-1:0] in, in_buf;

  assign in = {
    ctrl_qe_i,
    ctrl_phase_i,
    ctrl_err_storage_i,
    op_i,
    mode_i,
    cipher_op_i,
    sideload_i,
    prng_reseed_rate_i,
    manual_operation_i,
    key_touch_forces_reseed_i,
    start_i,
    key_iv_data_in_clear_i,
    data_out_clear_i,
    prng_reseed_i,
    mux_sel_err_i,
    sp_enc_err_i,
    lc_escalate_en_i,
    alert_fatal_i,
    key_sideload_valid_i,
    key_init_qe_i,
    iv_qe_i,
    data_in_qe_i,
    data_out_re_i,
    ctr_ready_ni,
    ctr_we_ni,
    cipher_in_ready_ni,
    cipher_out_valid_ni,
    cipher_crypt_ni,
    cipher_dec_key_gen_ni,
    cipher_prng_reseed_i,
    cipher_key_clear_i,
    cipher_data_out_clear_i,
    prng_data_ack_i,
    prng_reseed_ack_i,
    output_lost_i
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumInBufBits)
  ) u_prim_buf_in (
    .in_i(in),
    .out_o(in_buf)
  );

  logic                                    ctrl_qe;
  logic                                    ctrl_phase;
  logic                                    ctrl_err_storage;
  aes_op_e                                 op;
  aes_mode_e                               mode;
  ciph_op_e                                cipher_op;
  logic             [$bits(cipher_op)-1:0] cipher_op_raw;
  logic                                    sideload;
  prs_rate_e                               prng_reseed_rate;
  logic                                    manual_operation;
  logic                                    key_touch_forces_reseed;
  logic                                    start;
  logic                                    key_iv_data_in_clear;
  logic                                    data_out_clear;
  logic                                    prng_reseed_in_buf;
  logic                                    mux_sel_err;
  logic                                    sp_enc_err;
  lc_ctrl_pkg::lc_tx_t                     lc_escalate_en;
  logic                                    alert_fatal;
  logic                                    key_sideload_valid;
  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_qe;
  logic                    [NumRegsIv-1:0] iv_qe;
  logic                  [NumRegsData-1:0] data_in_qe;
  logic                  [NumRegsData-1:0] data_out_re;
  logic                                    ctr_ready_n;
  logic                 [NumSlicesCtr-1:0] ctr_we_n;
  logic                                    cipher_in_ready_n;
  logic                                    cipher_out_valid_n;
  logic                                    cipher_crypt_in_buf_n;
  logic                                    cipher_dec_key_gen_in_buf_n;
  logic                                    cipher_prng_reseed_in_buf;
  logic                                    cipher_key_clear_in_buf;
  logic                                    cipher_data_out_clear_in_buf;
  logic                                    prng_data_ack;
  logic                                    prng_reseed_ack;
  logic                                    output_lost_in_buf;

  assign {ctrl_qe,
          ctrl_phase,
          ctrl_err_storage,
          op,
          mode,
          cipher_op_raw,
          sideload,
          prng_reseed_rate,
          manual_operation,
          key_touch_forces_reseed,
          start,
          key_iv_data_in_clear,
          data_out_clear,
          prng_reseed_in_buf,
          mux_sel_err,
          sp_enc_err,
          lc_escalate_en,
          alert_fatal,
          key_sideload_valid,
          key_init_qe,
          iv_qe,
          data_in_qe,
          data_out_re,
          ctr_ready_n,
          ctr_we_n,
          cipher_in_ready_n,
          cipher_out_valid_n,
          cipher_crypt_in_buf_n,
          cipher_dec_key_gen_in_buf_n,
          cipher_prng_reseed_in_buf,
          cipher_key_clear_in_buf,
          cipher_data_out_clear_in_buf,
          prng_data_ack,
          prng_reseed_ack,
          output_lost_in_buf} = in_buf;

  assign cipher_op = ciph_op_e'(cipher_op_raw);

  // Intermediate output signals
  logic                                    ctrl_we;
  logic                                    alert;
  logic                                    data_in_we;
  logic                                    data_out_we;
  dip_sel_e                                data_in_prev_sel;
  logic                                    data_in_prev_we;
  si_sel_e                                 state_in_sel;
  add_si_sel_e                             add_state_in_sel;
  add_so_sel_e                             add_state_out_sel;
  logic                                    ctr_incr;
  logic                                    cipher_in_valid;
  logic                                    cipher_out_ready;
  logic                                    cipher_crypt_out_buf;
  logic                                    cipher_dec_key_gen_out_buf;
  logic                                    cipher_prng_reseed_out_buf;
  logic                                    cipher_key_clear_out_buf;
  logic                                    cipher_data_out_clear_out_buf;
  key_init_sel_e                           key_init_sel;
  logic [NumSharesKey-1:0][NumRegsKey-1:0] key_init_we;
  iv_sel_e                                 iv_sel;
  logic                 [NumSlicesCtr-1:0] iv_we;
  logic                                    prng_data_req;
  logic                                    prng_reseed_req;
  logic                                    start_we;
  logic                                    key_iv_data_in_clear_we;
  logic                                    data_out_clear_we;
  logic                                    prng_reseed_out_buf;
  logic                                    prng_reseed_we;
  logic                                    idle;
  logic                                    idle_we;
  logic                                    stall;
  logic                                    stall_we;
  logic                                    output_lost_out_buf;
  logic                                    output_lost_we;
  logic                                    output_valid;
  logic                                    output_valid_we;
  logic                                    input_ready;
  logic                                    input_ready_we;

  /////////////////
  // Regular FSM //
  /////////////////

  // The regular FSM operates on and produces the positive values of important control signals.
  // Invert *_n input signals here to get the positive values for the regular FSM. To obtain the
  // negated outputs, important output signals are inverted further below. Thanks to the prim_buf
  // synthesis optimization barriers, tools will push the inverters into the regular FSM.
  aes_control_fsm #(
    .SecMasking ( SecMasking )
  ) u_aes_control_fsm (
    .clk_i                     ( clk_i                         ),
    .rst_ni                    ( rst_ni                        ),

    .ctrl_qe_i                 ( ctrl_qe                       ),
    .ctrl_we_o                 ( ctrl_we                       ),
    .ctrl_phase_i              ( ctrl_phase                    ),
    .ctrl_err_storage_i        ( ctrl_err_storage              ),
    .op_i                      ( op                            ),
    .mode_i                    ( mode                          ),
    .cipher_op_i               ( cipher_op                     ),
    .sideload_i                ( sideload                      ),
    .prng_reseed_rate_i        ( prng_reseed_rate              ),
    .manual_operation_i        ( manual_operation              ),
    .key_touch_forces_reseed_i ( key_touch_forces_reseed       ),
    .start_i                   ( start                         ),
    .key_iv_data_in_clear_i    ( key_iv_data_in_clear          ),
    .data_out_clear_i          ( data_out_clear                ),
    .prng_reseed_i             ( prng_reseed_in_buf            ),
    .mux_sel_err_i             ( mux_sel_err                   ),
    .sp_enc_err_i              ( sp_enc_err                    ),
    .lc_escalate_en_i          ( lc_escalate_en                ),
    .alert_fatal_i             ( alert_fatal                   ),
    .alert_o                   ( alert                         ),

    .key_sideload_valid_i      ( key_sideload_valid            ),
    .key_init_qe_i             ( key_init_qe                   ),
    .iv_qe_i                   ( iv_qe                         ),
    .data_in_qe_i              ( data_in_qe                    ),
    .data_out_re_i             ( data_out_re                   ),
    .data_in_we_o              ( data_in_we                    ),
    .data_out_we_o             ( data_out_we                   ), // Invert below for _n output.

    .data_in_prev_sel_o        ( data_in_prev_sel              ),
    .data_in_prev_we_o         ( data_in_prev_we               ), // Invert below for _n output.

    .state_in_sel_o            ( state_in_sel                  ),
    .add_state_in_sel_o        ( add_state_in_sel              ),
    .add_state_out_sel_o       ( add_state_out_sel             ),

    .ctr_incr_o                ( ctr_incr                      ), // Invert below for _n output.
    .ctr_ready_i               ( ~ctr_ready_n                  ), // Invert for regular FSM.
    .ctr_we_i                  ( ~ctr_we_n                     ), // Invert for regular FSM.

    .cipher_in_valid_o         ( cipher_in_valid               ), // Invert below for _n output.
    .cipher_in_ready_i         ( ~cipher_in_ready_n            ), // Invert for regular FSM.
    .cipher_out_valid_i        ( ~cipher_out_valid_n           ), // Invert for regular FSM.
    .cipher_out_ready_o        ( cipher_out_ready              ), // Invert below for _n output.
    .cipher_crypt_o            ( cipher_crypt_out_buf          ), // Invert below for _n output.
    .cipher_crypt_i            ( ~cipher_crypt_in_buf_n        ), // Invert for regular FSM.
    .cipher_dec_key_gen_o      ( cipher_dec_key_gen_out_buf    ), // Invert below for _n output.
    .cipher_dec_key_gen_i      ( ~cipher_dec_key_gen_in_buf_n  ), // Invert for regular FSM.
    .cipher_prng_reseed_o      ( cipher_prng_reseed_out_buf    ),
    .cipher_prng_reseed_i      ( cipher_prng_reseed_in_buf     ),
    .cipher_key_clear_o        ( cipher_key_clear_out_buf      ),
    .cipher_key_clear_i        ( cipher_key_clear_in_buf       ),
    .cipher_data_out_clear_o   ( cipher_data_out_clear_out_buf ),
    .cipher_data_out_clear_i   ( cipher_data_out_clear_in_buf  ),

    .key_init_sel_o            ( key_init_sel                  ),
    .key_init_we_o             ( key_init_we                   ), // Invert below for _n output.

    .iv_sel_o                  ( iv_sel                        ),
    .iv_we_o                   ( iv_we                         ), // Invert below for _n output.

    .prng_data_req_o           ( prng_data_req                 ),
    .prng_data_ack_i           ( prng_data_ack                 ),
    .prng_reseed_req_o         ( prng_reseed_req               ),
    .prng_reseed_ack_i         ( prng_reseed_ack               ),

    .start_we_o                ( start_we                      ),
    .key_iv_data_in_clear_we_o ( key_iv_data_in_clear_we       ),
    .data_out_clear_we_o       ( data_out_clear_we             ),
    .prng_reseed_o             ( prng_reseed_out_buf           ),
    .prng_reseed_we_o          ( prng_reseed_we                ),

    .idle_o                    ( idle                          ),
    .idle_we_o                 ( idle_we                       ),
    .stall_o                   ( stall                         ),
    .stall_we_o                ( stall_we                      ),
    .output_lost_i             ( output_lost_in_buf            ),
    .output_lost_o             ( output_lost_out_buf           ),
    .output_lost_we_o          ( output_lost_we                ),
    .output_valid_o            ( output_valid                  ),
    .output_valid_we_o         ( output_valid_we               ),
    .input_ready_o             ( input_ready                   ),
    .input_ready_we_o          ( input_ready_we                )
  );

  //////////////////////
  // Output Buffering //
  //////////////////////

  localparam int NumOutBufBits = $bits({
    ctrl_we_o,
    alert_o,
    data_in_we_o,
    data_out_we_no,
    data_in_prev_sel_o,
    data_in_prev_we_no,
    state_in_sel_o,
    add_state_in_sel_o,
    add_state_out_sel_o,
    ctr_incr_no,
    cipher_in_valid_no,
    cipher_out_ready_no,
    cipher_crypt_no,
    cipher_dec_key_gen_no,
    cipher_prng_reseed_o,
    cipher_key_clear_o,
    cipher_data_out_clear_o,
    key_init_sel_o,
    key_init_we_no,
    iv_sel_o,
    iv_we_no,
    prng_data_req_o,
    prng_reseed_req_o,
    start_we_o,
    key_iv_data_in_clear_we_o,
    data_out_clear_we_o,
    prng_reseed_o,
    prng_reseed_we_o,
    idle_o,
    idle_we_o,
    stall_o,
    stall_we_o,
    output_lost_o,
    output_lost_we_o,
    output_valid_o,
    output_valid_we_o,
    input_ready_o,
    input_ready_we_o
  });

  logic [NumOutBufBits-1:0] out, out_buf;

  // Important output control signals need to be inverted here. Synthesis tools will push the
  // inverters back into the regular FSM.
  assign out = {
    ctrl_we,
    alert,
    data_in_we,
    ~data_out_we,
    data_in_prev_sel,
    ~data_in_prev_we,
    state_in_sel,
    add_state_in_sel,
    add_state_out_sel,
    ~ctr_incr,
    ~cipher_in_valid,
    ~cipher_out_ready,
    ~cipher_crypt_out_buf,
    ~cipher_dec_key_gen_out_buf,
    cipher_prng_reseed_out_buf,
    cipher_key_clear_out_buf,
    cipher_data_out_clear_out_buf,
    key_init_sel,
    ~key_init_we,
    iv_sel,
    ~iv_we,
    prng_data_req,
    prng_reseed_req,
    start_we,
    key_iv_data_in_clear_we,
    data_out_clear_we,
    prng_reseed_out_buf,
    prng_reseed_we,
    idle,
    idle_we,
    stall,
    stall_we,
    output_lost_out_buf,
    output_lost_we,
    output_valid,
    output_valid_we,
    input_ready,
    input_ready_we
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumOutBufBits)
  ) u_prim_buf_out (
    .in_i(out),
    .out_o(out_buf)
  );

  assign {ctrl_we_o,
          alert_o,
          data_in_we_o,
          data_out_we_no,
          data_in_prev_sel_o,
          data_in_prev_we_no,
          state_in_sel_o,
          add_state_in_sel_o,
          add_state_out_sel_o,
          ctr_incr_no,
          cipher_in_valid_no,
          cipher_out_ready_no,
          cipher_crypt_no,
          cipher_dec_key_gen_no,
          cipher_prng_reseed_o,
          cipher_key_clear_o,
          cipher_data_out_clear_o,
          key_init_sel_o,
          key_init_we_no,
          iv_sel_o,
          iv_we_no,
          prng_data_req_o,
          prng_reseed_req_o,
          start_we_o,
          key_iv_data_in_clear_we_o,
          data_out_clear_we_o,
          prng_reseed_o,
          prng_reseed_we_o,
          idle_o,
          idle_we_o,
          stall_o,
          stall_we_o,
          output_lost_o,
          output_lost_we_o,
          output_valid_o,
          output_valid_we_o,
          input_ready_o,
          input_ready_we_o} = out_buf;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES reg status
//
// This module tracks the collective status of multiple registers.

module aes_reg_status #(
  parameter int Width = 1
) (
  input  logic             clk_i,
  input  logic             rst_ni,

  input  logic [Width-1:0] we_i,
  input  logic             use_i,
  input  logic             clear_i,
  input  logic             arm_i,
  output logic             new_o,
  output logic             new_pulse_o,
  output logic             clean_o
);

  logic [Width-1:0] we_d, we_q;
  logic             armed_d, armed_q;
  logic             all_written;
  logic             none_written;
  logic             new_d, new_q;
  logic             clean_d, clean_q;

  // Collect write operations. Upon clear or use, we start over. If armed, the next write will
  // restart the tracking.
  assign we_d    = (clear_i || use_i) ? '0   :
                   (armed_q && |we_i) ? we_i : (we_q | we_i);
  assign armed_d = (clear_i || use_i) ? 1'b0 :
                   (armed_q && |we_i) ? 1'b0 : armed_q | arm_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_ops
    if (!rst_ni) begin
      we_q    <= '0;
      armed_q <= 1'b0;
    end else begin
      we_q    <= we_d;
      armed_q <= armed_d;
    end
  end

  // Status tracking
  assign all_written  =  &we_d;
  assign none_written = ~|we_d;

  // We have a complete new value if all registers have been written at least once.
  assign new_d   = (clear_i || use_i) ? 1'b0 : all_written;

  // We have a clean value, if either:
  // - all registers have been written at least once, or
  // - no registers have been written but the value was clean previsously.
  // A value is NOT clean, if either:
  // - we get a clear or reset, or
  // - some but not all registers have been written.
  assign clean_d =  clear_i      ? 1'b0    :
                    all_written  ? 1'b1    :
                    none_written ? clean_q : 1'b0;

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_status
    if (!rst_ni) begin
      new_q   <= 1'b0;
      clean_q <= 1'b0;
    end else begin
      new_q   <= new_d;
      clean_q <= clean_d;
    end
  end

  assign new_o       = new_q;
  assign new_pulse_o = new_d & ~new_q;
  assign clean_o     = clean_q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES mux selector buffer and checker
//
// When using sparse encodings for mux selector signals, this module can be used to:
// 1. Prevent aggressive synthesis optimizations on the selector signal, and
// 2. to check that the selector signal is valid, i.e., doesn't take on invalid values.
// Whenever the selector signal takes on an invalid value, an error is signaled.

`include "prim_assert.sv"

module aes_sel_buf_chk #(
  parameter int Num      = 2,
  parameter int Width    = 1,
  parameter bit EnSecBuf = 1'b0
) (
  input  logic             clk_i,  // Used for assertions only.
  input  logic             rst_ni, // Used for assertions only.
  input  logic [Width-1:0] sel_i,
  output logic [Width-1:0] sel_o,
  output logic             err_o
);

  import aes_pkg::*;

  // Tie off unused inputs.
  logic unused_clk;
  logic unused_rst;
  assign unused_clk = clk_i;
  assign unused_rst = rst_ni;

  ////////////
  // Buffer //
  ////////////

  if (EnSecBuf) begin : gen_sec_buf
    prim_sec_anchor_buf #(
      .Width ( Width )
    ) u_prim_buf_sel_i (
      .in_i  ( sel_i ),
      .out_o ( sel_o )
    );
  end else begin : gen_buf
    prim_buf  #(
      .Width ( Width )
    ) u_prim_buf_sel_i (
      .in_i  ( sel_i ),
      .out_o ( sel_o )
    );
  end

  /////////////
  // Checker //
  /////////////

  if (Num == 2) begin : gen_mux2_sel_chk
    // Cast to generic type.
    mux2_sel_e sel_chk;
    assign sel_chk = mux2_sel_e'(sel_o);

    // Actual checker
    always_comb begin : mux2_sel_chk
      unique case (sel_chk)
        MUX2_SEL_0,
        MUX2_SEL_1: err_o = 1'b0;
        default:    err_o = 1'b1;
      endcase
    end

    // Assertion
    `ASSERT(AesMux2SelValid, !err_o |-> sel_chk inside {
        MUX2_SEL_0,
        MUX2_SEL_1
        })

  end else if (Num == 3) begin : gen_mux3_sel_chk
    // Cast to generic type.
    mux3_sel_e sel_chk;
    assign sel_chk = mux3_sel_e'(sel_o);

    // Actual checker
    always_comb begin : mux3_sel_chk
      unique case (sel_chk)
        MUX3_SEL_0,
        MUX3_SEL_1,
        MUX3_SEL_2: err_o = 1'b0;
        default:    err_o = 1'b1;
      endcase
    end

    // Assertion
    `ASSERT(AesMux3SelValid, !err_o |-> sel_chk inside {
        MUX3_SEL_0,
        MUX3_SEL_1,
        MUX3_SEL_2
        })

  end else if (Num == 4) begin : gen_mux4_sel_chk
    // Cast to generic type.
    mux4_sel_e sel_chk;
    assign sel_chk = mux4_sel_e'(sel_o);

    // Actual checker
    always_comb begin : mux4_sel_chk
      unique case (sel_chk)
        MUX4_SEL_0,
        MUX4_SEL_1,
        MUX4_SEL_2,
        MUX4_SEL_3: err_o = 1'b0;
        default:    err_o = 1'b1;
      endcase
    end

    // Assertion
    `ASSERT(AesMux4SelValid, !err_o |-> sel_chk inside {
        MUX4_SEL_0,
        MUX4_SEL_1,
        MUX4_SEL_2,
        MUX4_SEL_3
        })

  end else if (Num == 6) begin : gen_mux6_sel_chk
    // Cast to generic type.
    mux6_sel_e sel_chk;
    assign sel_chk = mux6_sel_e'(sel_o);

    // Actual checker
    always_comb begin : mux6_sel_chk
      unique case (sel_chk)
        MUX6_SEL_0,
        MUX6_SEL_1,
        MUX6_SEL_2,
        MUX6_SEL_3,
        MUX6_SEL_4,
        MUX6_SEL_5: err_o = 1'b0;
        default:    err_o = 1'b1;
      endcase
    end

    // Assertion
    `ASSERT(AesMux6SelValid, !err_o |-> sel_chk inside {
        MUX6_SEL_0,
        MUX6_SEL_1,
        MUX6_SEL_2,
        MUX6_SEL_3,
        MUX6_SEL_4,
        MUX6_SEL_5
        })

  end else begin : gen_width_unsupported
    // Selected width not supported, signal error.
    assign err_o = 1'b1;
  end

  ////////////////
  // Assertions //
  ////////////////

  // We only have generic sparse encodings defined for certain mux input numbers (see aes_pkg.sv).
  `ASSERT_INIT(AesSelBufChkNum, Num inside {2, 3, 4, 6})

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES cipher core implementation
//
// This module contains the AES cipher core including, state register, full key and decryption key
// registers as well as key expand module and control unit.
//
//
// Masking
// -------
//
// If the parameter "Masking" is set to one, first-order masking is applied to the entire
// cipher core including key expand module. For details, see Rivain et al., "Provably secure
// higher-order masking of AES" available at https://eprint.iacr.org/2010/441.pdf .
//
//
// Details on the data formats
// ---------------------------
//
// This implementation uses 4-dimensional SystemVerilog arrays to represent the AES state:
//
//   logic [3:0][3:0][7:0] state_q [NumShares];
//
// The fourth dimension (unpacked) corresponds to the different shares. The first element holds the
// (masked) data share whereas the other elements hold the masks (masked implementation only).
// The three packed dimensions correspond to the 128-bit state matrix per share. This
// implementation uses the same encoding as the Advanced Encryption Standard (AES) FIPS Publication
// 197 available at https://www.nist.gov/publications/advanced-encryption-standard-aes (see Section
// 3.4). An input sequence of 16 bytes (128-bit, left most byte is the first one)
//
//   b0 b1 b2 b3 b4 b5 b6 b7 b8 b9 b10 b11 b12 b13 b14 b15
//
// is mapped to the state matrix as
//
//   [ b0  b4  b8  b12 ]
//   [ b1  b5  b9  b13 ]
//   [ b2  b6  b10 b14 ]
//   [ b3  b7  b11 b15 ] .
//
// This is mapped to three packed dimensions of SystemVerilog array as follows:
// - The first dimension corresponds to the rows. Thus, state_q[0] gives
//   - The first row of the state matrix       [ b0   b4  b8  b12 ], or
//   - A 32-bit packed SystemVerilog array 32h'{ b12, b8, b4, b0  }.
//
// - The second dimension corresponds to the columns. To access complete columns, the state matrix
//   must be transposed first. Thus state_transposed = aes_pkg::aes_transpose(state_q) and then
//   state_transposed[1] gives
//   - The second column of the state matrix   [ b4  b5  b6  b7 ], or
//   - A 32-bit packed SystemVerilog array 32h'{ b7, b6, b5, b4 }.
//
// - The third dimension corresponds to the bytes.
//
// Note that the CSRs are little-endian. The input sequence above is provided to 32-bit DATA_IN_0 -
// DATA_IN_3 registers as
//                   MSB            LSB
// - DATA_IN_0 32h'{ b3 , b2 , b1 , b0  }
// - DATA_IN_1 32h'{ b7 , b6 , b4 , b4  }
// - DATA_IN_2 32h'{ b11, b10, b9 , b8  }
// - DATA_IN_3 32h'{ b15, b14, b13, b12 } .
//
// The input state can thus be obtained by transposing the content of the DATA_IN_0 - DATA_IN_3
// registers.
//
// Similarly, the implementation uses a 3-dimensional array to represent the AES keys:
//
//   logic     [7:0][31:0] key_full_q [NumShares]
//
// The third dimension (unpacked) corresponds to the different shares. The first element holds the
// (masked) key share whereas the other elements hold the masks (masked implementation only).
// The two packed dimensions correspond to the 256-bit key per share. This implementation uses
// the same encoding as the Advanced Encryption Standard (AES) FIPS Publication
// 197 available at https://www.nist.gov/publications/advanced-encryption-standard-aes .
//
// The first packed dimension corresponds to the 8 key words. The second packed dimension
// corresponds to the 32 bits per key word. A key sequence of 32 bytes (256-bit, left most byte is
// the first one)
//
//   b0 b1 b2 b3 b4 b5 b6 b7 b8 b9 b10 b11 b12 b13 b14 b15 ... ... b28 b29 b30 b31
//
// is mapped to the key words and registers (little-endian) as
//                      MSB            LSB
// - KEY_SHARE0_0 32h'{ b3 , b2 , b1 , b0  }
// - KEY_SHARE0_1 32h'{ b7 , b6 , b4 , b4  }
// - KEY_SHARE0_2 32h'{ b11, b10, b9 , b8  }
// - KEY_SHARE0_3 32h'{ b15, b14, b13, b12 }
// - KEY_SHARE0_4 32h'{  .    .    .    .  }
// - KEY_SHARE0_5 32h'{  .    .    .    .  }
// - KEY_SHARE0_6 32h'{  .    .    .    .  }
// - KEY_SHARE0_7 32h'{ b31, b30, b29, b28 } .

`include "prim_assert.sv"

module aes_cipher_core import aes_pkg::*;
#(
  parameter bit          AES192Enable         = 1,
  parameter bit          SecMasking           = 1,
  parameter sbox_impl_e  SecSBoxImpl          = SBoxImplDom,
  parameter bit          SecAllowForcingMasks = 0,
  parameter bit          SecSkipPRNGReseeding = 0,
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,

  localparam int         NumShares            = SecMasking ? 2 : 1, // derived parameter

  parameter masking_lfsr_seed_t RndCnstMaskingLfsrSeed = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t RndCnstMaskingLfsrPerm = RndCnstMaskingLfsrPermDefault
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,

  // Input handshake signals
  input  sp2v_e                       in_valid_i,
  output sp2v_e                       in_ready_o,

  // Output handshake signals
  output sp2v_e                       out_valid_o,
  input  sp2v_e                       out_ready_i,

  // Control and sync signals
  input  logic                        cfg_valid_i, // Used for gating assertions only.
  input  ciph_op_e                    op_i,
  input  key_len_e                    key_len_i,
  input  sp2v_e                       crypt_i,
  output sp2v_e                       crypt_o,
  input  sp2v_e                       dec_key_gen_i,
  output sp2v_e                       dec_key_gen_o,
  input  logic                        prng_reseed_i,
  output logic                        prng_reseed_o,
  input  logic                        key_clear_i,
  output logic                        key_clear_o,
  input  logic                        data_out_clear_i, // Re-use the cipher core muxes.
  output logic                        data_out_clear_o,
  input  logic                        alert_fatal_i,
  output logic                        alert_o,

  // Pseudo-random data for register clearing
  input  logic [WidthPRDClearing-1:0] prd_clearing_i [NumShares],

  // Masking PRNG
  input  logic                        force_masks_i, // Useful for SCA only.
  output logic        [3:0][3:0][7:0] data_in_mask_o,
  output logic                        entropy_req_o,
  input  logic                        entropy_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_i,

  // I/O data & initial key
  input  logic        [3:0][3:0][7:0] state_init_i [NumShares],
  input  logic            [7:0][31:0] key_init_i [NumShares],
  output logic        [3:0][3:0][7:0] state_o [NumShares]
);

  // Signals
  logic               [3:0][3:0][7:0] state_d [NumShares];
  logic               [3:0][3:0][7:0] state_q [NumShares];
  sp2v_e                              state_we_ctrl;
  sp2v_e                              state_we;
  logic           [StateSelWidth-1:0] state_sel_raw;
  state_sel_e                         state_sel_ctrl;
  state_sel_e                         state_sel;
  logic                               state_sel_err;

  sp2v_e                              sub_bytes_en;
  logic                               sub_bytes_prd_we;
  sp2v_e                              sub_bytes_out_req;
  sp2v_e                              sub_bytes_out_ack;
  logic                               sub_bytes_err;
  logic               [3:0][3:0][7:0] sub_bytes_out;
  logic               [3:0][3:0][7:0] sb_in_mask;
  logic               [3:0][3:0][7:0] sb_out_mask;
  logic               [3:0][3:0][7:0] shift_rows_in [NumShares];
  logic               [3:0][3:0][7:0] shift_rows_out [NumShares];
  logic               [3:0][3:0][7:0] mix_columns_out [NumShares];
  logic               [3:0][3:0][7:0] add_round_key_in [NumShares];
  logic               [3:0][3:0][7:0] add_round_key_out [NumShares];
  logic           [AddRKSelWidth-1:0] add_rk_sel_raw;
  add_rk_sel_e                        add_rk_sel_ctrl;
  add_rk_sel_e                        add_rk_sel;
  logic                               add_rk_sel_err;

  logic                   [7:0][31:0] key_full_d [NumShares];
  logic                   [7:0][31:0] key_full_q [NumShares];
  sp2v_e                              key_full_we_ctrl;
  sp2v_e                              key_full_we;
  logic         [KeyFullSelWidth-1:0] key_full_sel_raw;
  key_full_sel_e                      key_full_sel_ctrl;
  key_full_sel_e                      key_full_sel;
  logic                               key_full_sel_err;
  logic                   [7:0][31:0] key_dec_d [NumShares];
  logic                   [7:0][31:0] key_dec_q [NumShares];
  sp2v_e                              key_dec_we_ctrl;
  sp2v_e                              key_dec_we;
  logic          [KeyDecSelWidth-1:0] key_dec_sel_raw;
  key_dec_sel_e                       key_dec_sel_ctrl;
  key_dec_sel_e                       key_dec_sel;
  logic                               key_dec_sel_err;
  logic                   [7:0][31:0] key_expand_out [NumShares];
  ciph_op_e                           key_expand_op;
  sp2v_e                              key_expand_en;
  logic                               key_expand_prd_we;
  sp2v_e                              key_expand_out_req;
  sp2v_e                              key_expand_out_ack;
  logic                               key_expand_err;
  logic                               key_expand_clear;
  logic                         [3:0] key_expand_round;
  logic        [KeyWordsSelWidth-1:0] key_words_sel_raw;
  key_words_sel_e                     key_words_sel_ctrl;
  key_words_sel_e                     key_words_sel;
  logic                               key_words_sel_err;
  logic                   [3:0][31:0] key_words [NumShares];
  logic               [3:0][3:0][7:0] key_bytes [NumShares];
  logic               [3:0][3:0][7:0] key_mix_columns_out [NumShares];
  logic               [3:0][3:0][7:0] round_key [NumShares];
  logic        [RoundKeySelWidth-1:0] round_key_sel_raw;
  round_key_sel_e                     round_key_sel_ctrl;
  round_key_sel_e                     round_key_sel;
  logic                               round_key_sel_err;

  logic                               cfg_valid;
  logic                               mux_sel_err;
  logic                               sp_enc_err_d, sp_enc_err_q;
  logic                               op_err;

  // Pseudo-random data for clearing and masking purposes
  logic                       [127:0] prd_clearing_128 [NumShares];
  logic                       [255:0] prd_clearing_256 [NumShares];

  logic         [WidthPRDMasking-1:0] prd_masking;
  logic  [3:0][3:0][WidthPRDSBox-1:0] prd_sub_bytes;
  logic             [WidthPRDKey-1:0] prd_key_expand;
  logic                               prd_masking_upd;
  logic                               prd_masking_rsd_req;
  logic                               prd_masking_rsd_ack;

  logic               [3:0][3:0][7:0] data_in_mask;

  // Generate clearing signals of appropriate widths. If masking is enabled, the two shares of
  // the registers must be cleared with different pseudo-random data.
  for (genvar s = 0; s < NumShares; s++) begin : gen_prd_clearing_shares
    for (genvar c = 0; c < NumChunksPRDClearing128; c++) begin : gen_prd_clearing_128
      assign prd_clearing_128[s][c * WidthPRDClearing +: WidthPRDClearing] = prd_clearing_i[s];
    end
    for (genvar c = 0; c < NumChunksPRDClearing256; c++) begin : gen_prd_clearing_256
      assign prd_clearing_256[s][c * WidthPRDClearing +: WidthPRDClearing] = prd_clearing_i[s];
    end
  end

  // op_i is one-hot encoded. Check the provided value and trigger an alert upon detecing invalid
  // encodings.
  assign op_err    = ~(op_i == CIPH_FWD || op_i == CIPH_INV);
  assign cfg_valid = cfg_valid_i & ~op_err;

  //////////
  // Data //
  //////////

  // SEC_CM: DATA_REG.SEC_WIPE
  // State registers
  always_comb begin : state_mux
    unique case (state_sel)
      STATE_INIT:  state_d = state_init_i;
      STATE_ROUND: state_d = add_round_key_out;
      STATE_CLEAR: state_d = prd_clearing_128;
      default:     state_d = prd_clearing_128;
    endcase
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : state_reg
    if (!rst_ni) begin
      state_q <= '{default: '0};
    end else if (state_we == SP2V_HIGH) begin
      state_q <= state_d;
    end
  end

  // Masking
  if (!SecMasking) begin : gen_no_masks
    // The masks are ignored anyway, they can be 0.
    assign sb_in_mask  = '0;
    assign prd_masking = '0;

    // Tie-off unused signals.
    logic unused_entropy_ack;
    logic [EntropyWidth-1:0] unused_entropy;
    assign unused_entropy_ack = entropy_ack_i;
    assign unused_entropy     = entropy_i;
    assign entropy_req_o      = 1'b0;

    logic unused_force_masks;
    logic unused_prd_masking_upd;
    logic unused_prd_masking_rsd_req;
    assign unused_force_masks         = force_masks_i;
    assign unused_prd_masking_upd     = prd_masking_upd;
    assign unused_prd_masking_rsd_req = prd_masking_rsd_req;
    assign prd_masking_rsd_ack        = 1'b0;

    logic [3:0][3:0][7:0] unused_sb_out_mask;
    assign unused_sb_out_mask = sb_out_mask;

  end else begin : gen_masks
    // The input mask is the mask share of the state.
    assign sb_in_mask  = state_q[1];

    // The masking PRNG generates:
    // - the pseudo-random data (PRD) required by SubBytes,
    // - the PRD required by the key expand module (has 4 S-Boxes internally).
    aes_prng_masking #(
      .Width                ( WidthPRDMasking        ),
      .ChunkSize            ( ChunkSizePRDMasking    ),
      .EntropyWidth         ( EntropyWidth           ),
      .SecAllowForcingMasks ( SecAllowForcingMasks   ),
      .SecSkipPRNGReseeding ( SecSkipPRNGReseeding   ),
      .RndCnstLfsrSeed      ( RndCnstMaskingLfsrSeed ),
      .RndCnstLfsrPerm      ( RndCnstMaskingLfsrPerm )
    ) u_aes_prng_masking (
      .clk_i         ( clk_i               ),
      .rst_ni        ( rst_ni              ),
      .force_masks_i ( force_masks_i       ),
      .data_update_i ( prd_masking_upd     ),
      .data_o        ( prd_masking         ),
      .reseed_req_i  ( prd_masking_rsd_req ),
      .reseed_ack_o  ( prd_masking_rsd_ack ),
      .entropy_req_o ( entropy_req_o       ),
      .entropy_ack_i ( entropy_ack_i       ),
      .entropy_i     ( entropy_i           )
    );
  end

  // Extract randomness for key expand module and SubBytes.
  //
  // The masking PRNG output has the following shape:
  // prd_masking = { prd_key_expand, prd_sub_bytes }
  assign prd_key_expand = prd_masking[WidthPRDMasking-1 -: WidthPRDKey];
  assign prd_sub_bytes  = prd_masking[WidthPRDData-1 -: WidthPRDData];

  // Extract randomness for masking the input data.
  //
  // The masking PRNG is used for generating both the PRD for the S-Boxes/SubBytes operation as
  // well as for the input data masks. When using any of the masked Canright S-Box implementations,
  // it is important that the SubBytes input masks (generated by the PRNG in Round X-1) and the
  // SubBytes output masks (generated by the PRNG in Round X) are independent. Inside the PRNG,
  // this is achieved by using multiple, separately re-seeded LFSR chunks and by selecting the
  // separate LFSR chunks in alternating fashion. Since the input data masks become the SubBytes
  // input masks in the first round, we select the same 8 bit lanes for the input data masks which
  // are also used to form the SubBytes output mask for the masked Canright S-Box implementations,
  // i.e., the 8 LSBs of the per S-Box PRD. In particular, we have:
  //
  // prd_masking = { prd_key_expand, ... , sb_prd[4], sb_out_mask[4], sb_prd[0], sb_out_mask[0] }
  //
  // Where sb_out_mask[x] contains the SubBytes output mask for byte x (when using a masked
  // Canright S-Box implementation) and sb_prd[x] contains additional PRD consumed by SubBytes for
  // byte x.
  //
  // When using a masked S-Box implementation other than Canright, we still select the 8 LSBs of
  // the per-S-Box PRD to form the input data mask of the corresponding byte. We do this to
  // distribute the input data masks over all LFSR chunks of the masking PRNG. We do the extraction
  // on a row basis.
  localparam int unsigned WidthPRDRow = 4*WidthPRDSBox;
  for (genvar i = 0; i < 4; i++) begin : gen_in_mask
    assign data_in_mask[i] = aes_prd_get_lsbs(prd_masking[i * WidthPRDRow +: WidthPRDRow]);
  end

  // Rotate the data input masks by two LFSR chunks to ensure the data input masks are independent
  // from the PRD fed to the S-Boxes/SubBytes operation.
  assign data_in_mask_o = {data_in_mask[1], data_in_mask[0], data_in_mask[3], data_in_mask[2]};

  // Make sure that whenever the data/mask inputs of the S-Boxes update, the internally buffered
  // PRD is updated in sync.
  assign sub_bytes_prd_we = (state_we == SP2V_HIGH) ? 1'b1 : 1'b0;

  // Cipher data path
  aes_sub_bytes #(
    .SecSBoxImpl ( SecSBoxImpl )
  ) u_aes_sub_bytes (
    .clk_i     ( clk_i             ),
    .rst_ni    ( rst_ni            ),
    .en_i      ( sub_bytes_en      ),
    .prd_we_i  ( sub_bytes_prd_we  ),
    .out_req_o ( sub_bytes_out_req ),
    .out_ack_i ( sub_bytes_out_ack ),
    .op_i      ( op_i              ),
    .data_i    ( state_q[0]        ),
    .mask_i    ( sb_in_mask        ),
    .prd_i     ( prd_sub_bytes     ),
    .data_o    ( sub_bytes_out     ),
    .mask_o    ( sb_out_mask       ),
    .err_o     ( sub_bytes_err     )
  );

  for (genvar s = 0; s < NumShares; s++) begin : gen_shares_shift_mix
    if (s == 0) begin : gen_shift_in_data
      // The (masked) data share
      assign shift_rows_in[s] = sub_bytes_out;
    end else begin : gen_shift_in_mask
      // The mask share
      assign shift_rows_in[s] = sb_out_mask;
    end

    aes_shift_rows u_aes_shift_rows (
      .op_i   ( op_i              ),
      .data_i ( shift_rows_in[s]  ),
      .data_o ( shift_rows_out[s] )
    );

    aes_mix_columns u_aes_mix_columns (
      .op_i   ( op_i               ),
      .data_i ( shift_rows_out[s]  ),
      .data_o ( mix_columns_out[s] )
    );
  end

  always_comb begin : add_round_key_in_mux
    unique case (add_rk_sel)
      ADD_RK_INIT:  add_round_key_in = state_q;
      ADD_RK_ROUND: add_round_key_in = mix_columns_out;
      ADD_RK_FINAL: add_round_key_in = shift_rows_out;
      default:      add_round_key_in = state_q;
    endcase
  end

  for (genvar s = 0; s < NumShares; s++) begin : gen_shares_add_round_key
    assign add_round_key_out[s] = add_round_key_in[s] ^ round_key[s];
  end

  /////////
  // Key //
  /////////

  // SEC_CM: KEY.SEC_WIPE
  // Full Key registers
  always_comb begin : key_full_mux
    unique case (key_full_sel)
      KEY_FULL_ENC_INIT: key_full_d = key_init_i;
      KEY_FULL_DEC_INIT: key_full_d = key_dec_q;
      KEY_FULL_ROUND:    key_full_d = key_expand_out;
      KEY_FULL_CLEAR:    key_full_d = prd_clearing_256;
      default:           key_full_d = prd_clearing_256;
    endcase
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : key_full_reg
    if (!rst_ni) begin
      key_full_q <= '{default: '0};
    end else if (key_full_we == SP2V_HIGH) begin
      key_full_q <= key_full_d;
    end
  end

  // SEC_CM: KEY.SEC_WIPE
  // Decryption Key registers
  always_comb begin : key_dec_mux
    unique case (key_dec_sel)
      KEY_DEC_EXPAND: key_dec_d = key_expand_out;
      KEY_DEC_CLEAR:  key_dec_d = prd_clearing_256;
      default:        key_dec_d = prd_clearing_256;
    endcase
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : key_dec_reg
    if (!rst_ni) begin
      key_dec_q <= '{default: '0};
    end else if (key_dec_we == SP2V_HIGH) begin
      key_dec_q <= key_dec_d;
    end
  end

  // Make sure that whenever the data/mask inputs of the S-Boxes update, the internally buffered
  // PRD is updated in sync.
  assign key_expand_prd_we = (key_full_we == SP2V_HIGH) ? 1'b1 : 1'b0;

  // Key expand data path
  aes_key_expand #(
    .AES192Enable ( AES192Enable ),
    .SecMasking   ( SecMasking   ),
    .SecSBoxImpl  ( SecSBoxImpl  )
  ) u_aes_key_expand (
    .clk_i       ( clk_i              ),
    .rst_ni      ( rst_ni             ),
    .cfg_valid_i ( cfg_valid          ),
    .op_i        ( key_expand_op      ),
    .en_i        ( key_expand_en      ),
    .prd_we_i    ( key_expand_prd_we  ),
    .out_req_o   ( key_expand_out_req ),
    .out_ack_i   ( key_expand_out_ack ),
    .clear_i     ( key_expand_clear   ),
    .round_i     ( key_expand_round   ),
    .key_len_i   ( key_len_i          ),
    .key_i       ( key_full_q         ),
    .key_o       ( key_expand_out     ),
    .prd_i       ( prd_key_expand     ),
    .err_o       ( key_expand_err     )
  );

  for (genvar s = 0; s < NumShares; s++) begin : gen_shares_round_key
    always_comb begin : key_words_mux
      unique case (key_words_sel)
        KEY_WORDS_0123: key_words[s] = key_full_q[s][3:0];
        KEY_WORDS_2345: key_words[s] = AES192Enable ? key_full_q[s][5:2] : '0;
        KEY_WORDS_4567: key_words[s] = key_full_q[s][7:4];
        KEY_WORDS_ZERO: key_words[s] = '0;
        default:        key_words[s] = '0;
      endcase
    end

    // Convert words to bytes (every key word contains one column).
    assign key_bytes[s] = aes_transpose(key_words[s]);

    aes_mix_columns u_aes_key_mix_columns (
      .op_i   ( CIPH_INV               ),
      .data_i ( key_bytes[s]           ),
      .data_o ( key_mix_columns_out[s] )
    );
  end

  always_comb begin : round_key_mux
    unique case (round_key_sel)
      ROUND_KEY_DIRECT: round_key = key_bytes;
      ROUND_KEY_MIXED:  round_key = key_mix_columns_out;
      default:          round_key = key_bytes;
    endcase
  end

  /////////////
  // Control //
  /////////////

  // Control
  aes_cipher_control #(
    .SecMasking  ( SecMasking  ),
    .SecSBoxImpl ( SecSBoxImpl )
  ) u_aes_cipher_control (
    .clk_i                ( clk_i               ),
    .rst_ni               ( rst_ni              ),

    .in_valid_i           ( in_valid_i          ),
    .in_ready_o           ( in_ready_o          ),

    .out_valid_o          ( out_valid_o         ),
    .out_ready_i          ( out_ready_i         ),

    .cfg_valid_i          ( cfg_valid           ),
    .op_i                 ( op_i                ),
    .key_len_i            ( key_len_i           ),
    .crypt_i              ( crypt_i             ),
    .crypt_o              ( crypt_o             ),
    .dec_key_gen_i        ( dec_key_gen_i       ),
    .dec_key_gen_o        ( dec_key_gen_o       ),
    .prng_reseed_i        ( prng_reseed_i       ),
    .prng_reseed_o        ( prng_reseed_o       ),
    .key_clear_i          ( key_clear_i         ),
    .key_clear_o          ( key_clear_o         ),
    .data_out_clear_i     ( data_out_clear_i    ),
    .data_out_clear_o     ( data_out_clear_o    ),
    .mux_sel_err_i        ( mux_sel_err         ),
    .sp_enc_err_i         ( sp_enc_err_q        ),
    .op_err_i             ( op_err              ),
    .alert_fatal_i        ( alert_fatal_i       ),
    .alert_o              ( alert_o             ),

    .prng_update_o        ( prd_masking_upd     ),
    .prng_reseed_req_o    ( prd_masking_rsd_req ),
    .prng_reseed_ack_i    ( prd_masking_rsd_ack ),

    .state_sel_o          ( state_sel_ctrl      ),
    .state_we_o           ( state_we_ctrl       ),
    .sub_bytes_en_o       ( sub_bytes_en        ),
    .sub_bytes_out_req_i  ( sub_bytes_out_req   ),
    .sub_bytes_out_ack_o  ( sub_bytes_out_ack   ),
    .add_rk_sel_o         ( add_rk_sel_ctrl     ),

    .key_expand_op_o      ( key_expand_op       ),
    .key_full_sel_o       ( key_full_sel_ctrl   ),
    .key_full_we_o        ( key_full_we_ctrl    ),
    .key_dec_sel_o        ( key_dec_sel_ctrl    ),
    .key_dec_we_o         ( key_dec_we_ctrl     ),
    .key_expand_en_o      ( key_expand_en       ),
    .key_expand_out_req_i ( key_expand_out_req  ),
    .key_expand_out_ack_o ( key_expand_out_ack  ),
    .key_expand_clear_o   ( key_expand_clear    ),
    .key_expand_round_o   ( key_expand_round    ),
    .key_words_sel_o      ( key_words_sel_ctrl  ),
    .round_key_sel_o      ( round_key_sel_ctrl  )
  );

  ///////////////
  // Selectors //
  ///////////////

  // We use sparse encodings for these mux selector signals and must ensure that:
  // 1. The synthesis tool doesn't optimize away the sparse encoding.
  // 2. The selector signal is always valid. More precisely, an alert or SVA is triggered if a
  //    selector signal takes on an invalid value.
  // 3. The alert signal remains asserted until reset even if the selector signal becomes valid
  //    again. This is achieved by driving the control FSM into the terminal error state whenever
  //    any mux selector signal becomes invalid.
  //
  // If any mux selector signal becomes invalid, the cipher core further immediately de-asserts
  // the out_valid_o signal to prevent any data from being released.

  aes_sel_buf_chk #(
    .Num      ( StateSelNum   ),
    .Width    ( StateSelWidth ),
    .EnSecBuf ( 1'b1          )
  ) u_aes_state_sel_buf_chk (
    .clk_i  ( clk_i          ),
    .rst_ni ( rst_ni         ),
    .sel_i  ( state_sel_ctrl ),
    .sel_o  ( state_sel_raw  ),
    .err_o  ( state_sel_err  )
  );
  assign state_sel = state_sel_e'(state_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( AddRKSelNum   ),
    .Width    ( AddRKSelWidth ),
    .EnSecBuf ( 1'b1          )
  ) u_aes_add_rk_sel_buf_chk (
    .clk_i  ( clk_i           ),
    .rst_ni ( rst_ni          ),
    .sel_i  ( add_rk_sel_ctrl ),
    .sel_o  ( add_rk_sel_raw  ),
    .err_o  ( add_rk_sel_err  )
  );
  assign add_rk_sel = add_rk_sel_e'(add_rk_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( KeyFullSelNum   ),
    .Width    ( KeyFullSelWidth ),
    .EnSecBuf ( 1'b1            )
  ) u_aes_key_full_sel_buf_chk (
    .clk_i  ( clk_i             ),
    .rst_ni ( rst_ni            ),
    .sel_i  ( key_full_sel_ctrl ),
    .sel_o  ( key_full_sel_raw  ),
    .err_o  ( key_full_sel_err  )
  );
  assign key_full_sel = key_full_sel_e'(key_full_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( KeyDecSelNum   ),
    .Width    ( KeyDecSelWidth ),
    .EnSecBuf ( 1'b1           )
  ) u_aes_key_dec_sel_buf_chk (
    .clk_i  ( clk_i            ),
    .rst_ni ( rst_ni           ),
    .sel_i  ( key_dec_sel_ctrl ),
    .sel_o  ( key_dec_sel_raw  ),
    .err_o  ( key_dec_sel_err  )
  );
  assign key_dec_sel = key_dec_sel_e'(key_dec_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( KeyWordsSelNum   ),
    .Width    ( KeyWordsSelWidth ),
    .EnSecBuf ( 1'b1             )
  ) u_aes_key_words_sel_buf_chk (
    .clk_i  ( clk_i              ),
    .rst_ni ( rst_ni             ),
    .sel_i  ( key_words_sel_ctrl ),
    .sel_o  ( key_words_sel_raw  ),
    .err_o  ( key_words_sel_err  )
  );
  assign key_words_sel = key_words_sel_e'(key_words_sel_raw);

  aes_sel_buf_chk #(
    .Num      ( RoundKeySelNum   ),
    .Width    ( RoundKeySelWidth ),
    .EnSecBuf ( 1'b1             )
  ) u_aes_round_key_sel_buf_chk (
    .clk_i  ( clk_i              ),
    .rst_ni ( rst_ni             ),
    .sel_i  ( round_key_sel_ctrl ),
    .sel_o  ( round_key_sel_raw  ),
    .err_o  ( round_key_sel_err  )
  );
  assign round_key_sel = round_key_sel_e'(round_key_sel_raw);

  // Signal invalid mux selector signals to control FSM which will lock up and trigger an alert.
  assign mux_sel_err = state_sel_err | add_rk_sel_err | key_full_sel_err |
      key_dec_sel_err | key_words_sel_err | round_key_sel_err;

  //////////////////////////////
  // Sparsely Encoded Signals //
  //////////////////////////////

  // We use sparse encodings for various critical signals and must ensure that:
  // 1. The synthesis tool doesn't optimize away the sparse encoding.
  // 2. The sparsely encoded signal is always valid. More precisely, an alert or SVA is triggered
  //    if a sparse signal takes on an invalid value.
  // 3. The alert signal remains asserted until reset even if the sparse signal becomes valid again
  //    This is achieved by driving the control FSM into the terminal error state whenever any
  //    sparsely encoded signal becomes invalid.
  //
  // If any sparsely encoded signal becomes invalid, the cipher core further immediately de-asserts
  // the out_valid_o signal to prevent any data from being released.

  // We use vectors of sparsely encoded signals to reduce code duplication.
  localparam int unsigned NumSp2VSig = 3;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig_chk;
  logic  [NumSp2VSig-1:0][Sp2VWidth-1:0] sp2v_sig_chk_raw;
  logic  [NumSp2VSig-1:0]                sp2v_sig_err;

  assign sp2v_sig[0] = state_we_ctrl;
  assign sp2v_sig[1] = key_full_we_ctrl;
  assign sp2v_sig[2] = key_dec_we_ctrl;

  // All signals inside sp2v_sig are eventually converted to single-rail signals.
  localparam bit [NumSp2VSig-1:0] Sp2VEnSecBuf = {NumSp2VSig{1'b1}};

  // Individually check sparsely encoded signals.
  for (genvar i = 0; i < NumSp2VSig; i++) begin : gen_sel_buf_chk
    aes_sel_buf_chk #(
      .Num      ( Sp2VNum         ),
      .Width    ( Sp2VWidth       ),
      .EnSecBuf ( Sp2VEnSecBuf[i] )
    ) u_aes_sp2v_sig_buf_chk_i (
      .clk_i  ( clk_i               ),
      .rst_ni ( rst_ni              ),
      .sel_i  ( sp2v_sig[i]         ),
      .sel_o  ( sp2v_sig_chk_raw[i] ),
      .err_o  ( sp2v_sig_err[i]     )
    );
    assign sp2v_sig_chk[i] = sp2v_e'(sp2v_sig_chk_raw[i]);
  end

  assign state_we    = sp2v_sig_chk[0];
  assign key_full_we = sp2v_sig_chk[1];
  assign key_dec_we  = sp2v_sig_chk[2];

  // Collect encoding errors.
  // We instantiate the checker modules as close as possible to where the sparsely encoded signals
  // are used. Here, we collect also encoding errors detected in other places of the cipher core.
  assign sp_enc_err_d = |sp2v_sig_err | sub_bytes_err | key_expand_err;

  // We need to register the collected error signal to avoid circular loops in the cipher core
  // controller related to out_valid_o and detecting errors in state_we_o and sub_bytes_out_ack.
  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_sp_enc_err
    if (!rst_ni) begin
      sp_enc_err_q <= 1'b0;
    end else if (sp_enc_err_d) begin
      sp_enc_err_q <= 1'b1;
    end
  end

  /////////////
  // Outputs //
  /////////////

  // The output of the last round is not stored into the state register but forwarded directly.
  assign state_o = add_round_key_out;

  ////////////////
  // Assertions //
  ////////////////

// Typically assertions already contain this macro, which ensures that assertions are only compiled
// in simulation and FPV. However, we wrap the entire assertion section with INC_ASSERT so that the
// helper logic below is not synthesized either, since that could cause issues in DC.
`ifdef INC_ASSERT
  //VCS coverage off
  // pragma coverage off

  // Create a lint error to reduce the risk of accidentally disabling the masking.
  `ASSERT_STATIC_LINT_ERROR(AesSecMaskingNonDefault, SecMasking == 1)

  // Cipher core masking requires a masked SBox and vice versa.
  `ASSERT_INIT(AesMaskedCoreAndSBox,
      (SecMasking &&
      (SecSBoxImpl == SBoxImplCanrightMasked ||
       SecSBoxImpl == SBoxImplCanrightMaskedNoreuse ||
       SecSBoxImpl == SBoxImplDom)) ||
      (!SecMasking &&
      (SecSBoxImpl == SBoxImplLut ||
       SecSBoxImpl == SBoxImplCanright)))

  // Signals used for assertions only.
  logic prd_clearing_equals_output, unused_prd_clearing_equals_output;
  assign prd_clearing_equals_output = (prd_clearing_128 == add_round_key_out);
  assign unused_prd_clearing_equals_output = prd_clearing_equals_output;

  // Ensure that the state register gets cleared with pseudo-random data at the end of the last
  // round. The following two scenarios are unlikely but not illegal:
  // 1. The newly loaded initial state matches the previous output (the round counter is only
  //    cleared upon loading the new initial state).
  // 2. The previous pseudo-random data is equal to the previous output.
  // Otherwise, we must see an alert e.g. because the state multiplexer got glitched.
  `ASSERT(AesSecCmDataRegKeySca, (state_we == SP2V_HIGH) &&
      ((key_len_i == AES_128 && u_aes_cipher_control.rnd_ctr == 4'd10) ||
       (key_len_i == AES_192 && u_aes_cipher_control.rnd_ctr == 4'd12) ||
       (key_len_i == AES_256 && u_aes_cipher_control.rnd_ctr == 4'd14)) |=>
      (state_q != $past(add_round_key_out)) ||
      (state_q == $past(state_init_i)) ||
      $past(prd_clearing_equals_output) || alert_o)

  if (SecMasking) begin : gen_sec_cm_key_masking_svas
      // The number of clock cycles a regular AES round takes - only used for assertions.
      localparam int unsigned NumCyclesPerRound = (SecSBoxImpl == SBoxImplDom) ? 5 : 1;
      logic unused_param;
      assign unused_param = (NumCyclesPerRound == 1);
      // Ensure that SubBytes gets fresh PRD input for every evaluation unless mask forcing is
      // enabled. We effectively check that the PRNG has been updated at least once within the
      // last NumCyclesPerRound cycles. This also holds for the very first round, as the PRNG
      // is always updated in the last cycle of the IDLE state and/or the first cycle of the
      // INIT state.
      `ASSERT(AesSecCmKeyMaskingPrdSubBytes,
          sub_bytes_en == SP2V_HIGH && ($past(sub_bytes_en) == SP2V_LOW ||
              ($past(sub_bytes_out_req) == SP2V_HIGH &&
               $past(sub_bytes_out_ack) == SP2V_HIGH)) |=>
          $past(prd_sub_bytes) != $past(prd_sub_bytes, NumCyclesPerRound + 1) ||
          SecAllowForcingMasks && force_masks_i)

      // Ensure that the PRNG has been updated between masking the input and starting the first
      // SubBytes evaluation/KeyExpand operation unless mask forcing is enabled. For AES-256,
      // we just spend 1 cycle in the INIT state and KeyExpand isn't evaluating its S-Boxes,
      // i.e., no fresh randomness is required. For the other key lengths, KeyExpand evaluates
      // its S-Boxes which takes NumCyclesPerRound cycles. When computing the start key for
      // decryption, the input isn't loaded and the PRNG is thus not advanced.
      `ASSERT(AesSecCmKeyMaskingInitialPrngUpdateSubBytes,
          sub_bytes_en == SP2V_HIGH && $past(sub_bytes_en) == SP2V_LOW |=>
          (key_len_i == AES_256 &&
              $past(prd_masking) != $past(prd_masking, 3)) ||
          ((key_len_i == AES_128 || key_len_i == AES_192) &&
              $past(prd_masking) != $past(prd_masking, NumCyclesPerRound + 2)) ||
          (SecAllowForcingMasks && force_masks_i))
      `ASSERT(AesSecCmKeyMaskingInitialPrngUpdateKeyExpand,
          key_expand_en == SP2V_HIGH && $past(key_expand_en) == SP2V_LOW |=>
          (key_len_i == AES_256 &&
              $past(prd_masking) != $past(prd_masking, 3)) ||
          ((key_len_i == AES_128 || key_len_i == AES_192) &&
              $past(prd_masking) != $past(prd_masking, 2)) ||
          (SecAllowForcingMasks && force_masks_i) || dec_key_gen_o == SP2V_HIGH)

      // Ensure none of the state shares keeps being constant during encryption/decryption
      // unless mask forcing is enabled. Even though unlikely it's not impossible that one
      // share remains constant throughout one round. The SVAs thus only fire if a share
      // remains constant across two rounds.
      for (genvar s = 0; s < NumShares; s++) begin : gen_sec_cm_key_masking_share_svas
        `ASSERT(AesSecCmKeyMaskingStateShare, state_we == SP2V_HIGH &&
            (crypt_i == SP2V_HIGH || crypt_o == SP2V_HIGH) |=>
            state_q[s] != $past(state_q[s], NumCyclesPerRound) ||
            $past(state_q[s], NumCyclesPerRound) != $past(state_q[s], 2*NumCyclesPerRound) ||
            (SecAllowForcingMasks && force_masks_i) || dec_key_gen_o == SP2V_HIGH)
        `ASSERT(AesSecCmKeyMaskingOutputShare,
            (out_valid_o == SP2V_HIGH && $past(out_valid_o) == SP2V_LOW) &&
            (crypt_o == SP2V_HIGH) |=>
            $past(state_o[s]) != $past(state_q[s], NumCyclesPerRound) ||
            $past(state_q[s], NumCyclesPerRound) != $past(state_q[s], 2*NumCyclesPerRound) ||
            (SecAllowForcingMasks && force_masks_i) || dec_key_gen_o == SP2V_HIGH)
      end
  end

  // Make sure the output of the masking PRNG is properly extracted without creating overlaps
  // in the data input masks, or between the PRD fed to the key expand module and SubBytes.
  if (WidthPRDSBox > 8) begin : gen_prd_extract_assert
    // For one row of the state matrix, extract the WidthPRDSBox-8 MSBs of the per-S-Box PRD from
    // the PRNG output.
    function automatic logic [3:0][(WidthPRDSBox-8)-1:0] aes_prd_get_msbs(
      logic [(4*WidthPRDSBox)-1:0] in
    );
      logic [3:0][(WidthPRDSBox-8)-1:0] prd_msbs;
      for (int i = 0; i < 4; i++) begin
        prd_msbs[i] = in[(i*WidthPRDSBox) + 8 +: (WidthPRDSBox-8)];
      end
      return prd_msbs;
    endfunction

    // For one row of the state matrix, undo the extraction of LSBs and MSBs of the per-S-Box PRD
    // from the PRNG output. This can be used to verify proper extraction (no overlap of output
    // masks and PRD for masked Canright S-Box implementations, no unused PRNG output).
    function automatic logic [4*WidthPRDSBox-1:0] aes_prd_concat_bits(
      logic [3:0]                 [7:0] prd_lsbs,
      logic [3:0][(WidthPRDSBox-8)-1:0] prd_msbs
    );
      logic [(4*WidthPRDSBox)-1:0] prd;
      for (int i = 0; i < 4; i++) begin
        prd[(i*WidthPRDSBox) +: WidthPRDSBox] = {prd_msbs[i], prd_lsbs[i]};
      end
      return prd;
    endfunction

    // Check for correct extraction of masking PRNG output without overlaps.
    logic            [WidthPRDMasking-1:0] unused_prd_masking;
    logic [3:0][3:0][(WidthPRDSBox-8)-1:0] unused_prd_msbs;
    for (genvar i = 0; i < 4; i++) begin : gen_unused_prd_msbs
      assign unused_prd_msbs[i] = aes_prd_get_msbs(prd_masking[i * WidthPRDRow +: WidthPRDRow]);
    end
    for (genvar i = 0; i < 4; i++) begin : gen_unused_prd_masking
      assign unused_prd_masking[i * WidthPRDRow +: WidthPRDRow] =
          aes_prd_concat_bits(data_in_mask[i], unused_prd_msbs[i]);
    end
    assign unused_prd_masking[WidthPRDMasking-1 -: WidthPRDKey] = prd_key_expand;
    `ASSERT(AesMskgPrdExtraction, prd_masking == unused_prd_masking)
  end
  //VCS coverage on
  // pragma coverage on
`endif

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES cipher core control
//
// This module controls the AES cipher core including the key expand module.

`include "prim_assert.sv"

module aes_cipher_control import aes_pkg::*;
#(
  parameter bit         SecMasking  = 0,
  parameter sbox_impl_e SecSBoxImpl = SBoxImplDom
) (
  input  logic                    clk_i,
  input  logic                    rst_ni,

  // Input handshake signals
  input  sp2v_e                   in_valid_i,
  output sp2v_e                   in_ready_o,

  // Output handshake signals
  output sp2v_e                   out_valid_o,
  input  sp2v_e                   out_ready_i,

  // Control and sync signals
  input  logic                    cfg_valid_i,
  input  ciph_op_e                op_i,
  input  key_len_e                key_len_i,
  input  sp2v_e                   crypt_i,
  output sp2v_e                   crypt_o,
  input  sp2v_e                   dec_key_gen_i,
  output sp2v_e                   dec_key_gen_o,
  input  logic                    prng_reseed_i,
  output logic                    prng_reseed_o,
  input  logic                    key_clear_i,
  output logic                    key_clear_o,
  input  logic                    data_out_clear_i,
  output logic                    data_out_clear_o,
  input  logic                    mux_sel_err_i,
  input  logic                    sp_enc_err_i,
  input  logic                    op_err_i,
  input  logic                    alert_fatal_i,
  output logic                    alert_o,

  // Control signals for masking PRNG
  output logic                    prng_update_o,
  output logic                    prng_reseed_req_o,
  input  logic                    prng_reseed_ack_i,

  // Control and sync signals for cipher data path
  output state_sel_e              state_sel_o,
  output sp2v_e                   state_we_o,
  output sp2v_e                   sub_bytes_en_o,
  input  sp2v_e                   sub_bytes_out_req_i,
  output sp2v_e                   sub_bytes_out_ack_o,
  output add_rk_sel_e             add_rk_sel_o,

  // Control and sync signals for key expand data path
  output ciph_op_e                key_expand_op_o,
  output key_full_sel_e           key_full_sel_o,
  output sp2v_e                   key_full_we_o,
  output key_dec_sel_e            key_dec_sel_o,
  output sp2v_e                   key_dec_we_o,
  output sp2v_e                   key_expand_en_o,
  input  sp2v_e                   key_expand_out_req_i,
  output sp2v_e                   key_expand_out_ack_o,
  output logic                    key_expand_clear_o,
  output logic [3:0]              key_expand_round_o,
  output key_words_sel_e          key_words_sel_o,
  output round_key_sel_e          round_key_sel_o
);

  // Signals
  logic                          [3:0] rnd_ctr;
  sp2v_e                               crypt_d, crypt_q;
  sp2v_e                               dec_key_gen_d, dec_key_gen_q;
  logic                                prng_reseed_d, prng_reseed_q;
  logic                                key_clear_d, key_clear_q;
  logic                                data_out_clear_d, data_out_clear_q;
  sp2v_e                               sub_bytes_out_req;
  sp2v_e                               key_expand_out_req;
  sp2v_e                               in_valid;
  sp2v_e                               out_ready;
  sp2v_e                               crypt;
  sp2v_e                               dec_key_gen;
  logic                                mux_sel_err;
  logic                                mr_err;
  logic                                sp_enc_err;
  logic                                rnd_ctr_err;

  // Sparsified FSM signals. These are needed for connecting the individual bits of the Sp2V
  // signals to the single-rail FSMs.
  logic           [Sp2VWidth-1:0]      sp_in_valid;
  logic           [Sp2VWidth-1:0]      sp_in_ready;
  logic           [Sp2VWidth-1:0]      sp_out_valid;
  logic           [Sp2VWidth-1:0]      sp_out_ready;
  logic           [Sp2VWidth-1:0]      sp_crypt;
  logic           [Sp2VWidth-1:0]      sp_dec_key_gen;
  logic           [Sp2VWidth-1:0]      sp_state_we;
  logic           [Sp2VWidth-1:0]      sp_sub_bytes_en;
  logic           [Sp2VWidth-1:0]      sp_sub_bytes_out_req;
  logic           [Sp2VWidth-1:0]      sp_sub_bytes_out_ack;
  logic           [Sp2VWidth-1:0]      sp_key_full_we;
  logic           [Sp2VWidth-1:0]      sp_key_dec_we;
  logic           [Sp2VWidth-1:0]      sp_key_expand_en;
  logic           [Sp2VWidth-1:0]      sp_key_expand_out_req;
  logic           [Sp2VWidth-1:0]      sp_key_expand_out_ack;
  logic           [Sp2VWidth-1:0]      sp_crypt_d;
  logic           [Sp2VWidth-1:0]      sp_crypt_q;
  logic           [Sp2VWidth-1:0]      sp_dec_key_gen_d;
  logic           [Sp2VWidth-1:0]      sp_dec_key_gen_q;

  // Multi-rail signals. These are outputs of the single-rail FSMs and need combining.
  logic           [Sp2VWidth-1:0]      mr_alert;
  logic           [Sp2VWidth-1:0]      mr_prng_update;
  logic           [Sp2VWidth-1:0]      mr_prng_reseed_req;
  logic           [Sp2VWidth-1:0]      mr_key_expand_clear;
  logic           [Sp2VWidth-1:0]      mr_prng_reseed_d;
  logic           [Sp2VWidth-1:0]      mr_key_clear_d;
  logic           [Sp2VWidth-1:0]      mr_data_out_clear_d;

  state_sel_e     [Sp2VWidth-1:0]      mr_state_sel;
  add_rk_sel_e    [Sp2VWidth-1:0]      mr_add_rk_sel;
  key_full_sel_e  [Sp2VWidth-1:0]      mr_key_full_sel;
  key_dec_sel_e   [Sp2VWidth-1:0]      mr_key_dec_sel;
  key_words_sel_e [Sp2VWidth-1:0]      mr_key_words_sel;
  round_key_sel_e [Sp2VWidth-1:0]      mr_round_key_sel;

  logic           [Sp2VWidth-1:0][3:0] mr_rnd_ctr;

  /////////
  // FSM //
  /////////

  // Convert sp2v_e signals to sparsified inputs.
  assign sp_in_valid           = {in_valid};
  assign sp_out_ready          = {out_ready};
  assign sp_crypt              = {crypt};
  assign sp_dec_key_gen        = {dec_key_gen};
  assign sp_sub_bytes_out_req  = {sub_bytes_out_req};
  assign sp_key_expand_out_req = {key_expand_out_req};
  assign sp_crypt_q            = {crypt_q};
  assign sp_dec_key_gen_q      = {dec_key_gen_q};

  // SEC_CM: CIPHER.FSM.REDUN
  // SEC_CM: CIPHER.CTR.REDUN
  // For every bit in the Sp2V signals, one separate rail is instantiated. The inputs and outputs
  // of every rail are buffered to prevent aggressive synthesis optimizations.
  for (genvar i = 0; i < Sp2VWidth; i++) begin : gen_fsm
    if (SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_fsm_p
      aes_cipher_control_fsm_p #(
        .SecMasking  ( SecMasking  ),
        .SecSBoxImpl ( SecSBoxImpl )
      ) u_aes_cipher_control_fsm_i (
        .clk_i                 ( clk_i                    ),
        .rst_ni                ( rst_ni                   ),

        .in_valid_i            ( sp_in_valid[i]           ), // Sparsified
        .in_ready_o            ( sp_in_ready[i]           ), // Sparsified

        .out_valid_o           ( sp_out_valid[i]          ), // Sparsified
        .out_ready_i           ( sp_out_ready[i]          ), // Sparsified

        .cfg_valid_i           ( cfg_valid_i              ),
        .op_i                  ( op_i                     ),
        .key_len_i             ( key_len_i                ),
        .crypt_i               ( sp_crypt[i]              ), // Sparsified
        .dec_key_gen_i         ( sp_dec_key_gen[i]        ), // Sparsified
        .prng_reseed_i         ( prng_reseed_i            ),
        .key_clear_i           ( key_clear_i              ),
        .data_out_clear_i      ( data_out_clear_i         ),
        .mux_sel_err_i         ( mux_sel_err              ),
        .sp_enc_err_i          ( sp_enc_err               ),
        .rnd_ctr_err_i         ( rnd_ctr_err              ),
        .op_err_i              ( op_err_i                 ),
        .alert_fatal_i         ( alert_fatal_i            ),
        .alert_o               ( mr_alert[i]              ), // OR-combine

        .prng_update_o         ( mr_prng_update[i]        ), // OR-combine
        .prng_reseed_req_o     ( mr_prng_reseed_req[i]    ), // OR-combine
        .prng_reseed_ack_i     ( prng_reseed_ack_i        ),

        .state_sel_o           ( mr_state_sel[i]          ), // OR-combine
        .state_we_o            ( sp_state_we[i]           ), // Sparsified
        .sub_bytes_en_o        ( sp_sub_bytes_en[i]       ), // Sparsified
        .sub_bytes_out_req_i   ( sp_sub_bytes_out_req[i]  ), // Sparsified
        .sub_bytes_out_ack_o   ( sp_sub_bytes_out_ack[i]  ), // Sparsified
        .add_rk_sel_o          ( mr_add_rk_sel[i]         ), // OR-combine

        .key_full_sel_o        ( mr_key_full_sel[i]       ), // OR-combine
        .key_full_we_o         ( sp_key_full_we[i]        ), // Sparsified
        .key_dec_sel_o         ( mr_key_dec_sel[i]        ), // OR-combine
        .key_dec_we_o          ( sp_key_dec_we[i]         ), // Sparsified
        .key_expand_en_o       ( sp_key_expand_en[i]      ), // Sparsified
        .key_expand_out_req_i  ( sp_key_expand_out_req[i] ), // Sparsified
        .key_expand_out_ack_o  ( sp_key_expand_out_ack[i] ), // Sparsified
        .key_expand_clear_o    ( mr_key_expand_clear[i]   ), // OR-combine
        .rnd_ctr_o             ( mr_rnd_ctr[i]            ), // OR-combine
        .key_words_sel_o       ( mr_key_words_sel[i]      ), // OR-combine
        .round_key_sel_o       ( mr_round_key_sel[i]      ), // OR-combine

        .crypt_q_i             ( sp_crypt_q[i]            ), // Sparsified
        .crypt_d_o             ( sp_crypt_d[i]            ), // Sparsified
        .dec_key_gen_q_i       ( sp_dec_key_gen_q[i]      ), // Sparsified
        .dec_key_gen_d_o       ( sp_dec_key_gen_d[i]      ), // Sparsified
        .prng_reseed_q_i       ( prng_reseed_q            ),
        .prng_reseed_d_o       ( mr_prng_reseed_d[i]      ), // AND-combine
        .key_clear_q_i         ( key_clear_q              ),
        .key_clear_d_o         ( mr_key_clear_d[i]        ), // AND-combine
        .data_out_clear_q_i    ( data_out_clear_q         ),
        .data_out_clear_d_o    ( mr_data_out_clear_d[i]   )  // AND-combine
      );
    end else begin : gen_fsm_n
      aes_cipher_control_fsm_n #(
        .SecMasking  ( SecMasking  ),
        .SecSBoxImpl ( SecSBoxImpl )
      ) u_aes_cipher_control_fsm_i (
        .clk_i                 ( clk_i                    ),
        .rst_ni                ( rst_ni                   ),

        .in_valid_ni           ( sp_in_valid[i]           ), // Sparsified
        .in_ready_no           ( sp_in_ready[i]           ), // Sparsified

        .out_valid_no          ( sp_out_valid[i]          ), // Sparsified
        .out_ready_ni          ( sp_out_ready[i]          ), // Sparsified

        .cfg_valid_i           ( cfg_valid_i              ),
        .op_i                  ( op_i                     ),
        .key_len_i             ( key_len_i                ),
        .crypt_ni              ( sp_crypt[i]              ), // Sparsified
        .dec_key_gen_ni        ( sp_dec_key_gen[i]        ), // Sparsified
        .prng_reseed_i         ( prng_reseed_i            ),
        .key_clear_i           ( key_clear_i              ),
        .data_out_clear_i      ( data_out_clear_i         ),
        .mux_sel_err_i         ( mux_sel_err              ),
        .sp_enc_err_i          ( sp_enc_err               ),
        .rnd_ctr_err_i         ( rnd_ctr_err              ),
        .op_err_i              ( op_err_i                 ),
        .alert_fatal_i         ( alert_fatal_i            ),
        .alert_o               ( mr_alert[i]              ), // OR-combine

        .prng_update_o         ( mr_prng_update[i]        ), // OR-combine
        .prng_reseed_req_o     ( mr_prng_reseed_req[i]    ), // OR-combine
        .prng_reseed_ack_i     ( prng_reseed_ack_i        ),

        .state_sel_o           ( mr_state_sel[i]          ), // OR-combine
        .state_we_no           ( sp_state_we[i]           ), // Sparsified
        .sub_bytes_en_no       ( sp_sub_bytes_en[i]       ), // Sparsified
        .sub_bytes_out_req_ni  ( sp_sub_bytes_out_req[i]  ), // Sparsified
        .sub_bytes_out_ack_no  ( sp_sub_bytes_out_ack[i]  ), // Sparsified
        .add_rk_sel_o          ( mr_add_rk_sel[i]         ), // OR-combine

        .key_full_sel_o        ( mr_key_full_sel[i]       ), // OR-combine
        .key_full_we_no        ( sp_key_full_we[i]        ), // Sparsified
        .key_dec_sel_o         ( mr_key_dec_sel[i]        ), // OR-combine
        .key_dec_we_no         ( sp_key_dec_we[i]         ), // Sparsified
        .key_expand_en_no      ( sp_key_expand_en[i]      ), // Sparsified
        .key_expand_out_req_ni ( sp_key_expand_out_req[i] ), // Sparsified
        .key_expand_out_ack_no ( sp_key_expand_out_ack[i] ), // Sparsified
        .key_expand_clear_o    ( mr_key_expand_clear[i]   ), // OR-combine
        .rnd_ctr_o             ( mr_rnd_ctr[i]            ), // OR-combine
        .key_words_sel_o       ( mr_key_words_sel[i]      ), // OR-combine
        .round_key_sel_o       ( mr_round_key_sel[i]      ), // OR-combine

        .crypt_q_ni            ( sp_crypt_q[i]            ), // Sparsified
        .crypt_d_no            ( sp_crypt_d[i]            ), // Sparsified
        .dec_key_gen_q_ni      ( sp_dec_key_gen_q[i]      ), // Sparsified
        .dec_key_gen_d_no      ( sp_dec_key_gen_d[i]      ), // Sparsified
        .prng_reseed_q_i       ( prng_reseed_q            ),
        .prng_reseed_d_o       ( mr_prng_reseed_d[i]      ), // AND-combine
        .key_clear_q_i         ( key_clear_q              ),
        .key_clear_d_o         ( mr_key_clear_d[i]        ), // AND-combine
        .data_out_clear_q_i    ( data_out_clear_q         ),
        .data_out_clear_d_o    ( mr_data_out_clear_d[i]   )  // AND-combine
      );
    end
  end

  // Convert sparsified outputs to sp2v_e type.
  assign in_ready_o           = sp2v_e'(sp_in_ready);
  assign out_valid_o          = sp2v_e'(sp_out_valid);
  assign state_we_o           = sp2v_e'(sp_state_we);
  assign sub_bytes_en_o       = sp2v_e'(sp_sub_bytes_en);
  assign sub_bytes_out_ack_o  = sp2v_e'(sp_sub_bytes_out_ack);
  assign key_full_we_o        = sp2v_e'(sp_key_full_we);
  assign key_dec_we_o         = sp2v_e'(sp_key_dec_we);
  assign key_expand_en_o      = sp2v_e'(sp_key_expand_en);
  assign key_expand_out_ack_o = sp2v_e'(sp_key_expand_out_ack);
  assign crypt_d              = sp2v_e'(sp_crypt_d);
  assign dec_key_gen_d        = sp2v_e'(sp_dec_key_gen_d);

  // Combine single-bit FSM outputs.
  // OR: One bit is sufficient to drive the corresponding output bit high.
  assign alert_o            = |mr_alert;
  assign prng_update_o      = |mr_prng_update;
  assign prng_reseed_req_o  = |mr_prng_reseed_req;
  assign key_expand_clear_o = |mr_key_expand_clear;
  // AND: Only if all bits are high, the corresponding status is signaled which will lead to
  // the clearing of these trigger bits.
  assign prng_reseed_d      = &mr_prng_reseed_d;
  assign key_clear_d        = &mr_key_clear_d;
  assign data_out_clear_d   = &mr_data_out_clear_d;

  // Combine multi-bit, sparse FSM outputs. We simply OR them together. If the FSMs don't provide
  // the same outputs, two cases are possible:
  // - An invalid encoding results: A downstream checker will fire, see mux_sel_err_i.
  // - A valid encoding results: The outputs are compared below to cover this case, see mr_err;
  always_comb begin : combine_sparse_signals
    state_sel_o     = state_sel_e'({StateSelWidth{1'b0}});
    add_rk_sel_o    = add_rk_sel_e'({AddRKSelWidth{1'b0}});
    key_full_sel_o  = key_full_sel_e'({KeyFullSelWidth{1'b0}});
    key_dec_sel_o   = key_dec_sel_e'({KeyDecSelWidth{1'b0}});
    key_words_sel_o = key_words_sel_e'({KeyWordsSelWidth{1'b0}});
    round_key_sel_o = round_key_sel_e'({RoundKeySelWidth{1'b0}});
    mr_err          = 1'b0;

    for (int i = 0; i < Sp2VWidth; i++) begin
      state_sel_o     = state_sel_e'({state_sel_o}         | {mr_state_sel[i]});
      add_rk_sel_o    = add_rk_sel_e'({add_rk_sel_o}       | {mr_add_rk_sel[i]});
      key_full_sel_o  = key_full_sel_e'({key_full_sel_o}   | {mr_key_full_sel[i]});
      key_dec_sel_o   = key_dec_sel_e'({key_dec_sel_o}     | {mr_key_dec_sel[i]});
      key_words_sel_o = key_words_sel_e'({key_words_sel_o} | {mr_key_words_sel[i]});
      round_key_sel_o = round_key_sel_e'({round_key_sel_o} | {mr_round_key_sel[i]});
    end

    for (int i = 0; i < Sp2VWidth; i++) begin
      if (state_sel_o     != mr_state_sel[i]     ||
          add_rk_sel_o    != mr_add_rk_sel[i]    ||
          key_full_sel_o  != mr_key_full_sel[i]  ||
          key_dec_sel_o   != mr_key_dec_sel[i]   ||
          key_words_sel_o != mr_key_words_sel[i] ||
          round_key_sel_o != mr_round_key_sel[i]) begin
        mr_err = 1'b1;
      end
    end
  end

  // Collect errors in mux selector signals.
  assign mux_sel_err = mux_sel_err_i | mr_err;

  // Combine counter signals. We simply OR them together. If the FSMs don't provide the same
  // outputs, rnd_ctr_err will be set.
  always_comb begin : combine_counter_signals
    rnd_ctr     = '0;
    rnd_ctr_err = 1'b0;
    for (int i = 0; i < Sp2VWidth; i++) begin
      rnd_ctr |= mr_rnd_ctr[i];
    end

    for (int i = 0; i < Sp2VWidth; i++) begin
      if (rnd_ctr != mr_rnd_ctr[i]) begin
        rnd_ctr_err = 1'b1;
      end
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_fsm
    if (!rst_ni) begin
      prng_reseed_q      <= 1'b0;
      key_clear_q        <= 1'b0;
      data_out_clear_q   <= 1'b0;
    end else begin
      prng_reseed_q      <= prng_reseed_d;
      key_clear_q        <= key_clear_d;
      data_out_clear_q   <= data_out_clear_d;
    end
  end

  // Use separate signal for key expand operation, forward round.
  assign key_expand_op_o    = (dec_key_gen_d == SP2V_HIGH ||
                               dec_key_gen_q == SP2V_HIGH) ? CIPH_FWD : op_i;
  assign key_expand_round_o = rnd_ctr;

  // Let the main controller know whate we are doing.
  assign crypt_o          = crypt_q;
  assign dec_key_gen_o    = dec_key_gen_q;
  assign prng_reseed_o    = prng_reseed_q;
  assign key_clear_o      = key_clear_q;
  assign data_out_clear_o = data_out_clear_q;


  //////////////////////////////
  // Sparsely Encoded Signals //
  //////////////////////////////

  // SEC_CM: CTRL.SPARSE
  // We use sparse encodings for various critical signals and must ensure that:
  // 1. The synthesis tool doesn't optimize away the sparse encoding.
  // 2. The sparsely encoded signal is always valid. More precisely, an alert or SVA is triggered
  //    if a sparse signal takes on an invalid value.
  // 3. The alert signal remains asserted until reset even if the sparse signal becomes valid again
  //    This is achieved by driving the control FSM into the terminal error state whenever any
  //    sparsely encoded signal becomes invalid.
  //
  // If any sparsely encoded signal becomes invalid, the cipher core further immediately de-asserts
  // the out_valid_o signal to prevent any data from being released.

  // The following primitives are used to place a size-only constraint on the
  // flops in order to prevent optimizations on these status signals.
  logic [Sp2VWidth-1:0] crypt_q_raw;
  prim_flop #(
    .Width      ( Sp2VWidth            ),
    .ResetValue ( Sp2VWidth'(SP2V_LOW) )
  ) u_crypt_regs (
    .clk_i  ( clk_i       ),
    .rst_ni ( rst_ni      ),
    .d_i    ( crypt_d     ),
    .q_o    ( crypt_q_raw )
  );

  logic [Sp2VWidth-1:0] dec_key_gen_q_raw;
  prim_flop #(
    .Width      ( Sp2VWidth            ),
    .ResetValue ( Sp2VWidth'(SP2V_LOW) )
  ) u_dec_key_gen_regs (
    .clk_i  ( clk_i             ),
    .rst_ni ( rst_ni            ),
    .d_i    ( dec_key_gen_d     ),
    .q_o    ( dec_key_gen_q_raw )
  );

  // We use vectors of sparsely encoded signals to reduce code duplication.
  localparam int unsigned NumSp2VSig = 8;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig;
  sp2v_e [NumSp2VSig-1:0]                sp2v_sig_chk;
  logic  [NumSp2VSig-1:0][Sp2VWidth-1:0] sp2v_sig_chk_raw;
  logic  [NumSp2VSig-1:0]                sp2v_sig_err;

  assign sp2v_sig[0] = in_valid_i;
  assign sp2v_sig[1] = out_ready_i;
  assign sp2v_sig[2] = crypt_i;
  assign sp2v_sig[3] = dec_key_gen_i;
  assign sp2v_sig[4] = sp2v_e'(crypt_q_raw);
  assign sp2v_sig[5] = sp2v_e'(dec_key_gen_q_raw);
  assign sp2v_sig[6] = sub_bytes_out_req_i;
  assign sp2v_sig[7] = key_expand_out_req_i;

  // All signals inside sp2v_sig except for sub_bytes/key_expand_out_req_i are driven and consumed
  // by multi-rail FSMs.
  localparam bit [NumSp2VSig-1:0] Sp2VEnSecBuf = 8'b1100_0000;

  // Individually check sparsely encoded signals.
  for (genvar i = 0; i < NumSp2VSig; i++) begin : gen_sel_buf_chk
    aes_sel_buf_chk #(
      .Num      ( Sp2VNum         ),
      .Width    ( Sp2VWidth       ),
      .EnSecBuf ( Sp2VEnSecBuf[i] )
    ) u_aes_sp2v_sig_buf_chk_i (
      .clk_i  ( clk_i               ),
      .rst_ni ( rst_ni              ),
      .sel_i  ( sp2v_sig[i]         ),
      .sel_o  ( sp2v_sig_chk_raw[i] ),
      .err_o  ( sp2v_sig_err[i]     )
    );
    assign sp2v_sig_chk[i] = sp2v_e'(sp2v_sig_chk_raw[i]);
  end

  assign in_valid           = sp2v_sig_chk[0];
  assign out_ready          = sp2v_sig_chk[1];
  assign crypt              = sp2v_sig_chk[2];
  assign dec_key_gen        = sp2v_sig_chk[3];
  assign crypt_q            = sp2v_sig_chk[4];
  assign dec_key_gen_q      = sp2v_sig_chk[5];
  assign sub_bytes_out_req  = sp2v_sig_chk[6];
  assign key_expand_out_req = sp2v_sig_chk[7];

  // Collect encoding errors.
  // We instantiate the checker modules as close as possible to where the sparsely encoded signals
  // are used. Here, we collect also encoding errors detected in other places of the cipher core.
  assign sp_enc_err = |sp2v_sig_err | sp_enc_err_i;

  ////////////////
  // Assertions //
  ////////////////

  // Selectors must be known/valid
  `ASSERT(AesCiphOpValid, cfg_valid_i |-> op_i inside {
      CIPH_FWD,
      CIPH_INV
      })

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES cipher core control FSM
//
// This module contains the AES cipher core control FSM.

`include "prim_assert.sv"

module aes_cipher_control_fsm import aes_pkg::*;
#(
  parameter bit         SecMasking  = 0,
  parameter sbox_impl_e SecSBoxImpl = SBoxImplDom
) (
  input  logic             clk_i,
  input  logic             rst_ni,

  // Input handshake signals
  input  logic             in_valid_i,           // Sparsify using multi-rail.
  output logic             in_ready_o,           // Sparsify using multi-rail.

  // Output handshake signals
  output logic             out_valid_o,          // Sparsify using multi-rail.
  input  logic             out_ready_i,          // Sparsify using multi-rail.

  // Control and sync signals
  input  logic             cfg_valid_i,          // Used for SVAs only.
  input  ciph_op_e         op_i,
  input  key_len_e         key_len_i,
  input  logic             crypt_i,              // Sparsify using multi-rail.
  input  logic             dec_key_gen_i,        // Sparsify using multi-rail.
  input  logic             prng_reseed_i,
  input  logic             key_clear_i,
  input  logic             data_out_clear_i,
  input  logic             mux_sel_err_i,
  input  logic             sp_enc_err_i,
  input  logic             rnd_ctr_err_i,
  input  logic             op_err_i,
  input  logic             alert_fatal_i,
  output logic             alert_o,

  // Control signals for masking PRNG
  output logic             prng_update_o,
  output logic             prng_reseed_req_o,
  input  logic             prng_reseed_ack_i,

  // Control and sync signals for cipher data path
  output state_sel_e       state_sel_o,
  output logic             state_we_o,           // Sparsify using multi-rail.
  output logic             sub_bytes_en_o,       // Sparsify using multi-rail.
  input  logic             sub_bytes_out_req_i,  // Sparsify using multi-rail.
  output logic             sub_bytes_out_ack_o,  // Sparsify using multi-rail.
  output add_rk_sel_e      add_rk_sel_o,

  // Control and sync signals for key expand data path
  output key_full_sel_e    key_full_sel_o,
  output logic             key_full_we_o,        // Sparsify using multi-rail.
  output key_dec_sel_e     key_dec_sel_o,
  output logic             key_dec_we_o,         // Sparsify using multi-rail.
  output logic             key_expand_en_o,      // Sparsify using multi-rail.
  input  logic             key_expand_out_req_i, // Sparsify using multi-rail.
  output logic             key_expand_out_ack_o, // Sparsify using multi-rail.
  output logic             key_expand_clear_o,
  output logic [3:0]       rnd_ctr_o,
  output key_words_sel_e   key_words_sel_o,
  output round_key_sel_e   round_key_sel_o,

  // Register signals
  input  logic             crypt_q_i,            // Sparsify using multi-rail.
  output logic             crypt_d_o,            // Sparsify using multi-rail.
  input  logic             dec_key_gen_q_i,      // Sparsify using multi-rail.
  output logic             dec_key_gen_d_o,      // Sparsify using multi-rail.
  input  logic             prng_reseed_q_i,
  output logic             prng_reseed_d_o,
  input  logic             key_clear_q_i,
  output logic             key_clear_d_o,
  input  logic             data_out_clear_q_i,
  output logic             data_out_clear_d_o
);

  // cfg_valid_i is used for SVAs only.
  logic unused_cfg_valid;
  assign unused_cfg_valid = cfg_valid_i;

  // Tie off unused inputs.
  if (!SecMasking) begin : gen_unused_prng_reseed
    logic unused_prng_reseed;
    assign unused_prng_reseed = prng_reseed_i;
  end

  // Signals
  aes_cipher_ctrl_e aes_cipher_ctrl_ns, aes_cipher_ctrl_cs;
  logic             advance;
  logic       [2:0] cyc_ctr_d, cyc_ctr_q;
  logic             cyc_ctr_expr;
  logic             prng_reseed_done_d, prng_reseed_done_q;
  logic       [3:0] rnd_ctr_d, rnd_ctr_q;
  logic       [3:0] num_rounds_d, num_rounds_q;
  logic       [3:0] num_rounds_regular;

  // Use separate signal for number of regular rounds.
  assign num_rounds_regular = num_rounds_q - 4'd1;

  // FSM
  always_comb begin : aes_cipher_ctrl_fsm

    // Handshake signals
    in_ready_o           = 1'b0;
    out_valid_o          = 1'b0;

    // Masking PRNG signals
    prng_update_o        = 1'b0;
    prng_reseed_req_o    = 1'b0;

    // Cipher data path
    state_sel_o          = STATE_ROUND;
    state_we_o           = 1'b0;
    add_rk_sel_o         = ADD_RK_ROUND;
    sub_bytes_en_o       = 1'b0;
    sub_bytes_out_ack_o  = 1'b0;

    // Key expand data path
    key_full_sel_o       = KEY_FULL_ROUND;
    key_full_we_o        = 1'b0;
    key_dec_sel_o        = KEY_DEC_EXPAND;
    key_dec_we_o         = 1'b0;
    key_expand_en_o      = 1'b0;
    key_expand_out_ack_o = 1'b0;
    key_expand_clear_o   = 1'b0;
    key_words_sel_o      = KEY_WORDS_ZERO;
    round_key_sel_o      = ROUND_KEY_DIRECT;

    // FSM
    aes_cipher_ctrl_ns   = aes_cipher_ctrl_cs;
    num_rounds_d         = num_rounds_q;
    rnd_ctr_d            = rnd_ctr_q;
    crypt_d_o            = crypt_q_i;
    dec_key_gen_d_o      = dec_key_gen_q_i;
    prng_reseed_d_o      = prng_reseed_q_i;
    key_clear_d_o        = key_clear_q_i;
    data_out_clear_d_o   = data_out_clear_q_i;
    prng_reseed_done_d   = prng_reseed_done_q | prng_reseed_ack_i;
    advance              = 1'b0;
    cyc_ctr_d            = (SecSBoxImpl == SBoxImplDom) ? cyc_ctr_q + 3'd1 : 3'd0;

    // Alert
    alert_o              = 1'b0;

    unique case (aes_cipher_ctrl_cs)

      CIPHER_CTRL_IDLE: begin
        cyc_ctr_d = 3'd0;

        // Signal that we are ready, wait for handshake.
        in_ready_o = 1'b1;
        if (in_valid_i) begin
          if (SecMasking && prng_reseed_i && !dec_key_gen_i && !crypt_i) begin
            // Reseed the masking PRNG without starting encryption/decryption or generation of the
            // start key for decryption.
            prng_reseed_d_o    = 1'b1;
            prng_reseed_done_d = 1'b0;
            aes_cipher_ctrl_ns = CIPHER_CTRL_PRNG_RESEED;

          end else if (key_clear_i || data_out_clear_i) begin
            // Clear internal key registers. The cipher core muxes are used to clear the data
            // output registers.
            key_clear_d_o      = key_clear_i;
            data_out_clear_d_o = data_out_clear_i;

            // To clear the data output registers, we must first clear the state.
            aes_cipher_ctrl_ns = data_out_clear_i ? CIPHER_CTRL_CLEAR_S : CIPHER_CTRL_CLEAR_KD;

          end else if (dec_key_gen_i || crypt_i) begin
            // Start encryption/decryption or generation of start key for decryption.
            crypt_d_o       = ~dec_key_gen_i & crypt_i;
            dec_key_gen_d_o =  dec_key_gen_i;

            // Latch whether we shall reseed the masking PRNG.
            prng_reseed_d_o = SecMasking & prng_reseed_i;

            // Load input data to state
            state_sel_o = dec_key_gen_i ? STATE_CLEAR : STATE_INIT;
            state_we_o  = 1'b1;

            // Make the masking PRNG advance. The current pseudo-random data is used to mask the
            // input data.
            prng_update_o = SecMasking;

            // Init key expand
            key_expand_clear_o = 1'b1;

            // Load full key
            key_full_sel_o = dec_key_gen_i ? KEY_FULL_ENC_INIT :
                        (op_i == CIPH_FWD) ? KEY_FULL_ENC_INIT :
                        (op_i == CIPH_INV) ? KEY_FULL_DEC_INIT :
                                             KEY_FULL_ENC_INIT;
            key_full_we_o  = 1'b1;

            // Load num_rounds, initialize round counter.
            num_rounds_d = (key_len_i == AES_128) ? 4'd10 :
                           (key_len_i == AES_192) ? 4'd12 :
                                                    4'd14;
            rnd_ctr_d          = '0;
            aes_cipher_ctrl_ns = CIPHER_CTRL_INIT;

          end else begin
            // Handshake without a valid command. We should never get here. If we do (e.g. via a
            // malicious glitch), error out immediately.
            aes_cipher_ctrl_ns = CIPHER_CTRL_ERROR;
          end
        end
      end

      CIPHER_CTRL_INIT: begin
        // Initial round: just add key to state
        add_rk_sel_o = ADD_RK_INIT;

        // Select key words for initial add_round_key
        key_words_sel_o = (dec_key_gen_q_i)            ? KEY_WORDS_ZERO :
            (key_len_i == AES_128)                     ? KEY_WORDS_0123 :
            (key_len_i == AES_192 && op_i == CIPH_FWD) ? KEY_WORDS_0123 :
            (key_len_i == AES_192 && op_i == CIPH_INV) ? KEY_WORDS_2345 :
            (key_len_i == AES_256 && op_i == CIPH_FWD) ? KEY_WORDS_0123 :
            (key_len_i == AES_256 && op_i == CIPH_INV) ? KEY_WORDS_4567 : KEY_WORDS_ZERO;

        // Clear masking PRNG reseed status.
        prng_reseed_done_d = 1'b0;

        // AES-256 has two round keys available right from beginning. Pseudo-random data is
        // required by KeyExpand only.
        if (key_len_i != AES_256) begin
          // Advance in sync with KeyExpand. Based on the S-Box implementation, it can take
          // multiple cycles to finish. Wait for handshake. The DOM S-Boxes consume fresh PRD
          // only in the first clock cycle. By requesting the PRNG update in any clock cycle
          // other than the last one, the PRD fed into the DOM S-Boxes is guaranteed to be stable.
          // This is better in terms of SCA resistance. Request the PRNG update in the first cycle.
          advance         = key_expand_out_req_i & cyc_ctr_expr;
          prng_update_o   = (SecSBoxImpl == SBoxImplDom) ? cyc_ctr_q == 3'd0 : SecMasking;
          key_expand_en_o = 1'b1;
          if (advance) begin
            key_expand_out_ack_o = 1'b1;
            state_we_o           = ~dec_key_gen_q_i;
            key_full_we_o        = 1'b1;
            rnd_ctr_d            = rnd_ctr_q + 4'b0001;
            cyc_ctr_d            = 3'd0;
            aes_cipher_ctrl_ns   = CIPHER_CTRL_ROUND;
          end
        end else begin
          prng_update_o      = SecMasking;
          state_we_o         = ~dec_key_gen_q_i;
          rnd_ctr_d          = rnd_ctr_q + 4'b0001;
          cyc_ctr_d          = 3'd0;
          aes_cipher_ctrl_ns = CIPHER_CTRL_ROUND;
        end
      end

      CIPHER_CTRL_ROUND: begin
        // Normal rounds

        // Select key words for add_round_key
        key_words_sel_o = (dec_key_gen_q_i)            ? KEY_WORDS_ZERO :
            (key_len_i == AES_128)                     ? KEY_WORDS_0123 :
            (key_len_i == AES_192 && op_i == CIPH_FWD) ? KEY_WORDS_2345 :
            (key_len_i == AES_192 && op_i == CIPH_INV) ? KEY_WORDS_0123 :
            (key_len_i == AES_256 && op_i == CIPH_FWD) ? KEY_WORDS_4567 :
            (key_len_i == AES_256 && op_i == CIPH_INV) ? KEY_WORDS_0123 : KEY_WORDS_ZERO;

        // Keep requesting PRNG reseeding until it is acknowledged.
        prng_reseed_req_o = SecMasking & prng_reseed_q_i & ~prng_reseed_done_q;

        // Select round key: direct or mixed (equivalent inverse cipher)
        round_key_sel_o = (op_i == CIPH_FWD) ? ROUND_KEY_DIRECT :
                          (op_i == CIPH_INV) ? ROUND_KEY_MIXED  : ROUND_KEY_DIRECT;

        // Advance in sync with SubBytes and KeyExpand. Based on the S-Box implementation, both can
        // take multiple cycles to finish. Wait for handshake. The DOM S-Boxes consume fresh PRD
        // only in the first clock cycle. By requesting the PRNG update in any clock cycle other
        // than the last one, the PRD fed into the DOM S-Boxes is guaranteed to be stable. This is
        // better in terms of SCA resistance. Request the PRNG update in the first cycle. Non-DOM
        // S-Boxes need fresh PRD in every clock cycle.
        advance = key_expand_out_req_i & cyc_ctr_expr & (dec_key_gen_q_i | sub_bytes_out_req_i);
        prng_update_o   = (SecSBoxImpl == SBoxImplDom) ? cyc_ctr_q == 3'd0 : SecMasking;
        sub_bytes_en_o  = ~dec_key_gen_q_i;
        key_expand_en_o = 1'b1;

        if (advance) begin
          sub_bytes_out_ack_o  = ~dec_key_gen_q_i;
          key_expand_out_ack_o = 1'b1;

          state_we_o    = ~dec_key_gen_q_i;
          key_full_we_o = 1'b1;

          // Update round
          rnd_ctr_d     = rnd_ctr_q + 4'b0001;
          cyc_ctr_d     = 3'd0;

          // Are we doing the last regular round?
          if (rnd_ctr_q >= num_rounds_regular) begin
            aes_cipher_ctrl_ns = CIPHER_CTRL_FINISH;

            if (dec_key_gen_q_i) begin
              // Write decryption key.
              key_dec_we_o = 1'b1;

              // Indicate that we are done, try to perform the handshake. But we don't wait here.
              // If we don't get the handshake now, we will wait in the finish state. When using
              // masking, we only finish if the masking PRNG has been reseeded.
              out_valid_o = SecMasking ? (prng_reseed_q_i ? prng_reseed_done_q : 1'b1) : 1'b1;
              if (out_valid_o && out_ready_i) begin
                // Go to idle state directly.
                dec_key_gen_d_o    = 1'b0;
                prng_reseed_d_o    = 1'b0;
                aes_cipher_ctrl_ns = CIPHER_CTRL_IDLE;
              end
            end
          end // rnd_ctr_q
        end // SubBytes/KeyExpand REQ/ACK
      end

      CIPHER_CTRL_FINISH: begin
        // Final round

        // Select key words for add_round_key
        key_words_sel_o = (dec_key_gen_q_i)            ? KEY_WORDS_ZERO :
            (key_len_i == AES_128)                     ? KEY_WORDS_0123 :
            (key_len_i == AES_192 && op_i == CIPH_FWD) ? KEY_WORDS_2345 :
            (key_len_i == AES_192 && op_i == CIPH_INV) ? KEY_WORDS_0123 :
            (key_len_i == AES_256 && op_i == CIPH_FWD) ? KEY_WORDS_4567 :
            (key_len_i == AES_256 && op_i == CIPH_INV) ? KEY_WORDS_0123 : KEY_WORDS_ZERO;

        // Skip mix_columns
        add_rk_sel_o = ADD_RK_FINAL;

        // Keep requesting PRNG reseeding until it is acknowledged.
        prng_reseed_req_o = SecMasking & prng_reseed_q_i & ~prng_reseed_done_q;

        // SEC_CM: DATA_REG.KEY.SCA
        // Once we're done, we won't need the state anymore. We actually clear it when progressing
        // to the next state.
        state_sel_o = STATE_CLEAR;

        // SEC_CM: DATA_REG.LOCAL_ESC
        // Advance in sync with SubBytes. Based on the S-Box implementation, it can take multiple
        // cycles to finish. Only indicate that we are done if:
        // - we have valid output (SubBytes finished),
        // - the masking PRNG has been reseeded (if masking is used),
        // - all mux selector signals are valid (don't release data in case of errors), and
        // - all sparsely encoded signals are valid (don't release data in case of errors).
        // Perform both handshakes simultaneously.
        advance        = (sub_bytes_out_req_i & cyc_ctr_expr) | dec_key_gen_q_i;
        sub_bytes_en_o = ~dec_key_gen_q_i;
        out_valid_o    = (mux_sel_err_i || sp_enc_err_i || op_err_i) ? 1'b0         :
            SecMasking ? (prng_reseed_q_i ? prng_reseed_done_q & advance : advance) : advance;

        // Stop updating the cycle counter once we have valid output.
        cyc_ctr_d =
            (SecSBoxImpl == SBoxImplDom) ? (!advance ? cyc_ctr_q + 3'd1 : cyc_ctr_q) : 3'd0;

        // The DOM S-Boxes consume fresh PRD only in the first clock cycle. By requesting the PRNG
        // update in any clock cycle other than the last one, the PRD fed into the DOM S-Boxes is
        // guaranteed to be stable. This is better in terms of SCA resistance. Request the PRNG
        // update in the first cycle. We update it only once and in the last cycle for non-DOM
        // S-Boxes where otherwise updating the PRNG while being stalled would cause the S-Boxes
        // to be re-evaluated, thereby creating additional SCA leakage.
        prng_update_o =
            (SecSBoxImpl == SBoxImplDom) ? cyc_ctr_q == 3'd0 : out_valid_o & out_ready_i;

        if (out_valid_o && out_ready_i) begin
          sub_bytes_out_ack_o = ~dec_key_gen_q_i;

          // Clear the state.
          state_we_o          = 1'b1;
          crypt_d_o           = 1'b0;
          cyc_ctr_d           = 3'd0;
          // If we were generating the decryption key and didn't get the handshake in the last
          // regular round, we should clear dec_key_gen now.
          dec_key_gen_d_o     = 1'b0;
          prng_reseed_d_o     = 1'b0;
          aes_cipher_ctrl_ns  = CIPHER_CTRL_IDLE;
        end
      end

      CIPHER_CTRL_PRNG_RESEED: begin
        // Keep requesting PRNG reseeding until it is acknowledged.
        prng_reseed_req_o = prng_reseed_q_i & ~prng_reseed_done_q;

        // Once we're done, wait for handshake.
        out_valid_o = prng_reseed_done_q;
        if (out_valid_o && out_ready_i) begin
          prng_reseed_d_o    = 1'b0;
          aes_cipher_ctrl_ns = CIPHER_CTRL_IDLE;
        end
      end

      CIPHER_CTRL_CLEAR_S: begin
        // Clear the state with pseudo-random data.
        state_we_o         = 1'b1;
        state_sel_o        = STATE_CLEAR;
        aes_cipher_ctrl_ns = CIPHER_CTRL_CLEAR_KD;
      end

      CIPHER_CTRL_CLEAR_KD: begin
        // Clear internal key registers and/or external data output registers.
        if (key_clear_q_i) begin
          key_full_sel_o = KEY_FULL_CLEAR;
          key_full_we_o  = 1'b1;
          key_dec_sel_o  = KEY_DEC_CLEAR;
          key_dec_we_o   = 1'b1;
        end
        if (data_out_clear_q_i) begin
          // Forward the state (previously cleared with psuedo-random data).
          // SEC_CM: DATA_REG.SEC_WIPE
          add_rk_sel_o    = ADD_RK_INIT;
          key_words_sel_o = KEY_WORDS_ZERO;
          round_key_sel_o = ROUND_KEY_DIRECT;
        end
        // Indicate that we are done, wait for handshake.
        out_valid_o = 1'b1;
        if (out_ready_i) begin
          key_clear_d_o      = 1'b0;
          data_out_clear_d_o = 1'b0;
          aes_cipher_ctrl_ns = CIPHER_CTRL_IDLE;
        end
      end

      CIPHER_CTRL_ERROR: begin
        // SEC_CM: CIPHER.FSM.LOCAL_ESC
        // Terminal error state
        alert_o = 1'b1;
      end

      // We should never get here. If we do (e.g. via a malicious glitch), error out immediately.
      default: begin
        aes_cipher_ctrl_ns = CIPHER_CTRL_ERROR;
        alert_o = 1'b1;
      end
    endcase

    // Unconditionally jump into the terminal error state in case a mux selector or a sparsely
    // encoded signal becomes invalid, in case we have detected a fault in the round counter,
    // or if a fatal alert has been triggered.
    if (mux_sel_err_i || sp_enc_err_i || rnd_ctr_err_i || op_err_i || alert_fatal_i) begin
      aes_cipher_ctrl_ns = CIPHER_CTRL_ERROR;
    end
  end

  // SEC_CM: CIPHER.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, aes_cipher_ctrl_ns,
      aes_cipher_ctrl_cs, aes_cipher_ctrl_e, CIPHER_CTRL_IDLE)

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_fsm
    if (!rst_ni) begin
      prng_reseed_done_q <= 1'b0;
      rnd_ctr_q          <= '0;
      num_rounds_q       <= '0;
    end else begin
      prng_reseed_done_q <= prng_reseed_done_d;
      rnd_ctr_q          <= rnd_ctr_d;
      num_rounds_q       <= num_rounds_d;
    end
  end

  assign rnd_ctr_o = rnd_ctr_q;

  if (SecSBoxImpl == SBoxImplDom) begin : gen_cyc_ctr
    always_ff @(posedge clk_i or negedge rst_ni) begin : reg_cyc_ctr
      if (!rst_ni) begin
        cyc_ctr_q <= 3'd0;
      end else begin
        cyc_ctr_q <= cyc_ctr_d;
      end
    end
    assign cyc_ctr_expr = cyc_ctr_q >= 3'd4;
  end else begin : gen_no_cyc_ctr
    logic [2:0] unused_cyc_ctr;
    assign cyc_ctr_q      = cyc_ctr_d;
    assign unused_cyc_ctr = cyc_ctr_q;
    assign cyc_ctr_expr   = 1'b1;
  end

  ////////////////
  // Assertions //
  ////////////////

  // Create a lint error to reduce the risk of accidentally disabling the masking.
  `ASSERT_STATIC_LINT_ERROR(AesCipherControlFsmSecMaskingNonDefault, SecMasking == 1)

  // Create a lint error to reduce the risk of accidentally using a less secure SBox
  // implementation.
  `ASSERT_STATIC_LINT_ERROR(AesCipherControlFsmSecSBoxImplNonDefault, SecSBoxImpl == SBoxImplDom)

  // Selectors must be known/valid
  `ASSERT(AesCiphOpValid, cfg_valid_i |-> op_i inside {
      CIPH_FWD,
      CIPH_INV
      })
  `ASSERT(AesKeyLenValid, cfg_valid_i |-> key_len_i inside {
      AES_128,
      AES_192,
      AES_256
      })
  `ASSERT(AesCipherControlStateValid, !alert_o |-> aes_cipher_ctrl_cs inside {
      CIPHER_CTRL_IDLE,
      CIPHER_CTRL_INIT,
      CIPHER_CTRL_ROUND,
      CIPHER_CTRL_FINISH,
      CIPHER_CTRL_PRNG_RESEED,
      CIPHER_CTRL_CLEAR_S,
      CIPHER_CTRL_CLEAR_KD
      })

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES cipher core control FSM
//
// This module contains the AES cipher core control FSM operating on
// and producing the positive values of important control signals.

module aes_cipher_control_fsm_p import aes_pkg::*;
#(
  parameter bit         SecMasking  = 0,
  parameter sbox_impl_e SecSBoxImpl = SBoxImplDom
) (
  input  logic             clk_i,
  input  logic             rst_ni,

  // Input handshake signals
  input  logic             in_valid_i,            // Sparsify using multi-rail.
  output logic             in_ready_o,            // Sparsify using multi-rail.

  // Output handshake signals
  output logic             out_valid_o,           // Sparsify using multi-rail.
  input  logic             out_ready_i,           // Sparsify using multi-rail.

  // Control and sync signals
  input  logic             cfg_valid_i,           // Used for SVAs only.
  input  ciph_op_e         op_i,
  input  key_len_e         key_len_i,
  input  logic             crypt_i,               // Sparsify using multi-rail.
  input  logic             dec_key_gen_i,         // Sparsify using multi-rail.
  input  logic             prng_reseed_i,
  input  logic             key_clear_i,
  input  logic             data_out_clear_i,
  input  logic             mux_sel_err_i,
  input  logic             sp_enc_err_i,
  input  logic             rnd_ctr_err_i,
  input  logic             op_err_i,
  input  logic             alert_fatal_i,
  output logic             alert_o,

  // Control signals for masking PRNG
  output logic             prng_update_o,
  output logic             prng_reseed_req_o,
  input  logic             prng_reseed_ack_i,

  // Control and sync signals for cipher data path
  output state_sel_e       state_sel_o,
  output logic             state_we_o,            // Sparsify using multi-rail.
  output logic             sub_bytes_en_o,        // Sparsify using multi-rail.
  input  logic             sub_bytes_out_req_i,   // Sparsify using multi-rail.
  output logic             sub_bytes_out_ack_o,   // Sparsify using multi-rail.
  output add_rk_sel_e      add_rk_sel_o,

  // Control and sync signals for key expand data path
  output key_full_sel_e    key_full_sel_o,
  output logic             key_full_we_o,         // Sparsify using multi-rail.
  output key_dec_sel_e     key_dec_sel_o,
  output logic             key_dec_we_o,          // Sparsify using multi-rail.
  output logic             key_expand_en_o,       // Sparsify using multi-rail.
  input  logic             key_expand_out_req_i,  // Sparsify using multi-rail.
  output logic             key_expand_out_ack_o,  // Sparsify using multi-rail.
  output logic             key_expand_clear_o,
  output logic [3:0]       rnd_ctr_o,
  output key_words_sel_e   key_words_sel_o,
  output round_key_sel_e   round_key_sel_o,

  // Register signals
  input  logic             crypt_q_i,             // Sparsify using multi-rail.
  output logic             crypt_d_o,             // Sparsify using multi-rail.
  input  logic             dec_key_gen_q_i,       // Sparsify using multi-rail.
  output logic             dec_key_gen_d_o,       // Sparsify using multi-rail.
  input  logic             prng_reseed_q_i,
  output logic             prng_reseed_d_o,
  input  logic             key_clear_q_i,
  output logic             key_clear_d_o,
  input  logic             data_out_clear_q_i,
  output logic             data_out_clear_d_o
);

  /////////////////////
  // Input Buffering //
  /////////////////////

  localparam int NumInBufBits = $bits({
    in_valid_i,
    out_ready_i,
    cfg_valid_i,
    op_i,
    key_len_i,
    crypt_i,
    dec_key_gen_i,
    prng_reseed_i,
    key_clear_i,
    data_out_clear_i,
    mux_sel_err_i,
    sp_enc_err_i,
    rnd_ctr_err_i,
    op_err_i,
    alert_fatal_i,
    prng_reseed_ack_i,
    sub_bytes_out_req_i,
    key_expand_out_req_i,
    crypt_q_i,
    dec_key_gen_q_i,
    prng_reseed_q_i,
    key_clear_q_i,
    data_out_clear_q_i
  });

  logic [NumInBufBits-1:0] in, in_buf;

  assign in = {
    in_valid_i,
    out_ready_i,
    cfg_valid_i,
    op_i,
    key_len_i,
    crypt_i,
    dec_key_gen_i,
    prng_reseed_i,
    key_clear_i,
    data_out_clear_i,
    mux_sel_err_i,
    sp_enc_err_i,
    rnd_ctr_err_i,
    op_err_i,
    alert_fatal_i,
    prng_reseed_ack_i,
    sub_bytes_out_req_i,
    key_expand_out_req_i,
    crypt_q_i,
    dec_key_gen_q_i,
    prng_reseed_q_i,
    key_clear_q_i,
    data_out_clear_q_i
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumInBufBits)
  ) u_prim_buf_in (
    .in_i(in),
    .out_o(in_buf)
  );

  logic                 in_valid;
  logic                 out_ready;
  logic                 cfg_valid;
  ciph_op_e             op;
  logic [$bits(op)-1:0] op_raw;
  key_len_e             key_len;
  logic                 crypt;
  logic                 dec_key_gen;
  logic                 prng_reseed;
  logic                 key_clear;
  logic                 data_out_clear;
  logic                 mux_sel_err;
  logic                 sp_enc_err;
  logic                 rnd_ctr_err;
  logic                 op_err;
  logic                 alert_fatal;
  logic                 prng_reseed_ack;
  logic                 sub_bytes_out_req;
  logic                 key_expand_out_req;
  logic                 crypt_q;
  logic                 dec_key_gen_q;
  logic                 prng_reseed_q;
  logic                 key_clear_q;
  logic                 data_out_clear_q;

  assign {in_valid,
          out_ready,
          cfg_valid,
          op_raw,
          key_len,
          crypt,
          dec_key_gen,
          prng_reseed,
          key_clear,
          data_out_clear,
          mux_sel_err,
          sp_enc_err,
          rnd_ctr_err,
          op_err,
          alert_fatal,
          prng_reseed_ack,
          sub_bytes_out_req,
          key_expand_out_req,
          crypt_q,
          dec_key_gen_q,
          prng_reseed_q,
          key_clear_q,
          data_out_clear_q} = in_buf;

  assign op = ciph_op_e'(op_raw);

  // Intermediate output signals
  logic             in_ready;
  logic             out_valid;
  logic             alert;
  logic             prng_update;
  logic             prng_reseed_req;
  state_sel_e       state_sel;
  logic             state_we;
  logic             sub_bytes_en;
  logic             sub_bytes_out_ack;
  add_rk_sel_e      add_rk_sel;
  key_full_sel_e    key_full_sel;
  logic             key_full_we;
  key_dec_sel_e     key_dec_sel;
  logic             key_dec_we;
  logic             key_expand_en;
  logic             key_expand_out_ack;
  logic             key_expand_clear;
  logic [3:0]       rnd_ctr;
  key_words_sel_e   key_words_sel;
  round_key_sel_e   round_key_sel;
  logic             crypt_d;
  logic             dec_key_gen_d;
  logic             prng_reseed_d;
  logic             key_clear_d;
  logic             data_out_clear_d;

  /////////////////
  // Regular FSM //
  /////////////////

  aes_cipher_control_fsm #(
    .SecMasking  ( SecMasking  ),
    .SecSBoxImpl ( SecSBoxImpl )
  ) u_aes_cipher_control_fsm (
    .clk_i                 ( clk_i                  ),
    .rst_ni                ( rst_ni                 ),

    .in_valid_i            ( in_valid               ),
    .in_ready_o            ( in_ready               ),

    .out_valid_o           ( out_valid              ),
    .out_ready_i           ( out_ready              ),

    .cfg_valid_i           ( cfg_valid              ),
    .op_i                  ( op                     ),
    .key_len_i             ( key_len                ),
    .crypt_i               ( crypt                  ),
    .dec_key_gen_i         ( dec_key_gen            ),
    .prng_reseed_i         ( prng_reseed            ),
    .key_clear_i           ( key_clear              ),
    .data_out_clear_i      ( data_out_clear         ),
    .mux_sel_err_i         ( mux_sel_err            ),
    .sp_enc_err_i          ( sp_enc_err             ),
    .rnd_ctr_err_i         ( rnd_ctr_err            ),
    .op_err_i              ( op_err                 ),
    .alert_fatal_i         ( alert_fatal            ),
    .alert_o               ( alert                  ),

    .prng_update_o         ( prng_update            ),
    .prng_reseed_req_o     ( prng_reseed_req        ),
    .prng_reseed_ack_i     ( prng_reseed_ack        ),

    .state_sel_o           ( state_sel              ),
    .state_we_o            ( state_we               ),
    .sub_bytes_en_o        ( sub_bytes_en           ),
    .sub_bytes_out_req_i   ( sub_bytes_out_req      ),
    .sub_bytes_out_ack_o   ( sub_bytes_out_ack      ),
    .add_rk_sel_o          ( add_rk_sel             ),

    .key_full_sel_o        ( key_full_sel           ),
    .key_full_we_o         ( key_full_we            ),
    .key_dec_sel_o         ( key_dec_sel            ),
    .key_dec_we_o          ( key_dec_we             ),
    .key_expand_en_o       ( key_expand_en          ),
    .key_expand_out_req_i  ( key_expand_out_req     ),
    .key_expand_out_ack_o  ( key_expand_out_ack     ),
    .key_expand_clear_o    ( key_expand_clear       ),
    .rnd_ctr_o             ( rnd_ctr                ),
    .key_words_sel_o       ( key_words_sel          ),
    .round_key_sel_o       ( round_key_sel          ),

    .crypt_q_i             ( crypt_q                ),
    .crypt_d_o             ( crypt_d                ),
    .dec_key_gen_q_i       ( dec_key_gen_q          ),
    .dec_key_gen_d_o       ( dec_key_gen_d          ),
    .key_clear_q_i         ( key_clear_q            ),
    .key_clear_d_o         ( key_clear_d            ),
    .prng_reseed_q_i       ( prng_reseed_q          ),
    .prng_reseed_d_o       ( prng_reseed_d          ),
    .data_out_clear_q_i    ( data_out_clear_q       ),
    .data_out_clear_d_o    ( data_out_clear_d       )
  );

  //////////////////////
  // Output Buffering //
  //////////////////////

  localparam int NumOutBufBits = $bits({
    in_ready_o,
    out_valid_o,
    alert_o,
    prng_update_o,
    prng_reseed_req_o,
    state_sel_o,
    state_we_o,
    sub_bytes_en_o,
    sub_bytes_out_ack_o,
    add_rk_sel_o,
    key_full_sel_o,
    key_full_we_o,
    key_dec_sel_o,
    key_dec_we_o,
    key_expand_en_o,
    key_expand_out_ack_o,
    key_expand_clear_o,
    rnd_ctr_o,
    key_words_sel_o,
    round_key_sel_o,
    crypt_d_o,
    dec_key_gen_d_o,
    key_clear_d_o,
    prng_reseed_d_o,
    data_out_clear_d_o
  });

  logic [NumOutBufBits-1:0] out, out_buf;

  assign out = {
    in_ready,
    out_valid,
    alert,
    prng_update,
    prng_reseed_req,
    state_sel,
    state_we,
    sub_bytes_en,
    sub_bytes_out_ack,
    add_rk_sel,
    key_full_sel,
    key_full_we,
    key_dec_sel,
    key_dec_we,
    key_expand_en,
    key_expand_out_ack,
    key_expand_clear,
    rnd_ctr,
    key_words_sel,
    round_key_sel,
    crypt_d,
    dec_key_gen_d,
    key_clear_d,
    prng_reseed_d,
    data_out_clear_d
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumOutBufBits)
  ) u_prim_buf_out (
    .in_i(out),
    .out_o(out_buf)
  );

  assign {in_ready_o,
          out_valid_o,
          alert_o,
          prng_update_o,
          prng_reseed_req_o,
          state_sel_o,
          state_we_o,
          sub_bytes_en_o,
          sub_bytes_out_ack_o,
          add_rk_sel_o,
          key_full_sel_o,
          key_full_we_o,
          key_dec_sel_o,
          key_dec_we_o,
          key_expand_en_o,
          key_expand_out_ack_o,
          key_expand_clear_o,
          rnd_ctr_o,
          key_words_sel_o,
          round_key_sel_o,
          crypt_d_o,
          dec_key_gen_d_o,
          key_clear_d_o,
          prng_reseed_d_o,
          data_out_clear_d_o} = out_buf;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES cipher core control FSM
//
// This module contains the AES cipher core control FSM operating on and producing the negated
// values of important control signals. This is achieved by:
// - instantiating the regular AES cipher core control FSM operating on and producing the positive
//   values of these signals, and
// - inverting these signals between the regular FSM and the prim_buf synthesis barriers.
// Synthesis tools will then push the inverters into the actual FSM.

module aes_cipher_control_fsm_n import aes_pkg::*;
#(
  parameter bit         SecMasking  = 0,
  parameter sbox_impl_e SecSBoxImpl = SBoxImplDom
) (
  input  logic             clk_i,
  input  logic             rst_ni,

  // Input handshake signals
  input  logic             in_valid_ni,           // Sparsify using multi-rail.
  output logic             in_ready_no,           // Sparsify using multi-rail.

  // Output handshake signals
  output logic             out_valid_no,          // Sparsify using multi-rail.
  input  logic             out_ready_ni,          // Sparsify using multi-rail.

  // Control and sync signals
  input  logic             cfg_valid_i,           // Used for SVAs only.
  input  ciph_op_e         op_i,
  input  key_len_e         key_len_i,
  input  logic             crypt_ni,              // Sparsify using multi-rail.
  input  logic             dec_key_gen_ni,        // Sparsify using multi-rail.
  input  logic             prng_reseed_i,
  input  logic             key_clear_i,
  input  logic             data_out_clear_i,
  input  logic             mux_sel_err_i,
  input  logic             sp_enc_err_i,
  input  logic             rnd_ctr_err_i,
  input  logic             op_err_i,
  input  logic             alert_fatal_i,
  output logic             alert_o,

  // Control signals for masking PRNG
  output logic             prng_update_o,
  output logic             prng_reseed_req_o,
  input  logic             prng_reseed_ack_i,

  // Control and sync signals for cipher data path
  output state_sel_e       state_sel_o,
  output logic             state_we_no,           // Sparsify using multi-rail.
  output logic             sub_bytes_en_no,       // Sparsify using multi-rail.
  input  logic             sub_bytes_out_req_ni,  // Sparsify using multi-rail.
  output logic             sub_bytes_out_ack_no,  // Sparsify using multi-rail.
  output add_rk_sel_e      add_rk_sel_o,

  // Control and sync signals for key expand data path
  output key_full_sel_e    key_full_sel_o,
  output logic             key_full_we_no,        // Sparsify using multi-rail.
  output key_dec_sel_e     key_dec_sel_o,
  output logic             key_dec_we_no,         // Sparsify using multi-rail.
  output logic             key_expand_en_no,      // Sparsify using multi-rail.
  input  logic             key_expand_out_req_ni, // Sparsify using multi-rail.
  output logic             key_expand_out_ack_no, // Sparsify using multi-rail.
  output logic             key_expand_clear_o,
  output logic [3:0]       rnd_ctr_o,
  output key_words_sel_e   key_words_sel_o,
  output round_key_sel_e   round_key_sel_o,

  // Register signals
  input  logic             crypt_q_ni,            // Sparsify using multi-rail.
  output logic             crypt_d_no,            // Sparsify using multi-rail.
  input  logic             dec_key_gen_q_ni,      // Sparsify using multi-rail.
  output logic             dec_key_gen_d_no,      // Sparsify using multi-rail.
  input  logic             prng_reseed_q_i,
  output logic             prng_reseed_d_o,
  input  logic             key_clear_q_i,
  output logic             key_clear_d_o,
  input  logic             data_out_clear_q_i,
  output logic             data_out_clear_d_o
);

  /////////////////////
  // Input Buffering //
  /////////////////////

  localparam int NumInBufBits = $bits({
    in_valid_ni,
    out_ready_ni,
    cfg_valid_i,
    op_i,
    key_len_i,
    crypt_ni,
    dec_key_gen_ni,
    prng_reseed_i,
    key_clear_i,
    data_out_clear_i,
    mux_sel_err_i,
    sp_enc_err_i,
    rnd_ctr_err_i,
    op_err_i,
    alert_fatal_i,
    prng_reseed_ack_i,
    sub_bytes_out_req_ni,
    key_expand_out_req_ni,
    crypt_q_ni,
    dec_key_gen_q_ni,
    prng_reseed_q_i,
    key_clear_q_i,
    data_out_clear_q_i
  });

  logic [NumInBufBits-1:0] in, in_buf;

  assign in = {
    in_valid_ni,
    out_ready_ni,
    cfg_valid_i,
    op_i,
    key_len_i,
    crypt_ni,
    dec_key_gen_ni,
    prng_reseed_i,
    key_clear_i,
    data_out_clear_i,
    mux_sel_err_i,
    sp_enc_err_i,
    rnd_ctr_err_i,
    op_err_i,
    alert_fatal_i,
    prng_reseed_ack_i,
    sub_bytes_out_req_ni,
    key_expand_out_req_ni,
    crypt_q_ni,
    dec_key_gen_q_ni,
    prng_reseed_q_i,
    key_clear_q_i,
    data_out_clear_q_i
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumInBufBits)
  ) u_prim_buf_in (
    .in_i(in),
    .out_o(in_buf)
  );

  logic                 in_valid_n;
  logic                 out_ready_n;
  logic                 cfg_valid;
  ciph_op_e             op;
  logic [$bits(op)-1:0] op_raw;
  key_len_e             key_len;
  logic                 crypt_n;
  logic                 dec_key_gen_n;
  logic                 prng_reseed;
  logic                 key_clear;
  logic                 data_out_clear;
  logic                 mux_sel_err;
  logic                 sp_enc_err;
  logic                 rnd_ctr_err;
  logic                 op_err;
  logic                 alert_fatal;
  logic                 prng_reseed_ack;
  logic                 sub_bytes_out_req_n;
  logic                 key_expand_out_req_n;
  logic                 crypt_q_n;
  logic                 dec_key_gen_q_n;
  logic                 prng_reseed_q;
  logic                 key_clear_q;
  logic                 data_out_clear_q;

  assign {in_valid_n,
          out_ready_n,
          cfg_valid,
          op_raw,
          key_len,
          crypt_n,
          dec_key_gen_n,
          prng_reseed,
          key_clear,
          data_out_clear,
          mux_sel_err,
          sp_enc_err,
          rnd_ctr_err,
          op_err,
          alert_fatal,
          prng_reseed_ack,
          sub_bytes_out_req_n,
          key_expand_out_req_n,
          crypt_q_n,
          dec_key_gen_q_n,
          prng_reseed_q,
          key_clear_q,
          data_out_clear_q} = in_buf;

  assign op = ciph_op_e'(op_raw);

  // Intermediate output signals
  logic             in_ready;
  logic             out_valid;
  logic             alert;
  logic             prng_update;
  logic             prng_reseed_req;
  state_sel_e       state_sel;
  logic             state_we;
  logic             sub_bytes_en;
  logic             sub_bytes_out_ack;
  add_rk_sel_e      add_rk_sel;
  key_full_sel_e    key_full_sel;
  logic             key_full_we;
  key_dec_sel_e     key_dec_sel;
  logic             key_dec_we;
  logic             key_expand_en;
  logic             key_expand_out_ack;
  logic             key_expand_clear;
  key_words_sel_e   key_words_sel;
  round_key_sel_e   round_key_sel;
  logic [3:0]       rnd_ctr;
  logic             crypt_d;
  logic             dec_key_gen_d;
  logic             prng_reseed_d;
  logic             key_clear_d;
  logic             data_out_clear_d;

  /////////////////
  // Regular FSM //
  /////////////////

  // The regular FSM operates on and produces the positive values of important control signals.
  // Invert *_n input signals here to get the positive values for the regular FSM. To obtain the
  // negated outputs, important output signals are inverted further below. Thanks to the prim_buf
  // synthesis optimization barriers, tools will push the inverters into the regular FSM.
  aes_cipher_control_fsm #(
    .SecMasking  ( SecMasking  ),
    .SecSBoxImpl ( SecSBoxImpl )
  ) u_aes_cipher_control_fsm (
    .clk_i                 ( clk_i                 ),
    .rst_ni                ( rst_ni                ),

    .in_valid_i            ( ~in_valid_n           ), // Invert for regular FSM.
    .in_ready_o            ( in_ready              ), // Invert below for negated output.

    .out_valid_o           ( out_valid             ), // Invert below for negated output.
    .out_ready_i           ( ~out_ready_n          ), // Invert for regular FSM.

    .cfg_valid_i           ( cfg_valid             ),
    .op_i                  ( op                    ),
    .key_len_i             ( key_len               ),
    .crypt_i               ( ~crypt_n              ), // Invert for regular FSM.
    .dec_key_gen_i         ( ~dec_key_gen_n        ), // Invert for regular FSM.
    .prng_reseed_i         ( prng_reseed           ),
    .key_clear_i           ( key_clear             ),
    .data_out_clear_i      ( data_out_clear        ),
    .mux_sel_err_i         ( mux_sel_err           ),
    .sp_enc_err_i          ( sp_enc_err            ),
    .rnd_ctr_err_i         ( rnd_ctr_err           ),
    .op_err_i              ( op_err                ),
    .alert_fatal_i         ( alert_fatal           ),
    .alert_o               ( alert                 ),

    .prng_update_o         ( prng_update           ),
    .prng_reseed_req_o     ( prng_reseed_req       ),
    .prng_reseed_ack_i     ( prng_reseed_ack       ),

    .state_sel_o           ( state_sel             ),
    .state_we_o            ( state_we              ), // Invert below for negated output.
    .sub_bytes_en_o        ( sub_bytes_en          ), // Invert below for negated output.
    .sub_bytes_out_req_i   ( ~sub_bytes_out_req_n  ), // Invert for regular FSM.
    .sub_bytes_out_ack_o   ( sub_bytes_out_ack     ), // Invert below for negated output.
    .add_rk_sel_o          ( add_rk_sel            ),

    .key_full_sel_o        ( key_full_sel          ),
    .key_full_we_o         ( key_full_we           ), // Invert below for negated output.
    .key_dec_sel_o         ( key_dec_sel           ),
    .key_dec_we_o          ( key_dec_we            ), // Invert below for negated output.
    .key_expand_en_o       ( key_expand_en         ), // Invert below for negated output.
    .key_expand_out_req_i  ( ~key_expand_out_req_n ), // Invert for regular FSM.
    .key_expand_out_ack_o  ( key_expand_out_ack    ), // Invert below for negated output.
    .key_expand_clear_o    ( key_expand_clear      ),
    .rnd_ctr_o             ( rnd_ctr               ),
    .key_words_sel_o       ( key_words_sel         ),
    .round_key_sel_o       ( round_key_sel         ),

    .crypt_q_i             ( ~crypt_q_n            ), // Invert for regular FSM.
    .crypt_d_o             ( crypt_d               ), // Invert below for negated output.
    .dec_key_gen_q_i       ( ~dec_key_gen_q_n      ), // Invert for regular FSM.
    .dec_key_gen_d_o       ( dec_key_gen_d         ), // Invert below for negated output.
    .key_clear_q_i         ( key_clear_q           ),
    .key_clear_d_o         ( key_clear_d           ),
    .prng_reseed_q_i       ( prng_reseed_q         ),
    .prng_reseed_d_o       ( prng_reseed_d         ),
    .data_out_clear_q_i    ( data_out_clear_q      ),
    .data_out_clear_d_o    ( data_out_clear_d      )
  );

  //////////////////////
  // Output Buffering //
  //////////////////////

  localparam int NumOutBufBits = $bits({
    in_ready_no,
    out_valid_no,
    alert_o,
    prng_update_o,
    prng_reseed_req_o,
    state_sel_o,
    state_we_no,
    sub_bytes_en_no,
    sub_bytes_out_ack_no,
    add_rk_sel_o,
    key_full_sel_o,
    key_full_we_no,
    key_dec_sel_o,
    key_dec_we_no,
    key_expand_en_no,
    key_expand_out_ack_no,
    key_expand_clear_o,
    rnd_ctr_o,
    key_words_sel_o,
    round_key_sel_o,
    crypt_d_no,
    dec_key_gen_d_no,
    key_clear_d_o,
    prng_reseed_d_o,
    data_out_clear_d_o
  });

  logic [NumOutBufBits-1:0] out, out_buf;

  // Important output control signals need to be inverted here. Synthesis tools will push the
  // inverters back into the regular FSM.
  assign out = {
    ~in_ready,
    ~out_valid,
    alert,
    prng_update,
    prng_reseed_req,
    state_sel,
    ~state_we,
    ~sub_bytes_en,
    ~sub_bytes_out_ack,
    add_rk_sel,
    key_full_sel,
    ~key_full_we,
    key_dec_sel,
    ~key_dec_we,
    ~key_expand_en,
    ~key_expand_out_ack,
    key_expand_clear,
    rnd_ctr,
    key_words_sel,
    round_key_sel,
    ~crypt_d,
    ~dec_key_gen_d,
    key_clear_d,
    prng_reseed_d,
    data_out_clear_d
  };

  // This primitive is used to place a size-only constraint on the
  // buffers to act as a synthesis optimization barrier.
  prim_buf #(
    .Width(NumOutBufBits)
  ) u_prim_buf_out (
    .in_i(out),
    .out_o(out_buf)
  );

  assign {in_ready_no,
          out_valid_no,
          alert_o,
          prng_update_o,
          prng_reseed_req_o,
          state_sel_o,
          state_we_no,
          sub_bytes_en_no,
          sub_bytes_out_ack_no,
          add_rk_sel_o,
          key_full_sel_o,
          key_full_we_no,
          key_dec_sel_o,
          key_dec_we_no,
          key_expand_en_no,
          key_expand_out_ack_no,
          key_expand_clear_o,
          rnd_ctr_o,
          key_words_sel_o,
          round_key_sel_o,
          crypt_d_no,
          dec_key_gen_d_no,
          key_clear_d_o,
          prng_reseed_d_o,
          data_out_clear_d_o} = out_buf;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES SubBytes

module aes_sub_bytes import aes_pkg::*;
#(
  parameter sbox_impl_e SecSBoxImpl = SBoxImplDom
) (
  input  logic                              clk_i,
  input  logic                              rst_ni,
  input  sp2v_e                             en_i,
  input  logic                              prd_we_i,
  output sp2v_e                             out_req_o,
  input  sp2v_e                             out_ack_i,
  input  ciph_op_e                          op_i,
  input  logic              [3:0][3:0][7:0] data_i,
  input  logic              [3:0][3:0][7:0] mask_i,
  input  logic [3:0][3:0][WidthPRDSBox-1:0] prd_i,
  output logic              [3:0][3:0][7:0] data_o,
  output logic              [3:0][3:0][7:0] mask_o,
  output logic                              err_o
);

  sp2v_e           en;
  logic            en_err;
  logic [3:0][3:0] out_req;
  sp2v_e           out_ack;
  logic            out_ack_err;

  // Every DOM S-Box instance consumes 28 bits of randomness but itself produces 20 bits for use in
  // another S-Box instance. For other S-Box implementations, only the bits corresponding to prd_i
  // are used. Other bits are ignored and tied to 0.
  logic [3:0][3:0][WidthPRDSBox+19:0] in_prd;
  logic [3:0][3:0]             [19:0] out_prd;

  // SEC_CM: CTRL.SPARSE
  // Check sparsely encoded signals.
  logic [Sp2VWidth-1:0] en_raw;
  aes_sel_buf_chk #(
    .Num      ( Sp2VNum   ),
    .Width    ( Sp2VWidth ),
    .EnSecBuf ( 1'b1      )
  ) u_aes_sb_en_buf_chk (
    .clk_i  ( clk_i  ),
    .rst_ni ( rst_ni ),
    .sel_i  ( en_i   ),
    .sel_o  ( en_raw ),
    .err_o  ( en_err )
  );
  assign en = sp2v_e'(en_raw);

  logic [Sp2VWidth-1:0] out_ack_raw;
  aes_sel_buf_chk #(
    .Num      ( Sp2VNum   ),
    .Width    ( Sp2VWidth ),
    .EnSecBuf ( 1'b1      )
  ) u_aes_sb_out_ack_buf_chk (
    .clk_i  ( clk_i       ),
    .rst_ni ( rst_ni      ),
    .sel_i  ( out_ack_i   ),
    .sel_o  ( out_ack_raw ),
    .err_o  ( out_ack_err )
  );
  assign out_ack = sp2v_e'(out_ack_raw);

  // Individually substitute bytes.
  for (genvar j = 0; j < 4; j++) begin : gen_sbox_j
    for (genvar i = 0; i < 4; i++) begin : gen_sbox_i

      // Rotate the randomness produced by the S-Boxes over the columns but not across rows as
      // MixColumns will operate across rows. The LSBs are taken from the masking PRNG (prd_i)
      // whereas the MSBs are produced by the other S-Box instances.
      assign in_prd[i][j] = {out_prd[i][aes_rot_int(j,4)], prd_i[i][j]};

      aes_sbox #(
        .SecSBoxImpl ( SecSBoxImpl )
      ) u_aes_sbox_ij (
        .clk_i     ( clk_i                ),
        .rst_ni    ( rst_ni               ),
        .en_i      ( en == SP2V_HIGH      ),
        .prd_we_i  ( prd_we_i             ),
        .out_req_o ( out_req[i][j]        ),
        .out_ack_i ( out_ack == SP2V_HIGH ),
        .op_i      ( op_i                 ),
        .data_i    ( data_i[i][j]         ),
        .mask_i    ( mask_i[i][j]         ),
        .prd_i     ( in_prd[i][j]         ),
        .data_o    ( data_o[i][j]         ),
        .mask_o    ( mask_o[i][j]         ),
        .prd_o     ( out_prd[i][j]        )
      );
    end
  end

  // Collect REQ signals.
  assign out_req_o = &out_req ? SP2V_HIGH : SP2V_LOW;

  // Collect encoding errors.
  assign err_o = en_err | out_ack_err;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES SBox

`include "prim_assert.sv"

module aes_sbox import aes_pkg::*;
#(
  parameter sbox_impl_e SecSBoxImpl = SBoxImplLut
) (
  input  logic                     clk_i,
  input  logic                     rst_ni,
  input  logic                     en_i,
  input  logic                     prd_we_i,
  output logic                     out_req_o,
  input  logic                     out_ack_i,
  input  ciph_op_e                 op_i,
  input  logic               [7:0] data_i,
  input  logic               [7:0] mask_i,
  input  logic [WidthPRDSBox+19:0] prd_i,
  output logic               [7:0] data_o,
  output logic               [7:0] mask_o,
  output logic              [19:0] prd_o
);

  // Create a lint error to reduce the risk of accidentally using a less secure SBox
  // implementation.
  `ASSERT_STATIC_LINT_ERROR(AesSBoxSecSBoxImplNonDefault, SecSBoxImpl == SBoxImplDom)

  localparam bit SBoxMasked = (SecSBoxImpl == SBoxImplCanrightMasked ||
                               SecSBoxImpl == SBoxImplCanrightMaskedNoreuse ||
                               SecSBoxImpl == SBoxImplDom) ? 1'b1 : 1'b0;

  localparam bit SBoxSingleCycle = (SecSBoxImpl == SBoxImplDom) ? 1'b0 : 1'b1;

  if (!SBoxMasked) begin : gen_sbox_unmasked
    // Tie off unused inputs.
    logic                     unused_clk;
    logic                     unused_rst;
    logic               [7:0] unused_mask;
    logic [WidthPRDSBox+19:0] unused_prd;
    assign unused_clk  = clk_i;
    assign unused_rst  = rst_ni;
    assign unused_mask = mask_i;
    assign unused_prd  = prd_i;

    if (SecSBoxImpl == SBoxImplCanright) begin : gen_sbox_canright
      aes_sbox_canright u_aes_sbox (
        .op_i   ( op_i   ),
        .data_i ( data_i ),
        .data_o ( data_o )
      );

    end else begin : gen_sbox_lut // SecSBoxImpl == SBoxImplLut
      aes_sbox_lut u_aes_sbox (
        .op_i   ( op_i   ),
        .data_i ( data_i ),
        .data_o ( data_o )
      );
    end

    assign mask_o = '0;
    assign prd_o  = '0;

  end else begin : gen_sbox_masked

    // SEC_CM: KEY.MASKING
    if (SecSBoxImpl == SBoxImplDom) begin : gen_sbox_dom

      aes_sbox_dom u_aes_sbox (
        .clk_i      ( clk_i       ),
        .rst_ni     ( rst_ni      ),
        .en_i       ( en_i        ),
        .prd_we_i   ( prd_we_i    ),
        .out_req_o  ( out_req_o   ),
        .out_ack_i  ( out_ack_i   ),
        .op_i       ( op_i        ),
        .data_i     ( data_i      ),
        .mask_i     ( mask_i      ),
        .prd_i      ( prd_i[27:0] ),
        .data_o     ( data_o      ),
        .mask_o     ( mask_o      ),
        .prd_o      ( prd_o       )
      );

      `ASSERT_INIT(AesWidthPRDSBox, WidthPRDSBox == 8)

    end else if (SecSBoxImpl == SBoxImplCanrightMaskedNoreuse) begin :
        gen_sbox_canright_masked_noreuse
      // Tie off unused inputs.
      logic        unused_clk;
      logic        unused_rst;
      logic [19:0] unused_prd;
      assign unused_clk = clk_i;
      assign unused_rst = rst_ni;
      assign unused_prd = prd_i[WidthPRDSBox+19:WidthPRDSBox];

      aes_sbox_canright_masked_noreuse u_aes_sbox (
        .op_i   ( op_i        ),
        .data_i ( data_i      ),
        .mask_i ( mask_i      ),
        .prd_i  ( prd_i[17:0] ),
        .data_o ( data_o      ),
        .mask_o ( mask_o      )
      );

      assign prd_o = '0;

      `ASSERT_INIT(AesWidthPRDSBox, WidthPRDSBox == 18)

    end else begin : gen_sbox_canright_masked // SecSBoxImpl == SBoxImplCanrightMasked
      // Tie off unused inputs.
      logic        unused_clk;
      logic        unused_rst;
      logic [19:0] unused_prd;
      assign unused_clk = clk_i;
      assign unused_rst = rst_ni;
      assign unused_prd = prd_i[WidthPRDSBox+19:WidthPRDSBox];

      aes_sbox_canright_masked u_aes_sbox (
        .op_i   ( op_i       ),
        .data_i ( data_i     ),
        .mask_i ( mask_i     ),
        .prd_i  ( prd_i[7:0] ),
        .data_o ( data_o     ),
        .mask_o ( mask_o     )
      );

      assign prd_o = '0;

      `ASSERT_INIT(AesWidthPRDSBox, WidthPRDSBox == 8)
    end
  end

  if (SBoxSingleCycle) begin : gen_req_singlecycle
    // Tie off unused inputs.
    logic unused_out_ack;
    logic unused_prd_we;
    assign unused_out_ack = out_ack_i;
    assign unused_prd_we  = prd_we_i;

    // Signal that we have valid output right away.
    assign out_req_o = en_i;
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES LUT-based SBox

module aes_sbox_lut (
  input  aes_pkg::ciph_op_e op_i,
  input  logic [7:0]        data_i,
  output logic [7:0]        data_o
);

  import aes_pkg::*;

  // Define the LUTs
  localparam logic [7:0] SBOX_FWD [256] = '{
    8'h63, 8'h7C, 8'h77, 8'h7B, 8'hF2, 8'h6B, 8'h6F, 8'hC5,
    8'h30, 8'h01, 8'h67, 8'h2B, 8'hFE, 8'hD7, 8'hAB, 8'h76,

    8'hCA, 8'h82, 8'hC9, 8'h7D, 8'hFA, 8'h59, 8'h47, 8'hF0,
    8'hAD, 8'hD4, 8'hA2, 8'hAF, 8'h9C, 8'hA4, 8'h72, 8'hC0,

    8'hB7, 8'hFD, 8'h93, 8'h26, 8'h36, 8'h3F, 8'hF7, 8'hCC,
    8'h34, 8'hA5, 8'hE5, 8'hF1, 8'h71, 8'hD8, 8'h31, 8'h15,

    8'h04, 8'hC7, 8'h23, 8'hC3, 8'h18, 8'h96, 8'h05, 8'h9A,
    8'h07, 8'h12, 8'h80, 8'hE2, 8'hEB, 8'h27, 8'hB2, 8'h75,

    8'h09, 8'h83, 8'h2C, 8'h1A, 8'h1B, 8'h6E, 8'h5A, 8'hA0,
    8'h52, 8'h3B, 8'hD6, 8'hB3, 8'h29, 8'hE3, 8'h2F, 8'h84,

    8'h53, 8'hD1, 8'h00, 8'hED, 8'h20, 8'hFC, 8'hB1, 8'h5B,
    8'h6A, 8'hCB, 8'hBE, 8'h39, 8'h4A, 8'h4C, 8'h58, 8'hCF,

    8'hD0, 8'hEF, 8'hAA, 8'hFB, 8'h43, 8'h4D, 8'h33, 8'h85,
    8'h45, 8'hF9, 8'h02, 8'h7F, 8'h50, 8'h3C, 8'h9F, 8'hA8,

    8'h51, 8'hA3, 8'h40, 8'h8F, 8'h92, 8'h9D, 8'h38, 8'hF5,
    8'hBC, 8'hB6, 8'hDA, 8'h21, 8'h10, 8'hFF, 8'hF3, 8'hD2,

    8'hCD, 8'h0C, 8'h13, 8'hEC, 8'h5F, 8'h97, 8'h44, 8'h17,
    8'hC4, 8'hA7, 8'h7E, 8'h3D, 8'h64, 8'h5D, 8'h19, 8'h73,

    8'h60, 8'h81, 8'h4F, 8'hDC, 8'h22, 8'h2A, 8'h90, 8'h88,
    8'h46, 8'hEE, 8'hB8, 8'h14, 8'hDE, 8'h5E, 8'h0B, 8'hDB,

    8'hE0, 8'h32, 8'h3A, 8'h0A, 8'h49, 8'h06, 8'h24, 8'h5C,
    8'hC2, 8'hD3, 8'hAC, 8'h62, 8'h91, 8'h95, 8'hE4, 8'h79,

    8'hE7, 8'hC8, 8'h37, 8'h6D, 8'h8D, 8'hD5, 8'h4E, 8'hA9,
    8'h6C, 8'h56, 8'hF4, 8'hEA, 8'h65, 8'h7A, 8'hAE, 8'h08,

    8'hBA, 8'h78, 8'h25, 8'h2E, 8'h1C, 8'hA6, 8'hB4, 8'hC6,
    8'hE8, 8'hDD, 8'h74, 8'h1F, 8'h4B, 8'hBD, 8'h8B, 8'h8A,

    8'h70, 8'h3E, 8'hB5, 8'h66, 8'h48, 8'h03, 8'hF6, 8'h0E,
    8'h61, 8'h35, 8'h57, 8'hB9, 8'h86, 8'hC1, 8'h1D, 8'h9E,

    8'hE1, 8'hF8, 8'h98, 8'h11, 8'h69, 8'hD9, 8'h8E, 8'h94,
    8'h9B, 8'h1E, 8'h87, 8'hE9, 8'hCE, 8'h55, 8'h28, 8'hDF,

    8'h8C, 8'hA1, 8'h89, 8'h0D, 8'hBF, 8'hE6, 8'h42, 8'h68,
    8'h41, 8'h99, 8'h2D, 8'h0F, 8'hB0, 8'h54, 8'hBB, 8'h16
  };

  localparam logic [7:0] SBOX_INV [256] = '{
    8'h52, 8'h09, 8'h6a, 8'hd5, 8'h30, 8'h36, 8'ha5, 8'h38,
    8'hbf, 8'h40, 8'ha3, 8'h9e, 8'h81, 8'hf3, 8'hd7, 8'hfb,

    8'h7c, 8'he3, 8'h39, 8'h82, 8'h9b, 8'h2f, 8'hff, 8'h87,
    8'h34, 8'h8e, 8'h43, 8'h44, 8'hc4, 8'hde, 8'he9, 8'hcb,

    8'h54, 8'h7b, 8'h94, 8'h32, 8'ha6, 8'hc2, 8'h23, 8'h3d,
    8'hee, 8'h4c, 8'h95, 8'h0b, 8'h42, 8'hfa, 8'hc3, 8'h4e,

    8'h08, 8'h2e, 8'ha1, 8'h66, 8'h28, 8'hd9, 8'h24, 8'hb2,
    8'h76, 8'h5b, 8'ha2, 8'h49, 8'h6d, 8'h8b, 8'hd1, 8'h25,

    8'h72, 8'hf8, 8'hf6, 8'h64, 8'h86, 8'h68, 8'h98, 8'h16,
    8'hd4, 8'ha4, 8'h5c, 8'hcc, 8'h5d, 8'h65, 8'hb6, 8'h92,

    8'h6c, 8'h70, 8'h48, 8'h50, 8'hfd, 8'hed, 8'hb9, 8'hda,
    8'h5e, 8'h15, 8'h46, 8'h57, 8'ha7, 8'h8d, 8'h9d, 8'h84,

    8'h90, 8'hd8, 8'hab, 8'h00, 8'h8c, 8'hbc, 8'hd3, 8'h0a,
    8'hf7, 8'he4, 8'h58, 8'h05, 8'hb8, 8'hb3, 8'h45, 8'h06,

    8'hd0, 8'h2c, 8'h1e, 8'h8f, 8'hca, 8'h3f, 8'h0f, 8'h02,
    8'hc1, 8'haf, 8'hbd, 8'h03, 8'h01, 8'h13, 8'h8a, 8'h6b,

    8'h3a, 8'h91, 8'h11, 8'h41, 8'h4f, 8'h67, 8'hdc, 8'hea,
    8'h97, 8'hf2, 8'hcf, 8'hce, 8'hf0, 8'hb4, 8'he6, 8'h73,

    8'h96, 8'hac, 8'h74, 8'h22, 8'he7, 8'had, 8'h35, 8'h85,
    8'he2, 8'hf9, 8'h37, 8'he8, 8'h1c, 8'h75, 8'hdf, 8'h6e,

    8'h47, 8'hf1, 8'h1a, 8'h71, 8'h1d, 8'h29, 8'hc5, 8'h89,
    8'h6f, 8'hb7, 8'h62, 8'h0e, 8'haa, 8'h18, 8'hbe, 8'h1b,

    8'hfc, 8'h56, 8'h3e, 8'h4b, 8'hc6, 8'hd2, 8'h79, 8'h20,
    8'h9a, 8'hdb, 8'hc0, 8'hfe, 8'h78, 8'hcd, 8'h5a, 8'hf4,

    8'h1f, 8'hdd, 8'ha8, 8'h33, 8'h88, 8'h07, 8'hc7, 8'h31,
    8'hb1, 8'h12, 8'h10, 8'h59, 8'h27, 8'h80, 8'hec, 8'h5f,

    8'h60, 8'h51, 8'h7f, 8'ha9, 8'h19, 8'hb5, 8'h4a, 8'h0d,
    8'h2d, 8'he5, 8'h7a, 8'h9f, 8'h93, 8'hc9, 8'h9c, 8'hef,

    8'ha0, 8'he0, 8'h3b, 8'h4d, 8'hae, 8'h2a, 8'hf5, 8'hb0,
    8'hc8, 8'heb, 8'hbb, 8'h3c, 8'h83, 8'h53, 8'h99, 8'h61,

    8'h17, 8'h2b, 8'h04, 8'h7e, 8'hba, 8'h77, 8'hd6, 8'h26,
    8'he1, 8'h69, 8'h14, 8'h63, 8'h55, 8'h21, 8'h0c, 8'h7d
  };

  // Drive output
  assign data_o = (op_i == CIPH_FWD) ? SBOX_FWD[data_i] :
                  (op_i == CIPH_INV) ? SBOX_INV[data_i] : SBOX_FWD[data_i];

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES Canright SBox package
//
// For details, see the following documents:
// - Canright, "A very compact Rijndael S-box", technical report
//   available at https://hdl.handle.net/10945/25608
// - Canright, "A very compact 'perfectly masked' S-box for AES (corrected)", paper
//   available at https://eprint.iacr.org/2009/011.pdf

package aes_sbox_canright_pkg;

  // Multiplication in GF(2^2), using normal basis [Omega^2, Omega]
  // (see Figure 14 in the technical report)
  function automatic logic [1:0] aes_mul_gf2p2(logic [1:0] g, logic [1:0] d);
    logic [1:0] f;
    logic       a, b, c;
    a    = g[1] & d[1];
    b    = (^g) & (^d);
    c    = g[0] & d[0];
    f[1] = a ^ b;
    f[0] = c ^ b;
    return f;
  endfunction

  // Scale by Omega^2 = N in GF(2^2), using normal basis [Omega^2, Omega]
  // (see Figure 16 in the technical report)
  function automatic logic [1:0] aes_scale_omega2_gf2p2(logic [1:0] g);
    logic [1:0] d;
    d[1] = g[0];
    d[0] = g[1] ^ g[0];
    return d;
  endfunction

  // Scale by Omega = N^2 in GF(2^2), using normal basis [Omega^2, Omega]
  // (see Figure 15 in the technical report)
  function automatic logic [1:0] aes_scale_omega_gf2p2(logic [1:0] g);
    logic [1:0] d;
    d[1] = g[1] ^ g[0];
    d[0] = g[1];
    return d;
  endfunction

  // Square in GF(2^2), using normal basis [Omega^2, Omega]
  // (see Figures 8 and 10 in the technical report)
  function automatic logic [1:0] aes_square_gf2p2(logic [1:0] g);
    logic [1:0] d;
    d[1] = g[0];
    d[0] = g[1];
    return d;
  endfunction

  // Multiplication in GF(2^4), using normal basis [alpha^8, alpha^2]
  // (see Figure 13 in the technical report)
  function automatic logic [3:0] aes_mul_gf2p4(logic [3:0] gamma, logic [3:0] delta);
    logic [3:0] theta;
    logic [1:0] a, b, c;
    a          = aes_mul_gf2p2(gamma[3:2], delta[3:2]);
    b          = aes_mul_gf2p2(gamma[3:2] ^ gamma[1:0], delta[3:2] ^ delta[1:0]);
    c          = aes_mul_gf2p2(gamma[1:0], delta[1:0]);
    theta[3:2] = a ^ aes_scale_omega2_gf2p2(b);
    theta[1:0] = c ^ aes_scale_omega2_gf2p2(b);
    return theta;
  endfunction

  // Square and scale by nu in GF(2^4)/GF(2^2), using normal basis [alpha^8, alpha^2]
  // (see Figure 19 as well as Appendix A of the technical report)
  function automatic logic [3:0] aes_square_scale_gf2p4_gf2p2(logic [3:0] gamma);
    logic [3:0] delta;
    logic [1:0] a, b;
    a          = gamma[3:2] ^ gamma[1:0];
    b          = aes_square_gf2p2(gamma[1:0]);
    delta[3:2] = aes_square_gf2p2(a);
    delta[1:0] = aes_scale_omega_gf2p2(b);
    return delta;
  endfunction

  // Basis conversion matrices to convert between polynomial basis A, normal basis X
  // and basis S incorporating the bit matrix of the SBox. More specifically,
  // multiplication by X2X performs the transformation from normal basis X into
  // polynomial basis A, followed by the affine transformation (substep 2). Likewise,
  // multiplication by S2X performs the inverse affine transformation followed by the
  // transformation from polynomial basis A to normal basis X.
  // (see Appendix A of the technical report)
  parameter logic [7:0] A2X [8] = '{8'h98, 8'hf3, 8'hf2, 8'h48, 8'h09, 8'h81, 8'ha9, 8'hff};
  parameter logic [7:0] X2A [8] = '{8'h64, 8'h78, 8'h6e, 8'h8c, 8'h68, 8'h29, 8'hde, 8'h60};
  parameter logic [7:0] X2S [8] = '{8'h58, 8'h2d, 8'h9e, 8'h0b, 8'hdc, 8'h04, 8'h03, 8'h24};
  parameter logic [7:0] S2X [8] = '{8'h8c, 8'h79, 8'h05, 8'heb, 8'h12, 8'h04, 8'h51, 8'h53};

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES Canright SBox #4
//
// For details, see the technical report: Canright, "A very compact Rijndael S-box"
// available at https://hdl.handle.net/10945/25608

module aes_sbox_canright (
  input  aes_pkg::ciph_op_e op_i,
  input  logic [7:0]        data_i,
  output logic [7:0]        data_o
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  ///////////////
  // Functions //
  ///////////////

  // Inverse in GF(2^4), using normal basis [alpha^8, alpha^2]
  // (see Figure 12 in the technical report)
  function automatic logic [3:0] aes_inverse_gf2p4(logic [3:0] gamma);
    logic [3:0] delta;
    logic [1:0] a, b, c, d;
    a          = gamma[3:2] ^ gamma[1:0];
    b          = aes_mul_gf2p2(gamma[3:2], gamma[1:0]);
    c          = aes_scale_omega2_gf2p2(aes_square_gf2p2(a));
    d          = aes_square_gf2p2(c ^ b);
    delta[3:2] = aes_mul_gf2p2(d, gamma[1:0]);
    delta[1:0] = aes_mul_gf2p2(d, gamma[3:2]);
    return delta;
  endfunction

  // Inverse in GF(2^8), using normal basis [d^16, d]
  // (see Figure 11 in the technical report)
  function automatic logic [7:0] aes_inverse_gf2p8(logic [7:0] gamma);
    logic [7:0] delta;
    logic [3:0] a, b, c, d;
    a          = gamma[7:4] ^ gamma[3:0];
    b          = aes_mul_gf2p4(gamma[7:4], gamma[3:0]);
    c          = aes_square_scale_gf2p4_gf2p2(a);
    d          = aes_inverse_gf2p4(c ^ b);
    delta[7:4] = aes_mul_gf2p4(d, gamma[3:0]);
    delta[3:0] = aes_mul_gf2p4(d, gamma[7:4]);
    return delta;
  endfunction

  ///////////////////
  // Canright SBox //
  ///////////////////

  logic [7:0] data_basis_x, data_inverse;

  // Convert to normal basis X.
  assign data_basis_x = (op_i == CIPH_FWD) ? aes_mvm(data_i, A2X)         :
                        (op_i == CIPH_INV) ? aes_mvm(data_i ^ 8'h63, S2X) :
                                             aes_mvm(data_i, A2X);

  // Do the inversion in normal basis X.
  assign data_inverse = aes_inverse_gf2p8(data_basis_x);

  // Convert to basis S or A.
  assign data_o       = (op_i == CIPH_FWD) ? aes_mvm(data_inverse, X2S) ^ 8'h63 :
                        (op_i == CIPH_INV) ? aes_mvm(data_inverse, X2A) :
                                             aes_mvm(data_inverse, X2S) ^ 8'h63;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES Masked Canright SBox without Mask Re-Use
//
// For details, see the following paper:
// Canright, "A very compact 'perfectly masked' S-box for AES (corrected)"
// available at https://eprint.iacr.org/2009/011.pdf
//
// Note: This module implements the original masked inversion algorithm without re-using masks.
// For details, see Section 2.2 of the paper. In addition, a formal analysis using REBECCA (stable
// mode) shows that the intermediate masks cannot be created by re-using bits from the input and
// output masks. Instead, fresh random bits need to be used for these intermediate masks. Still,
// the implmentation cannot be made to pass formal analysis in transient mode. It's usage is thus
// discouraged. It's included here mainly for reference.
//
// For details on the REBECCA tool, see the following paper:
// Bloem, "Formal verification of masked hardware implementations in the presence of glitches"
// available at https://eprint.iacr.org/2017/897.pdf

///////////////////////////////////////////////////////////////////////////////////////////////////
// IMPORTANT NOTE:                                                                               //
//                            DO NOT USE THIS FOR SYNTHESIS BLINDLY!                             //
//                                                                                               //
// This implementation relies on primitive cells like prim_buf containing tool-specific          //
// synthesis attributes to enforce the correct ordering of operations and avoid aggressive       //
// optimization. Without the proper primitives, synthesis tools might heavily optimize the       //
// design. The result is likely insecure. Use with care.                                         //
///////////////////////////////////////////////////////////////////////////////////////////////////

// Masked inverse in GF(2^4), using normal basis [z^4, z]
// (see Formulas 6, 13, 14, 15, 16, 17 in the paper)
module aes_masked_inverse_gf2p4_noreuse (
  input  logic [3:0] b,
  input  logic [3:0] q,
  input  logic [1:0] r,
  input  logic [3:0] t,
  output logic [3:0] b_inv
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  logic [1:0] b1, b0, q1, q0, c_inv, r_sq, t1, t0;
  assign b1 = b[3:2];
  assign b0 = b[1:0];
  assign q1 = q[3:2];
  assign q0 = q[1:0];
  assign t1 = t[3:2];
  assign t0 = t[1:0];

  ////////////////
  // Formula 13 //
  ////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // c = r ^ aes_scale_omega2_gf2p2(aes_square_gf2p2(b1 ^ b0))
  //       ^ aes_scale_omega2_gf2p2(aes_square_gf2p2(q1 ^ q0))
  //       ^ aes_mul_gf2p2(b1, b0)
  //       ^ aes_mul_gf2p2(b1, q0) ^ aes_mul_gf2p2(b0, q1) ^ aes_mul_gf2p2(q1, q0);

  // Get intermediate terms.
  logic [1:0] scale_omega2_b, scale_omega2_q;
  logic [1:0] mul_b1_b0, mul_b1_q0, mul_b0_q1, mul_q1_q0;
  assign scale_omega2_b = aes_scale_omega2_gf2p2(aes_square_gf2p2(b1 ^ b0));
  assign scale_omega2_q = aes_scale_omega2_gf2p2(aes_square_gf2p2(q1 ^ q0));
  assign mul_b1_b0 = aes_mul_gf2p2(b1, b0);
  assign mul_b1_q0 = aes_mul_gf2p2(b1, q0);
  assign mul_b0_q1 = aes_mul_gf2p2(b0, q1);
  assign mul_q1_q0 = aes_mul_gf2p2(q1, q0);

  // These terms are added to other terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [1:0] scale_omega2_b_buf, scale_omega2_q_buf;
  prim_buf #(
    .Width ( 4 )
  ) u_prim_buf_scale_omega2_bq (
    .in_i  ( {scale_omega2_b,     scale_omega2_q}     ),
    .out_o ( {scale_omega2_b_buf, scale_omega2_q_buf} )
  );
  logic [1:0] mul_b1_b0_buf, mul_b1_q0_buf, mul_b0_q1_buf, mul_q1_q0_buf;
  prim_buf #(
    .Width ( 8 )
  ) u_prim_buf_mul_bq01 (
    .in_i  ( {mul_b1_b0,     mul_b1_q0,     mul_b0_q1,     mul_q1_q0}     ),
    .out_o ( {mul_b1_b0_buf, mul_b1_q0_buf, mul_b0_q1_buf, mul_q1_q0_buf} )
  );

  // Generate c step by step.
  logic [1:0] c [6];
  logic [1:0] c_buf [6];
  assign c[0] = r        ^ scale_omega2_b_buf;
  assign c[1] = c_buf[0] ^ scale_omega2_q_buf;
  assign c[2] = c_buf[1] ^ mul_b1_b0_buf;
  assign c[3] = c_buf[2] ^ mul_b1_q0_buf;
  assign c[4] = c_buf[3] ^ mul_b0_q1_buf;
  assign c[5] = c_buf[4] ^ mul_q1_q0_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 6; i++) begin : gen_c_buf
    prim_buf #(
      .Width ( 2 )
    ) u_prim_buf_c_i (
      .in_i  ( c[i]     ),
      .out_o ( c_buf[i] )
    );
  end

  ////////////////////////
  // Formulas 14 and 15 //
  ////////////////////////
  // Note: aes_square_gf2p2 contains no logic, it's just a bit swap. There is no need to insert
  // additional buffers to stop aggressive synthesis optimizations here.
  assign c_inv = aes_square_gf2p2(c_buf[5]);
  assign r_sq  = aes_square_gf2p2(r);

  ////////////////////////
  // Formulas 16 and 17 //
  ////////////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // b1_inv = t1 ^ aes_mul_gf2p2(b0, c_inv)
  //             ^ aes_mul_gf2p2(b0, r_sq) ^ aes_mul_gf2p2(q0, c_inv) ^ aes_mul_gf2p2(q0, r_sq);
  // b0_inv = t0 ^ aes_mul_gf2p2(b1, c_inv)
  //             ^ aes_mul_gf2p2(b1, r_sq) ^ aes_mul_gf2p2(q1, c_inv) ^ aes_mul_gf2p2(q1, r_sq);

  // Get intermediate terms.
  logic [1:0] mul_b0_r_sq, mul_q0_c_inv, mul_q0_r_sq;
  logic [1:0] mul_b1_r_sq, mul_q1_c_inv, mul_q1_r_sq;
  assign mul_b0_r_sq  = aes_mul_gf2p2(b0, r_sq);
  assign mul_q0_c_inv = aes_mul_gf2p2(q0, c_inv);
  assign mul_q0_r_sq  = aes_mul_gf2p2(q0, r_sq);
  assign mul_b1_r_sq  = aes_mul_gf2p2(b1, r_sq);
  assign mul_q1_c_inv = aes_mul_gf2p2(q1, c_inv);
  assign mul_q1_r_sq  = aes_mul_gf2p2(q1, r_sq);

  // The multiplier outputs are added to terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [1:0] mul_b0_r_sq_buf, mul_q0_c_inv_buf, mul_q0_r_sq_buf;
  prim_buf #(
    .Width ( 6 )
  ) u_prim_buf_mul_bq0 (
    .in_i  ( {mul_b0_r_sq,     mul_q0_c_inv,     mul_q0_r_sq}     ),
    .out_o ( {mul_b0_r_sq_buf, mul_q0_c_inv_buf, mul_q0_r_sq_buf} )
  );
  logic [1:0] mul_b1_r_sq_buf, mul_q1_c_inv_buf, mul_q1_r_sq_buf;
  prim_buf #(
    .Width ( 6 )
  ) u_prim_buf_mul_bq1 (
    .in_i  ( {mul_b1_r_sq,     mul_q1_c_inv,     mul_q1_r_sq}     ),
    .out_o ( {mul_b1_r_sq_buf, mul_q1_c_inv_buf, mul_q1_r_sq_buf} )
  );

  // Generate b1_inv and b0_inv step by step.
  logic [1:0] b1_inv [4];
  logic [1:0] b1_inv_buf [4];
  logic [1:0] b0_inv [4];
  logic [1:0] b0_inv_buf [4];
  assign b1_inv[0] = t1            ^ aes_mul_gf2p2(b0, c_inv); // t1 does not depend on b0, c_inv.
  assign b1_inv[1] = b1_inv_buf[0] ^ mul_b0_r_sq_buf;
  assign b1_inv[2] = b1_inv_buf[1] ^ mul_q0_c_inv_buf;
  assign b1_inv[3] = b1_inv_buf[2] ^ mul_q0_r_sq_buf;
  assign b0_inv[0] = t0            ^ aes_mul_gf2p2(b1, c_inv); // t0 does not depend on b1, c_inv.
  assign b0_inv[1] = b0_inv_buf[0] ^ mul_b1_r_sq_buf;
  assign b0_inv[2] = b0_inv_buf[1] ^ mul_q1_c_inv_buf;
  assign b0_inv[3] = b0_inv_buf[2] ^ mul_q1_r_sq_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 4; i++) begin : gen_a01_inv_buf
    prim_buf #(
      .Width ( 2 )
    ) u_prim_buf_b1_inv_i (
      .in_i  ( b1_inv[i]     ),
      .out_o ( b1_inv_buf[i] )
    );
    prim_buf #(
      .Width ( 2 )
    ) u_prim_buf_b0_inv_i (
      .in_i  ( b0_inv[i]     ),
      .out_o ( b0_inv_buf[i] )
    );
  end

  // Note: b_inv is masked by t, b was masked by q.
  assign b_inv = {b1_inv_buf[3], b0_inv_buf[3]};

endmodule

// Masked inverse in GF(2^8), using normal basis [y^16, y]
// (see Formulas 3, 12, 18 and 19 in the paper)
module aes_masked_inverse_gf2p8_noreuse (
  input  logic [7:0] a,    // input data masked by m
  input  logic [7:0] m,    // input mask
  input  logic [7:0] n,    // output mask
  input  logic [9:0] prd,  // pseudo-random data, e.g. for intermediate masks
  output logic [7:0] a_inv // output data masked by n
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  logic [3:0] a1, a0, m1, m0, q, b_inv, s1, s0, t;
  logic [1:0] r;

  assign a1 = a[7:4];
  assign a0 = a[3:0];
  assign m1 = m[7:4];
  assign m0 = m[3:0];

  ////////////////////
  // Notes on masks //
  ////////////////////
  // The paper states the following.
  // r:
  // - must be independent of q,
  // - it is suggested to re-use bits of m,
  // - but further analysis shows that this is not sufficient (see below).
  //
  // q:
  // - must be independent of m.
  //
  // t:
  // - must be independent of r,
  // - must be independent of m (for the final steps involving s),
  // - t1 must be independent of q0, t0 must be independent of q1,
  // - it is suggested to use t = q,
  // - but further analysis shows that this is not sufficient (see below).
  //
  // s:
  // - must be independent of t,
  // - s1 must be independent of m0, s0 must be independent of m1,
  // - it is suggested to use s = m,
  // - but further analysis shows that this is not sufficient (see below).
  //
  // Formally analyzing the implementation with REBECCA reveals that:
  // 1. Fresh random bits are required for r, q and t. Any re-use of other mask bits from m or n
  //    causes the static check to fail.
  // 2. s can be the specified output mask n.
  assign r  = prd[1:0];
  assign q  = prd[5:2];
  assign t  = prd[9:6];
  assign s1 = n[7:4];
  assign s0 = n[3:0];

  ////////////////
  // Formula 12 //
  ////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // b = q ^ aes_square_scale_gf2p4_gf2p2(a1 ^ a0)
  //       ^ aes_square_scale_gf2p4_gf2p2(m1 ^ m0)
  //       ^ aes_mul_gf2p4(a1, a0)
  //       ^ aes_mul_gf2p4(a1, m0) ^ aes_mul_gf2p4(a0, m1) ^ aes_mul_gf2p4(m0, m1);

  // Get intermediate terms.
  logic [3:0] ss_a1_a0, ss_m1_m0;
  assign ss_a1_a0 = aes_square_scale_gf2p4_gf2p2(a1 ^ a0);
  assign ss_m1_m0 = aes_square_scale_gf2p4_gf2p2(m1 ^ m0);

  logic [3:0] mul_a1_a0, mul_a1_m0, mul_a0_m1, mul_m0_m1;
  assign mul_a1_a0 = aes_mul_gf2p4(a1, a0);
  assign mul_a1_m0 = aes_mul_gf2p4(a1, m0);
  assign mul_a0_m1 = aes_mul_gf2p4(a0, m1);
  assign mul_m0_m1 = aes_mul_gf2p4(m0, m1);

  // The multiplier outputs are added to terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [3:0] mul_a1_a0_buf, mul_a1_m0_buf, mul_a0_m1_buf, mul_m0_m1_buf;
  prim_buf #(
    .Width ( 16 )
  ) u_prim_buf_mul_am01 (
    .in_i  ( {mul_a1_a0,     mul_a1_m0,     mul_a0_m1,     mul_m0_m1}     ),
    .out_o ( {mul_a1_a0_buf, mul_a1_m0_buf, mul_a0_m1_buf, mul_m0_m1_buf} )
  );

  // Generate b step by step.
  logic [3:0] b [6];
  logic [3:0] b_buf [6];
  assign b[0] = q        ^ ss_a1_a0; // q does not depend on a1, a0.
  assign b[1] = b_buf[0] ^ ss_m1_m0; // b[0] does not depend on m1, m0.
  assign b[2] = b_buf[1] ^ mul_a1_a0_buf;
  assign b[3] = b_buf[2] ^ mul_a1_m0_buf;
  assign b[4] = b_buf[3] ^ mul_a0_m1_buf;
  assign b[5] = b_buf[4] ^ mul_m0_m1_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 6; i++) begin : gen_b_buf
    prim_buf #(
      .Width ( 4 )
    ) u_prim_buf_b_i (
      .in_i  ( b[i]     ),
      .out_o ( b_buf[i] )
    );
  end

  //////////////////////
  // GF(2^4) Inverter //
  //////////////////////

  // b is masked by q, b_inv is masked by t.
  aes_masked_inverse_gf2p4_noreuse u_aes_masked_inverse_gf2p4 (
    .b     ( b_buf[5] ),
    .q     ( q        ),
    .r     ( r        ),
    .t     ( t        ),
    .b_inv ( b_inv    )
  );

  // The output of the inverse over GF(2^4) and signals derived from that are again recombined
  // with inputs to the GF(2^4) inverter. Aggressive synthesis optimizations across the GF(2^4)
  // inverter may result in SCA leakage and should be avoided.
  logic [3:0] b_inv_buf;
  prim_buf #(
    .Width ( 4 )
  ) u_prim_buf_b_inv (
    .in_i  ( b_inv     ),
    .out_o ( b_inv_buf )
  );

  ////////////////////////
  // Formulas 18 and 19 //
  ////////////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // a1_inv = s1 ^ aes_mul_gf2p4(a0, b_inv)
  //             ^ aes_mul_gf2p4(a0, t) ^ aes_mul_gf2p4(m0, b_inv) ^ aes_mul_gf2p4(m0, t);
  // a0_inv = s0 ^ aes_mul_gf2p4(a1, b_inv)
  //             ^ aes_mul_gf2p4(a1, t) ^ aes_mul_gf2p4(m1, b_inv) ^ aes_mul_gf2p4(m1, t);

  // Get intermediate terms.
  logic [3:0] mul_a0_b_inv, mul_a0_t, mul_m0_b_inv, mul_m0_t;
  logic [3:0] mul_a1_b_inv, mul_a1_t, mul_m1_b_inv, mul_m1_t;
  assign mul_a0_b_inv = aes_mul_gf2p4(a0, b_inv_buf);
  assign mul_a0_t     = aes_mul_gf2p4(a0, t);
  assign mul_m0_b_inv = aes_mul_gf2p4(m0, b_inv_buf);
  assign mul_m0_t     = aes_mul_gf2p4(m0, t);
  assign mul_a1_b_inv = aes_mul_gf2p4(a1, b_inv_buf);
  assign mul_a1_t     = aes_mul_gf2p4(a1, t);
  assign mul_m1_b_inv = aes_mul_gf2p4(m1, b_inv_buf);
  assign mul_m1_t     = aes_mul_gf2p4(m1, t);

  // The multiplier outputs are added to terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [3:0] mul_a0_b_inv_buf, mul_a0_t_buf, mul_m0_b_inv_buf, mul_m0_t_buf;
  prim_buf #(
    .Width ( 16 )
  ) u_prim_buf_mul_am0 (
    .in_i  ( {mul_a0_b_inv,     mul_a0_t,     mul_m0_b_inv,     mul_m0_t}     ),
    .out_o ( {mul_a0_b_inv_buf, mul_a0_t_buf, mul_m0_b_inv_buf, mul_m0_t_buf} )
  );
  logic [3:0] mul_a1_b_inv_buf, mul_a1_t_buf, mul_m1_b_inv_buf, mul_m1_t_buf;
  prim_buf #(
    .Width ( 16 )
  ) u_prim_buf_mul_am1 (
    .in_i  ( {mul_a1_b_inv,     mul_a1_t,     mul_m1_b_inv,     mul_m1_t}     ),
    .out_o ( {mul_a1_b_inv_buf, mul_a1_t_buf, mul_m1_b_inv_buf, mul_m1_t_buf} )
  );

  // Generate a1_inv and a0_inv step by step.
  logic [3:0] a1_inv [4];
  logic [3:0] a1_inv_buf [4];
  logic [3:0] a0_inv [4];
  logic [3:0] a0_inv_buf [4];
  assign a1_inv[0] = s1            ^ mul_a0_b_inv_buf;
  assign a1_inv[1] = a1_inv_buf[0] ^ mul_a0_t_buf;
  assign a1_inv[2] = a1_inv_buf[1] ^ mul_m0_b_inv_buf;
  assign a1_inv[3] = a1_inv_buf[2] ^ mul_m0_t_buf;
  assign a0_inv[0] = s0            ^ mul_a1_b_inv_buf;
  assign a0_inv[1] = a0_inv_buf[0] ^ mul_a1_t_buf;
  assign a0_inv[2] = a0_inv_buf[1] ^ mul_m1_b_inv_buf;
  assign a0_inv[3] = a0_inv_buf[2] ^ mul_m1_t_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 4; i++) begin : gen_a01_inv_buf
    prim_buf #(
      .Width ( 4 )
    ) u_prim_buf_a1_inv_i (
      .in_i  ( a1_inv[i]     ),
      .out_o ( a1_inv_buf[i] )
    );
    prim_buf #(
      .Width ( 4 )
    ) u_prim_buf_a0_inv_i (
      .in_i  ( a0_inv[i]     ),
      .out_o ( a0_inv_buf[i] )
    );
  end

  // Note: a_inv is masked by s (= n), a was masked by m.
  assign a_inv = {a1_inv_buf[3], a0_inv_buf[3]};

endmodule

// SEC_CM: KEY.MASKING
module aes_sbox_canright_masked_noreuse (
  input  aes_pkg::ciph_op_e op_i,
  input  logic        [7:0] data_i, // masked, the actual input data is data_i ^ mask_i
  input  logic        [7:0] mask_i, // input mask, independent from actual input data
  input  logic       [17:0] prd_i,  // pseudo-random data, for remasking and for intermediate
                                    // masks, must be independent of input mask
  output logic        [7:0] data_o, // masked, the actual output data is data_o ^ mask_o
  output logic        [7:0] mask_o  // output mask
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  //////////////////////////
  // Masked Canright SBox //
  //////////////////////////

  logic [7:0] in_data_basis_x, out_data_basis_x;
  logic [7:0] in_mask_basis_x, out_mask_basis_x;

  // Convert data to normal basis X.
  assign in_data_basis_x = (op_i == CIPH_FWD) ? aes_mvm(data_i, A2X)         :
                           (op_i == CIPH_INV) ? aes_mvm(data_i ^ 8'h63, S2X) :
                                                aes_mvm(data_i, A2X);

  // For the masked Canright SBox with no re-use, the output mask directly corresponds to the
  // LSBs of the pseduo-random data provided as input.
  assign mask_o = prd_i[7:0];

  // The remaining bits are used for intermediate masks.
  logic [9:0] prd_masking;
  assign prd_masking = prd_i[17:8];

  // Convert masks to normal basis X.
  // The addition of constant 8'h63 following the affine transformation is skipped.
  assign in_mask_basis_x  = (op_i == CIPH_FWD) ? aes_mvm(mask_i, A2X) :
                            (op_i == CIPH_INV) ? aes_mvm(mask_i, S2X) :
                                                 aes_mvm(mask_i, A2X);

  // The output mask is converted in the opposite direction.
  assign out_mask_basis_x = (op_i == CIPH_INV) ? aes_mvm(mask_o, A2X) :
                            (op_i == CIPH_FWD) ? aes_mvm(mask_o, S2X) :
                                                 aes_mvm(mask_o, S2X);

  // Do the inversion in normal basis X.
  aes_masked_inverse_gf2p8_noreuse u_aes_masked_inverse_gf2p8 (
    .a     ( in_data_basis_x  ), // input
    .m     ( in_mask_basis_x  ), // input
    .n     ( out_mask_basis_x ), // input
    .prd   ( prd_masking      ), // input
    .a_inv ( out_data_basis_x )  // output
  );

  // Convert to basis S or A.
  assign data_o = (op_i == CIPH_FWD) ? (aes_mvm(out_data_basis_x, X2S) ^ 8'h63) :
                  (op_i == CIPH_INV) ? (aes_mvm(out_data_basis_x, X2A))         :
                                       (aes_mvm(out_data_basis_x, X2S) ^ 8'h63);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES Masked Canright SBox with Mask Re-Use
//
// For details, see the following paper:
// Canright, "A very compact 'perfectly masked' S-box for AES (corrected)"
// available at https://eprint.iacr.org/2009/011.pdf
//
// Note: This module implements the masked inversion algorithm with re-using masks.
// For details, see Section 2.3 of the paper. Re-using masks may make the implementation more
// vulnerable to higher-order differential side-channel analysis, but it remains secure against
// first-order attacks. This implementation is commonly referred to as THE Canright Masked SBox.
//
// A formal analysis using REBECCA (stable and transient mode) shows that this implementation is
// not secure. It's usage is thus discouraged. It's included here mainly for reference.
//
// For details on the REBECCA tool, see the following paper:
// Bloem, "Formal verification of masked hardware implementations in the presence of glitches"
// available at https://eprint.iacr.org/2017/897.pdf

///////////////////////////////////////////////////////////////////////////////////////////////////
// IMPORTANT NOTE:                                                                               //
//                            DO NOT USE THIS FOR SYNTHESIS BLINDLY!                             //
//                                                                                               //
// This implementation relies on primitive cells like prim_buf/xor2 containing tool-specific     //
// synthesis attributes to enforce the correct ordering of operations and avoid aggressive       //
// optimization. Without the proper primitives, synthesis tools might heavily optimize the       //
// design. The result is likely insecure. Use with care.                                         //
///////////////////////////////////////////////////////////////////////////////////////////////////

// Masked inverse in GF(2^4), using normal basis [z^4, z]
// (see Formulas 6, 13, 14, 15, 21, 22, 23, 24 in the paper)
module aes_masked_inverse_gf2p4 (
  input  logic [3:0] b,
  input  logic [3:0] q,
  input  logic [1:0] r,
  input  logic [3:0] m1,
  output logic [3:0] b_inv
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  logic [1:0] b1, b0, q1, q0, c_inv, r_sq, m11, m10;
  assign b1  = b[3:2];
  assign b0  = b[1:0];
  assign q1  = q[3:2];
  assign q0  = q[1:0];
  assign m11 = m1[3:2];
  assign m10 = m1[1:0];

  // Get re-usable intermediate results.
  logic [1:0] mul_b0_q1, mul_b1_q0, mul_q1_q0;
  assign mul_b0_q1 = aes_mul_gf2p2(b0, q1);
  assign mul_b1_q0 = aes_mul_gf2p2(b1, q0);
  assign mul_q1_q0 = aes_mul_gf2p2(q1, q0);

  // Avoid aggressive synthesis optimizations.
  logic [1:0] mul_b0_q1_buf, mul_b1_q0_buf, mul_q1_q0_buf;
  prim_buf #(
    .Width ( 6 )
  ) u_prim_buf_mul_bq01 (
    .in_i  ( {mul_b0_q1,     mul_b1_q0,     mul_q1_q0}     ),
    .out_o ( {mul_b0_q1_buf, mul_b1_q0_buf, mul_q1_q0_buf} )
  );

  ////////////////
  // Formula 13 //
  ////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // c = r ^ aes_scale_omega2_gf2p2(aes_square_gf2p2(b1 ^ b0))
  //       ^ aes_scale_omega2_gf2p2(aes_square_gf2p2(q1 ^ q0))
  //       ^ aes_mul_gf2p2(b1, b0)
  //       ^ mul_b1_q0 ^ mul_b0_q1 ^ mul_q0_q1;

  // Get intermediate terms.
  logic [1:0] scale_omega2_b, scale_omega2_q;
  logic [1:0] mul_b1_b0;
  assign scale_omega2_b = aes_scale_omega2_gf2p2(aes_square_gf2p2(b1 ^ b0));
  assign scale_omega2_q = aes_scale_omega2_gf2p2(aes_square_gf2p2(q1 ^ q0));
  assign mul_b1_b0 = aes_mul_gf2p2(b1, b0);

  // These terms are added to other terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [1:0] scale_omega2_b_buf, scale_omega2_q_buf;
  prim_buf #(
    .Width ( 4 )
  ) u_prim_buf_scale_omega2_bq (
    .in_i  ( {scale_omega2_b,     scale_omega2_q}     ),
    .out_o ( {scale_omega2_b_buf, scale_omega2_q_buf} )
  );
  logic [1:0] mul_b1_b0_buf;
  prim_buf #(
    .Width ( 2 )
  ) u_prim_buf_mul_b1_b0 (
    .in_i  ( mul_b1_b0     ),
    .out_o ( mul_b1_b0_buf )
  );

  // Generate c step by step.
  logic [1:0] c [6];
  logic [1:0] c_buf [6];
  assign c[0] = r        ^ scale_omega2_b_buf;
  assign c[1] = c_buf[0] ^ scale_omega2_q_buf;
  assign c[2] = c_buf[1] ^ mul_b1_b0_buf;
  assign c[3] = c_buf[2] ^ mul_b1_q0_buf;
  assign c[4] = c_buf[3] ^ mul_b0_q1_buf;
  assign c[5] = c_buf[4] ^ mul_q1_q0_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 6; i++) begin : gen_c_buf
    prim_buf #(
      .Width ( 2 )
    ) u_prim_buf_c_i (
      .in_i  ( c[i]     ),
      .out_o ( c_buf[i] )
    );
  end

  ////////////////////////
  // Formulas 14 and 15 //
  ////////////////////////
  // Note: aes_square_gf2p2 contains no logic, it's just a bit swap. There is no need to insert
  // additional buffers to stop aggressive synthesis optimizations here.
  assign c_inv = aes_square_gf2p2(c_buf[5]);
  assign r_sq  = aes_square_gf2p2(r);

  ////////////////////////
  // Formulas 21 and 23 //
  ////////////////////////
  // Re-masking c_inv
  // IMPORTANT: First combine the masks (ops in parens) then apply to c_inv:
  // c_inv  = c_inv ^ (q1 ^ r_sq);
  // c2_inv = c_inv ^ (q0 ^ q1);

  // Get intermediate terms.
  logic [1:0] xor_q1_r_sq, xor_q0_q1, c1_inv, c2_inv;
  prim_xor2 #(
    .Width ( 2 )
  ) u_prim_xor_q1_r_sq (
    .in0_i ( q1          ),
    .in1_i ( r_sq        ),
    .out_o ( xor_q1_r_sq )
  );
  prim_xor2 #(
    .Width ( 2 )
  ) u_prim_xor_q0_q1 (
    .in0_i ( q0        ),
    .in1_i ( q1        ),
    .out_o ( xor_q0_q1 )
  );

  // Generate c1_inv and c2_inv.
  prim_xor2 #(
    .Width ( 2 )
  ) u_prim_c1_inv (
    .in0_i ( xor_q1_r_sq ),
    .in1_i ( c_inv       ),
    .out_o ( c1_inv      )
  );
  prim_xor2 #(
    .Width ( 2 )
  ) u_prim_c2_inv (
    .in0_i ( c1_inv    ),
    .in1_i ( xor_q0_q1 ),
    .out_o ( c2_inv    )
  );

  ////////////////////////
  // Formulas 22 and 24 //
  ////////////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // b1_inv = m11 ^ aes_mul_gf2p2(b0, c1_inv)
  //              ^ mul_b0_q1 ^ aes_mul_gf2p2(q0, c1_inv) ^ mul_q0_q1;
  // b0_inv = m10 ^ aes_mul_gf2p2(b1, c2_inv)
  //              ^ mul_b1_q0 ^ aes_mul_gf2p2(q1, c2_inv) ^ mul_q0_q1;

  // Get intermediate terms.
  logic [1:0] mul_b0_c1_inv, mul_q0_c1_inv, mul_b1_c2_inv, mul_q1_c2_inv;
  assign mul_b0_c1_inv = aes_mul_gf2p2(b0, c1_inv);
  assign mul_q0_c1_inv = aes_mul_gf2p2(q0, c1_inv);
  assign mul_b1_c2_inv = aes_mul_gf2p2(b1, c2_inv);
  assign mul_q1_c2_inv = aes_mul_gf2p2(q1, c2_inv);

  // The multiplier outputs are added to terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [1:0] mul_b0_c1_inv_buf, mul_q0_c1_inv_buf, mul_b1_c2_inv_buf, mul_q1_c2_inv_buf;
  prim_buf #(
    .Width ( 8 )
  ) u_prim_buf_mul_bq01_c12_inv (
    .in_i  ( {mul_b0_c1_inv,     mul_q0_c1_inv,     mul_b1_c2_inv,     mul_q1_c2_inv}     ),
    .out_o ( {mul_b0_c1_inv_buf, mul_q0_c1_inv_buf, mul_b1_c2_inv_buf, mul_q1_c2_inv_buf} )
  );

  // Generate b1_inv and b0_inv step by step.
  logic [1:0] b1_inv [4];
  logic [1:0] b1_inv_buf [4];
  logic [1:0] b0_inv [4];
  logic [1:0] b0_inv_buf [4];
  assign b1_inv[0] = m11           ^ mul_b0_c1_inv_buf;
  assign b1_inv[1] = b1_inv_buf[0] ^ mul_b0_q1_buf;
  assign b1_inv[2] = b1_inv_buf[1] ^ mul_q0_c1_inv_buf;
  assign b1_inv[3] = b1_inv_buf[2] ^ mul_q1_q0_buf;
  assign b0_inv[0] = m10           ^ mul_b1_c2_inv_buf;
  assign b0_inv[1] = b0_inv_buf[0] ^ mul_b1_q0_buf;
  assign b0_inv[2] = b0_inv_buf[1] ^ mul_q1_c2_inv_buf;
  assign b0_inv[3] = b0_inv_buf[2] ^ mul_q1_q0_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 4; i++) begin : gen_a01_inv_buf
    prim_buf #(
      .Width ( 2 )
    ) u_prim_buf_b1_inv_i (
      .in_i  ( b1_inv[i]     ),
      .out_o ( b1_inv_buf[i] )
    );
    prim_buf #(
      .Width ( 2 )
    ) u_prim_buf_b0_inv_i (
      .in_i  ( b0_inv[i]     ),
      .out_o ( b0_inv_buf[i] )
    );
  end

  // Note: b_inv is masked by m1, b was masked by q.
  assign b_inv = {b1_inv_buf[3], b0_inv_buf[3]};
endmodule

// Masked inverse in GF(2^8), using normal basis [y^16, y]
// (see Formulas 3, 12, 25, 26 and 27 in the paper)
module aes_masked_inverse_gf2p8 (
  input  logic [7:0] a,
  input  logic [7:0] m,
  input  logic [7:0] n,
  output logic [7:0] a_inv
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  logic [3:0] a1, a0, m1, m0, q, b_inv, s1, s0;
  logic [1:0] r;

  assign a1 = a[7:4];
  assign a0 = a[3:0];
  assign m1 = m[7:4];
  assign m0 = m[3:0];

  ////////////////////
  // Notes on masks //
  ////////////////////
  // The paper states the following.
  // - r must be independent of q.
  // - q must be independent of m.
  // - s is the specified output mask n.
  assign r = m1[3:2];
  assign q = n[7:4];
  assign s1 = n[7:4];
  assign s0 = n[3:0];

  // Get re-usable intermediate results.
  logic [3:0] mul_a0_m1, mul_a1_m0, mul_m0_m1;
  assign mul_a0_m1 = aes_mul_gf2p4(a0, m1);
  assign mul_a1_m0 = aes_mul_gf2p4(a1, m0);
  assign mul_m0_m1 = aes_mul_gf2p4(m0, m1);

  // Avoid aggressive synthesis optimizations.
  logic [3:0] mul_a0_m1_buf, mul_a1_m0_buf, mul_m0_m1_buf;
  prim_buf #(
    .Width ( 12 )
  ) u_prim_buf_mul_bq01 (
    .in_i  ( {mul_a0_m1,     mul_a1_m0,     mul_m0_m1}     ),
    .out_o ( {mul_a0_m1_buf, mul_a1_m0_buf, mul_m0_m1_buf} )
  );

  ////////////////
  // Formula 12 //
  ////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // b = q ^ aes_square_scale_gf2p4_gf2p2(a1 ^ a0)
  //       ^ aes_square_scale_gf2p4_gf2p2(m1 ^ m0)
  //       ^ aes_mul_gf2p4(a1, a0)
  //       ^ mul_a1_m0 ^ mul_a0_m1 ^ mul_m0_m1;

  // Get intermediate terms.
  logic [3:0] ss_a1_a0, ss_m1_m0;
  assign ss_a1_a0 = aes_square_scale_gf2p4_gf2p2(a1 ^ a0);
  assign ss_m1_m0 = aes_square_scale_gf2p4_gf2p2(m1 ^ m0);

  logic [3:0] mul_a1_a0;
  assign mul_a1_a0 = aes_mul_gf2p4(a1, a0);

  // The multiplier output is added to terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [3:0] mul_a1_a0_buf;
  prim_buf #(
    .Width ( 4 )
  ) u_prim_buf_mul_am01 (
    .in_i  ( mul_a1_a0     ),
    .out_o ( mul_a1_a0_buf )
  );

  // Generate b step by step.
  logic [3:0] b [6];
  logic [3:0] b_buf [6];
  assign b[0] = q        ^ ss_a1_a0; // q does not depend on a1, a0.
  assign b[1] = b_buf[0] ^ ss_m1_m0; // b[0] does not depend on m1, m0.
  assign b[2] = b_buf[1] ^ mul_a1_a0_buf;
  assign b[3] = b_buf[2] ^ mul_a1_m0_buf;
  assign b[4] = b_buf[3] ^ mul_a0_m1_buf;
  assign b[5] = b_buf[4] ^ mul_m0_m1_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 6; i++) begin : gen_b_buf
    prim_buf #(
      .Width ( 4 )
    ) u_prim_buf_b_i (
      .in_i  ( b[i]     ),
      .out_o ( b_buf[i] )
    );
  end

  //////////////////////
  // GF(2^4) Inverter //
  //////////////////////

  // b is masked by q, b_inv is masked by m1.
  aes_masked_inverse_gf2p4 u_aes_masked_inverse_gf2p4 (
    .b     ( b_buf[5] ),
    .q     ( q        ),
    .r     ( r        ),
    .m1    ( m1       ),
    .b_inv ( b_inv    )
  );

  // The output of the inverse over GF(2^4) and signals derived from that are again recombined
  // with inputs to the GF(2^4) inverter. Aggressive synthesis optimizations across the GF(2^4)
  // inverter may result in SCA leakage and should be avoided.
  logic [3:0] b_inv_buf;
  prim_buf #(
    .Width ( 4 )
  ) u_prim_buf_b_inv (
    .in_i  ( b_inv     ),
    .out_o ( b_inv_buf )
  );

  ////////////////
  // Formula 26 //
  ////////////////
  // IMPORTANT: First combine the masks (ops in parens) then apply to b_inv:
  // b2_inv = b_inv ^ (m1 ^ m0);

  // Generate b2_inv step by step.
  logic [3:0] xor_m1_m0, b2_inv;
  prim_xor2 #(
    .Width ( 4 )
  ) u_prim_xor_m1_m0 (
    .in0_i ( m1        ),
    .in1_i ( m0        ),
    .out_o ( xor_m1_m0 )
  );
  prim_xor2 #(
    .Width ( 4 )
  ) u_prim_xor_b2_inv (
    .in0_i ( b_inv_buf ),
    .in1_i ( xor_m1_m0 ),
    .out_o ( b2_inv    )
  );

  ////////////////////////
  // Formulas 25 and 27 //
  ////////////////////////
  // IMPORTANT: The following ops must be executed in order (left to right):
  // a1_inv = s1 ^ aes_mul_gf2p4(a0, b_inv)
  //             ^ mul_a0_m1 ^ aes_mul_gf2p4(m0, b_inv)  ^ mul_m0_m1;
  // a0_inv = s0 ^ aes_mul_gf2p4(a1, b2_inv)
  //             ^ mul_a1_m0 ^ aes_mul_gf2p4(m1, b2_inv) ^ mul_m0_m1;

  // Get intermediate terms.
  logic [3:0] mul_a0_b_inv, mul_m0_b_inv, mul_a1_b2_inv, mul_m1_b2_inv;
  assign mul_a0_b_inv  = aes_mul_gf2p4(a0, b_inv_buf);
  assign mul_m0_b_inv  = aes_mul_gf2p4(m0, b_inv_buf);
  assign mul_a1_b2_inv = aes_mul_gf2p4(a1, b2_inv);
  assign mul_m1_b2_inv = aes_mul_gf2p4(m1, b2_inv);

  // The multiplier outputs are added to terms that depend on the same inputs.
  // Avoid aggressive synthesis optimizations.
  logic [3:0] mul_a0_b_inv_buf, mul_m0_b_inv_buf, mul_a1_b2_inv_buf, mul_m1_b2_inv_buf;
  prim_buf #(
    .Width ( 16 )
  ) u_prim_buf_mul_bq01_c12_inv (
    .in_i  ( {mul_a0_b_inv,     mul_m0_b_inv,     mul_a1_b2_inv,     mul_m1_b2_inv}     ),
    .out_o ( {mul_a0_b_inv_buf, mul_m0_b_inv_buf, mul_a1_b2_inv_buf, mul_m1_b2_inv_buf} )
  );

  // Generate a1_inv and a0_inv step by step.
  logic [3:0] a1_inv [4];
  logic [3:0] a1_inv_buf [4];
  logic [3:0] a0_inv [4];
  logic [3:0] a0_inv_buf [4];
  assign a1_inv[0] = s1            ^ mul_a0_b_inv_buf;
  assign a1_inv[1] = a1_inv_buf[0] ^ mul_a0_m1_buf;
  assign a1_inv[2] = a1_inv_buf[1] ^ mul_m0_b_inv_buf;
  assign a1_inv[3] = a1_inv_buf[2] ^ mul_m0_m1_buf;
  assign a0_inv[0] = s0            ^ mul_a1_b2_inv_buf; // s0 doesn't depend on a1, b2_inv.
  assign a0_inv[1] = a0_inv_buf[0] ^ mul_a1_m0_buf;
  assign a0_inv[2] = a0_inv_buf[1] ^ mul_m1_b2_inv_buf;
  assign a0_inv[3] = a0_inv_buf[2] ^ mul_m0_m1_buf;

  // Avoid aggressive synthesis optimizations.
  for (genvar i = 0; i < 4; i++) begin : gen_a01_inv_buf
    prim_buf #(
      .Width ( 4 )
    ) u_prim_buf_a1_inv_i (
      .in_i  ( a1_inv[i]     ),
      .out_o ( a1_inv_buf[i] )
    );
    prim_buf #(
      .Width ( 4 )
    ) u_prim_buf_a0_inv_i (
      .in_i  ( a0_inv[i]     ),
      .out_o ( a0_inv_buf[i] )
    );
  end

  // Note: a_inv is masked by s (= n), a was masked by m.
  assign a_inv = {a1_inv_buf[3], a0_inv_buf[3]};

endmodule

// SEC_CM: KEY.MASKING
module aes_sbox_canright_masked (
  input  aes_pkg::ciph_op_e op_i,
  input  logic [7:0]        data_i, // masked, the actual input data is data_i ^ mask_i
  input  logic [7:0]        mask_i, // input mask, independent from actual input data
  input  logic [7:0]        prd_i,  // pseudo-random data for remasking, independent of input mask
  output logic [7:0]        data_o, // masked, the actual output data is data_o ^ mask_o
  output logic [7:0]        mask_o  // output mask
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  //////////////////////////
  // Masked Canright SBox //
  //////////////////////////

  logic [7:0] in_data_basis_x, out_data_basis_x;
  logic [7:0] in_mask_basis_x, out_mask_basis_x;

  // Convert data to normal basis X.
  assign in_data_basis_x = (op_i == CIPH_FWD) ? aes_mvm(data_i, A2X)         :
                           (op_i == CIPH_INV) ? aes_mvm(data_i ^ 8'h63, S2X) :
                                                aes_mvm(data_i, A2X);

  // For the masked Canright SBox, the output mask directly corresponds to the pseduo-random data
  // provided as input.
  assign mask_o = prd_i;

  // Convert masks to normal basis X.
  // The addition of constant 8'h63 following the affine transformation is skipped.
  assign in_mask_basis_x  = (op_i == CIPH_FWD) ? aes_mvm(mask_i, A2X) :
                            (op_i == CIPH_INV) ? aes_mvm(mask_i, S2X) :
                                                 aes_mvm(mask_i, A2X);

  // The output mask is converted in the opposite direction.
  assign out_mask_basis_x = (op_i == CIPH_INV) ? aes_mvm(mask_o, A2X) :
                            (op_i == CIPH_FWD) ? aes_mvm(mask_o, S2X) :
                                                 aes_mvm(mask_o, S2X);

  // Do the inversion in normal basis X.
  aes_masked_inverse_gf2p8 u_aes_masked_inverse_gf2p8 (
    .a     ( in_data_basis_x  ), // input
    .m     ( in_mask_basis_x  ), // input
    .n     ( out_mask_basis_x ), // input
    .a_inv ( out_data_basis_x )  // output
  );

  // Convert to basis S or A.
  assign data_o = (op_i == CIPH_FWD) ? (aes_mvm(out_data_basis_x, X2S) ^ 8'h63) :
                  (op_i == CIPH_INV) ? (aes_mvm(out_data_basis_x, X2A))         :
                                       (aes_mvm(out_data_basis_x, X2S) ^ 8'h63);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES S-Box with First-Order Domain-Oriented Masking
//
// This is the unpipelined version using DOM-dep multipliers. It has a latency of 5 clock cycles
// and requires 28 bits of pseudo-random data per evaluation. Pipelining would only be beneficial
// when using
// - either a cipher core architecture with a data path smaller than 128 bit, i.e., where the
//   individual S-Boxes are evaluated more than once per round, or
// - a fully unrolled cipher core architecture for maximum throughput.
//
// Note: The DOM AES S-Box is built on top of the Canright masked S-Box without mask re-use.
//
// For details, see the following papers and reports:
// [1] Gross, "Domain-Oriented Masking: Compact Masked Hardware Implementations with Arbitrary
//     Protection Order" available at https://eprint.iacr.org/2016/486.pdf
// [2] Canright, "A very compact 'perfectly masked' S-box for AES (corrected)" available at
//     https://eprint.iacr.org/2009/011.pdf
// [3] Canright, "A very compact Rijndael S-box" available at https://hdl.handle.net/10945/25608
//
// Using the Coco-Alma tool in transient mode, this implementation has been formally verified to be
// secure against first-order side-channel analysis (SCA). For more information on the tool,
// refer to the following papers:
// [4] Gigerl, "COCO: Co-design and co-verification of masked software implementations on CPUs"
//     available at https://eprint.iacr.org/2020/1294.pdf
// [5] Bloem, "Formal verification of masked hardware implementations in the presence of glitches"
//     available at https://eprint.iacr.org/2017/897.pdf

///////////////////////////////////////////////////////////////////////////////////////////////////
// IMPORTANT NOTE:                                                                               //
//                            DO NOT USE THIS FOR SYNTHESIS BLINDLY!                             //
//                                                                                               //
// This implementation relies on primitive cells like prim_buf/flop_en containing tool-specific  //
// synthesis attributes to prevent the synthesis tool from optimizing away/re-ordering registers //
// and to enforce the correct ordering of operations. Without the proper primitives, synthesis   //
// tools might heavily optimize the design. The result is likely insecure. Use with care.        //
///////////////////////////////////////////////////////////////////////////////////////////////////

`include "prim_assert.sv"

// Packed struct for pseudo-random data (PRD) input. Stages 1, 3 and 4 require 8 bits each. Stage 2
// requires just 4 bits.
typedef struct packed {
  logic [7:0] prd_1;
  logic [3:0] prd_2;
  logic [7:0] prd_3;
  logic [7:0] prd_4;
} prd_in_t;

// Packed struct for pseudo-random data (PRD) output. Stages 2 and 3 produce 8 bits each. Stage 1
// produces just 4 bits.
typedef struct packed {
  logic [3:0] prd_1;
  logic [7:0] prd_2;
  logic [7:0] prd_3;
} prd_out_t;

// DOM-indep GF(2^N) multiplier, first-order masked.
// Computes (a_q ^ b_q) = (a_x ^ b_x) * (a_y ^ b_y), i.e. q = x * y using first-order
// domain-oriented masking. The sharings of x and y are required to be uniformly random and
// independent from each other.
// See Fig. 2 in [1].
module aes_dom_indep_mul_gf2pn #(
  parameter int unsigned NPower   = 4,
  parameter bit          Pipeline = 1'b0
) (
  input  logic              clk_i,
  input  logic              rst_ni,
  input  logic              we_i,
  input  logic [NPower-1:0] a_x,    // Share a of x
  input  logic [NPower-1:0] a_y,    // Share a of y
  input  logic [NPower-1:0] b_x,    // Share b of x
  input  logic [NPower-1:0] b_y,    // Share b of y
  input  logic [NPower-1:0] z_0,    // Randomness for resharing
  output logic [NPower-1:0] a_q,    // Share a of q
  output logic [NPower-1:0] b_q     // Share b of q
);

  import aes_sbox_canright_pkg::*;

  /////////////////
  // Calculation //
  /////////////////
  // Inner-domain terms
  logic [NPower-1:0] mul_ax_ay_d, mul_bx_by_d;
  if (NPower == 4) begin : gen_inner_mul_gf2p4
    assign mul_ax_ay_d = aes_mul_gf2p4(a_x, a_y);
    assign mul_bx_by_d = aes_mul_gf2p4(b_x, b_y);

  end else begin : gen_inner_mul_gf2p2
    assign mul_ax_ay_d = aes_mul_gf2p2(a_x, a_y);
    assign mul_bx_by_d = aes_mul_gf2p2(b_x, b_y);
  end

  // Cross-domain terms
  logic [NPower-1:0] mul_ax_by, mul_ay_bx;
  if (NPower == 4) begin : gen_cross_mul_gf2p4
    assign mul_ax_by = aes_mul_gf2p4(a_x, b_y);
    assign mul_ay_bx = aes_mul_gf2p4(a_y, b_x);

  end else begin : gen_cross_mul_gf2p2
    assign mul_ax_by = aes_mul_gf2p2(a_x, b_y);
    assign mul_ay_bx = aes_mul_gf2p2(a_y, b_x);
  end

  ///////////////
  // Resharing //
  ///////////////
  // Resharing of cross-domain terms
  logic [NPower-1:0] aq_z0_d, bq_z0_d;
  logic [NPower-1:0] aq_z0_q, bq_z0_q;
  assign aq_z0_d = z_0 ^ mul_ax_by;
  assign bq_z0_d = z_0 ^ mul_ay_bx;

  // Registers
  prim_flop_en #(
    .Width      ( 2*NPower ),
    .ResetValue ( '0       )
  ) u_prim_flop_abq_z0 (
    .clk_i  ( clk_i              ),
    .rst_ni ( rst_ni             ),
    .en_i   ( we_i               ),
    .d_i    ( {aq_z0_d, bq_z0_d} ),
    .q_o    ( {aq_z0_q, bq_z0_q} )
  );

  /////////////////////////
  // Optional Pipelining //
  /////////////////////////
  logic [NPower-1:0] mul_ax_ay, mul_bx_by;

  if (Pipeline == 1'b1) begin : gen_pipeline
    // Add pipeline registers on inner-domain terms prior to integration. This allows accepting new
    // input data every clock cycle and prevents SCA leakage occurring due to the integration of
    // reshared cross-domain terms with inner-domain terms derived from different input data.

    logic [NPower-1:0] mul_ax_ay_q, mul_bx_by_q;
    prim_flop_en #(
      .Width      ( 2*NPower ),
      .ResetValue ( '0       )
    ) u_prim_flop_mul_abx_aby (
      .clk_i  ( clk_i                      ),
      .rst_ni ( rst_ni                     ),
      .en_i   ( we_i                       ),
      .d_i    ( {mul_ax_ay_d, mul_bx_by_d} ),
      .q_o    ( {mul_ax_ay_q, mul_bx_by_q} )
    );

    assign mul_ax_ay = mul_ax_ay_q;
    assign mul_bx_by = mul_bx_by_q;

  end else begin : gen_no_pipeline
    // Do not add the optional pipeline registers on the inner-domain terms. This allows to save
    // some area in case the multiplier does not need to accept new data in every cycle. However,
    // this can cause SCA leakage as during the clock cycle in which new data arrives, the new
    // inner-domain terms are integrated with the previous, reshared cross-domain terms.

    // Avoid aggressive synthesis optimizations.
    logic [NPower-1:0] mul_ax_ay_buf, mul_bx_by_buf;
    prim_buf #(
      .Width  ( 2*NPower )
    ) u_prim_buf_mul_abx_aby (
      .in_i  ( {mul_ax_ay_d,   mul_bx_by_d}   ),
      .out_o ( {mul_ax_ay_buf, mul_bx_by_buf} )
    );

    assign mul_ax_ay = mul_ax_ay_buf;
    assign mul_bx_by = mul_bx_by_buf;
  end

  /////////////////
  // Integration //
  /////////////////
  assign a_q = mul_ax_ay ^ aq_z0_q;
  assign b_q = mul_bx_by ^ bq_z0_q;

  // Only GF(2^4) and GF(2^2) is supported.
  `ASSERT_INIT(AesDomIndepMulPower, NPower == 4 || NPower == 2)

endmodule

// DOM-dep GF(2^N) multiplier, first-order masked.
// Computes (a_q ^ b_q) = (a_x ^ b_x) * (a_y ^ b_y), i.e. q = x * y using first-order
// domain-oriented masking. The sharings of x and y are NOT required to be independent from each
// other. This is the un-optimized version consuming 3 times N bits of randomness for blinding and
// resharing. It is not used in the design but we keep it for reference.
// See Fig. 4 and Formulas 8 - 11 in [1].
module aes_dom_dep_mul_gf2pn_unopt #(
  parameter int unsigned NPower   = 4,
  parameter bit          Pipeline = 1'b0
) (
  input  logic              clk_i,
  input  logic              rst_ni,
  input  logic              we_i,
  input  logic [NPower-1:0] a_x,    // Share a of x
  input  logic [NPower-1:0] a_y,    // Share a of y
  input  logic [NPower-1:0] b_x,    // Share b of x
  input  logic [NPower-1:0] b_y,    // Share b of y
  input  logic [NPower-1:0] a_z,    // Randomness for blinding
  input  logic [NPower-1:0] b_z,    // Randomness for blinding
  input  logic [NPower-1:0] z_0,    // Randomness for resharing
  output logic [NPower-1:0] a_q,    // Share a of q
  output logic [NPower-1:0] b_q     // Share b of q
);

  import aes_sbox_canright_pkg::*;

  //////////////
  // Blinding //
  //////////////
  // Blinding of y by z.
  logic [NPower-1:0] a_yz_d, b_yz_d;
  logic [NPower-1:0] a_yz_q, b_yz_q;
  assign a_yz_d = a_y ^ a_z;
  assign b_yz_d = b_y ^ b_z;

  // Registers
  prim_flop_en #(
    .Width      ( 2*NPower ),
    .ResetValue ( '0       )
  ) u_prim_flop_ab_yz (
    .clk_i  ( clk_i            ),
    .rst_ni ( rst_ni           ),
    .en_i   ( we_i             ),
    .d_i    ( {a_yz_d, b_yz_d} ),
    .q_o    ( {a_yz_q, b_yz_q} )
  );

  ////////////////
  // Correction //
  ////////////////
  logic [NPower-1:0] a_mul_x_z, b_mul_x_z;
  aes_dom_indep_mul_gf2pn #(
    .NPower   ( NPower   ),
    .Pipeline ( Pipeline )
  ) u_aes_dom_indep_mul_gf2pn (
    .clk_i  ( clk_i     ),
    .rst_ni ( rst_ni    ),
    .we_i   ( we_i      ),
    .a_x    ( a_x       ), // Share a of x
    .a_y    ( a_z       ), // Share a of z
    .b_x    ( b_x       ), // Share b of x
    .b_y    ( b_z       ), // Share b of z
    .z_0    ( z_0       ), // Randomness for resharing
    .a_q    ( a_mul_x_z ), // Share a of x * z
    .b_q    ( b_mul_x_z )  // Share b of x * z
  );

  /////////////////////////
  // Optional Pipelining //
  /////////////////////////
  logic [NPower-1:0] a_x_calc, b_x_calc;

  if (Pipeline == 1'b1) begin : gen_pipeline
    // Add pipeline registers for input x. This allows accepting new input data every clock cycle
    // and prevents SCA leakage occurring due to the multiplication of input x with b belonging to
    // different clock cycles.

    logic [NPower-1:0] a_x_q, b_x_q;
    prim_flop_en #(
      .Width      ( 2*NPower ),
      .ResetValue ( '0       )
    ) u_prim_flop_ab_x (
      .clk_i  ( clk_i          ),
      .rst_ni ( rst_ni         ),
      .en_i   ( we_i           ),
      .d_i    ( {a_x,   b_x}   ),
      .q_o    ( {a_x_q, b_x_q} )
    );

    assign a_x_calc = a_x_q;
    assign b_x_calc = b_x_q;

  end else begin : gen_no_pipeline
    // Do not add the optional pipeline registers for input x. This allows to save some area in
    // case the multiplier does not need to accept new data in every cycle. However, this can cause
    // SCA leakage as during the clock cycle in which new data arrives, the new x input is
    // multiplied with the previous b.

    assign a_x_calc = a_x;
    assign b_x_calc = b_x;
  end

  /////////////////
  // Calculation //
  /////////////////
  // Combine shares of blinded y to obtain b.
  logic [NPower-1:0] b;
  assign b = a_yz_q ^ b_yz_q;

  logic [NPower-1:0] a_mul_ax_b, b_mul_bx_b;
  if (NPower == 4) begin : gen_mul_gf2p4
    assign a_mul_ax_b = aes_mul_gf2p4(a_x_calc, b);
    assign b_mul_bx_b = aes_mul_gf2p4(b_x_calc, b);

  end else begin : gen_mul_gf2p2
    assign a_mul_ax_b = aes_mul_gf2p2(a_x_calc, b);
    assign b_mul_bx_b = aes_mul_gf2p2(b_x_calc, b);
  end

  /////////////////
  // Integration //
  /////////////////
  assign a_q = a_mul_x_z ^ a_mul_ax_b;
  assign b_q = b_mul_x_z ^ b_mul_bx_b;

  // Only GF(2^4) and GF(2^2) is supported.
  `ASSERT_INIT(AesDomDepMulUnoptPower, NPower == 4 || NPower == 2)

endmodule

// DOM-dep GF(2^N) multiplier, first-order masked.
// Computes (a_q ^ b_q) = (a_x ^ b_x) * (a_y ^ b_y), i.e. q = x * y using first-order
// domain-oriented masking. The sharings of x and y are NOT required to be independent from each
// other. This is the optimized version consuming 2 instead of 3 times N bits of randomness for
// blinding and resharing.
// See Formula 12 in [1].
module aes_dom_dep_mul_gf2pn #(
  parameter int unsigned NPower      = 4,
  parameter bit          Pipeline    = 1'b0,
  parameter bit          PreDomIndep = 1'b0 // 1'b0: Not followed by an un-pipelined DOM-indep
                                            //       multiplier, this enables additional area
                                            //       optimizations
                                            // 1'b1: Directly followed by an un-pipelined
                                            //       DOM-indep multiplier, this is the version
                                            //       discussed in [1].
) (
  input  logic                clk_i,
  input  logic                rst_ni,
  input  logic                we_i,
  input  logic   [NPower-1:0] a_x,    // Share a of x
  input  logic   [NPower-1:0] a_y,    // Share a of y
  input  logic   [NPower-1:0] b_x,    // Share b of x
  input  logic   [NPower-1:0] b_y,    // Share b of y
  input  logic   [NPower-1:0] a_x_q,  // Share a of x, pipelined (for Pipeline=1 or PreDomIndep=1)
  input  logic   [NPower-1:0] a_y_q,  // Share a of y, pipelined (for Pipeline=1)
  input  logic   [NPower-1:0] b_x_q,  // Share b of x, pipelined (for Pipeline=1 or PreDomIndep=1)
  input  logic   [NPower-1:0] b_y_q,  // Share b of y, pipelined (for Pipeline=1)
  input  logic   [NPower-1:0] z_0,    // Randomness for blinding
  input  logic   [NPower-1:0] z_1,    // Randomness for resharing
  output logic   [NPower-1:0] a_q,    // Share a of q
  output logic   [NPower-1:0] b_q,    // Share b of q
  output logic [2*NPower-1:0] prd_o   // Randomness for use in another S-Box instance
);

  import aes_sbox_canright_pkg::*;

  //////////////
  // Blinding //
  //////////////
  // Blinding of y by z_0.
  logic [NPower-1:0] a_yz0_d, b_yz0_d;
  logic [NPower-1:0] a_yz0_q, b_yz0_q;
  assign a_yz0_d = a_y ^ z_0;
  assign b_yz0_d = b_y ^ z_0;

  // Registers
  prim_flop_en #(
    .Width      ( 2*NPower ),
    .ResetValue ( '0       )
  ) u_prim_flop_ab_yz0 (
    .clk_i  ( clk_i              ),
    .rst_ni ( rst_ni             ),
    .en_i   ( we_i               ),
    .d_i    ( {a_yz0_d, b_yz0_d} ),
    .q_o    ( {a_yz0_q, b_yz0_q} )
  );

  ////////////////
  // Correction //
  ////////////////
  // Basically, this a DOM-indep multiplier with:
  // - a_x = a_x, b_x = b_x, and
  // - a_y = z_0, b_y = 0 (constant),
  // which allows for further optimizations.

  // Calculation
  logic [NPower-1:0] mul_ax_z0, mul_bx_z0;
  if (NPower == 4) begin : gen_corr_mul_gf2p4
    assign mul_ax_z0 = aes_mul_gf2p4(a_x, z_0);
    assign mul_bx_z0 = aes_mul_gf2p4(b_x, z_0);

  end else begin : gen_corr_mul_gf2p2
    assign mul_ax_z0 = aes_mul_gf2p2(a_x, z_0);
    assign mul_bx_z0 = aes_mul_gf2p2(b_x, z_0);
  end

  // Avoid aggressive synthesis optimizations.
  logic [NPower-1:0] mul_ax_z0_buf, mul_bx_z0_buf;
  prim_buf #(
    .Width ( 2*NPower )
  ) u_prim_buf_mul_abx_z0 (
    .in_i  ( {mul_ax_z0,     mul_bx_z0}     ),
    .out_o ( {mul_ax_z0_buf, mul_bx_z0_buf} )
  );

  // Resharing
  logic [NPower-1:0] axz0_z1_d, bxz0_z1_d;
  logic [NPower-1:0] axz0_z1_q, bxz0_z1_q;
  assign axz0_z1_d = mul_ax_z0_buf ^ z_1;
  assign bxz0_z1_d = mul_bx_z0_buf ^ z_1;

  // Registers
  prim_flop_en #(
    .Width      ( 2*NPower ),
    .ResetValue ( '0       )
  ) u_prim_flop_abxz0_z1 (
    .clk_i  ( clk_i                  ),
    .rst_ni ( rst_ni                 ),
    .en_i   ( we_i                   ),
    .d_i    ( {axz0_z1_d, bxz0_z1_d} ),
    .q_o    ( {axz0_z1_q, bxz0_z1_q} )
  );

  // Use intermediate results for generating PRD for another S-Box instance.
  // Use one share only. Directly use output of flops updating with we_i.
  // These intermediate results are obtained by remasking b_y and mul_bx_z0 with z_0 and z_1,
  // respectively. Since z_0/1 are uniformly distributed and independent of b_y and mul_bx_z0,
  // the intermediate results are also uniformly distributed and independent of b_y and mul_bx_z0.
  // For details, see Lemma 1 in [2].
  assign prd_o = {b_yz0_q, bxz0_z1_q};

  /////////////////////////
  // Optional Pipelining //
  /////////////////////////
  logic [NPower-1:0] a_x_calc, b_x_calc, a_y_calc, b_y_calc;

  if (Pipeline == 1'b1 && PreDomIndep != 1'b1) begin : gen_pipeline_use
    // Use pipelined inputs x and y. This allows accepting new input data every clock cycle and
    // prevents SCA leakage occurring due to the multiplication of inputs x and y with d_b
    // belonging to different clock cycles.
    //
    // The PreDomIndep variant uses the pipelined inputs directly.

    assign a_x_calc = a_x_q;
    assign b_x_calc = b_x_q;
    assign a_y_calc = a_y_q;
    assign b_y_calc = b_y_q;

  end else begin : gen_no_pipeline_use
    // Do not use pipelined inputs x and y. This allows to save some area in case the multiplier
    // does not need to accept new data in every cycle. However, this can cause SCA leakage as
    // during the clock cycle in which new data arrives, the new x and y inputs are multiplied
    // with the previous d_b.

    assign a_x_calc = a_x;
    assign b_x_calc = b_x;
    assign a_y_calc = a_y;
    assign b_y_calc = b_y;

    // Tie off unused signals.
    if (PreDomIndep != 1'b1) begin : gen_ab_x_q
      logic [NPower-1:0] unused_a_x_q, unused_b_x_q;
      assign unused_a_x_q = a_x_q;
      assign unused_b_x_q = b_x_q;
    end
    logic [NPower-1:0] unused_a_y_q, unused_b_y_q;
    assign unused_a_y_q = a_y_q;
    assign unused_b_y_q = b_y_q;
  end

  ///////////////////////////////
  // Calculation & Integration //
  ///////////////////////////////
  // Compute b. Note that unlike for the unoptimized implementation, we don't combine the blinded
  // shares of y to obtain a single b value. Intstead, every domain d gets its own version of b:
  //
  //   d_b = d_y ^ _D_y_z0
  //
  // where _D_y_z0 corresponds to the sum of all domains of y except for domain d, each
  // individually blinded by z0 (needs to happen before the register bank). This optimization
  // is only suitable for first-order masking.
  // See Formula 12 in [1].

  if (PreDomIndep == 1'b1) begin : gen_pre_dom_indep
    // This DOM-dep multiplier is directly followed by an un-pipelined DOM-indep multiplier. To
    // prevent SCA leakage in the un-pipelined DOM-indep multiplier, the d_y and _D_y_z0 parts of
    // d_b need to be individually multiplied with input x and then the results need to be
    // integrated (summed up) on a per-domain basis.

    // d_y part: Inner-domain terms of x * y
    logic [NPower-1:0] mul_ax_ay_d, mul_bx_by_d;
    logic [NPower-1:0] mul_ax_ay_q, mul_bx_by_q;
    if (NPower == 4) begin : gen_inner_mul_gf2p4
      assign mul_ax_ay_d = aes_mul_gf2p4(a_x_calc, a_y_calc);
      assign mul_bx_by_d = aes_mul_gf2p4(b_x_calc, b_y_calc);

    end else begin : gen_inner_mul_gf2p2
      assign mul_ax_ay_d = aes_mul_gf2p2(a_x_calc, a_y_calc);
      assign mul_bx_by_d = aes_mul_gf2p2(b_x_calc, b_y_calc);
    end

    // Registers
    prim_flop_en #(
      .Width      ( 2*NPower ),
      .ResetValue ( '0       )
    ) u_prim_flop_mul_abx_aby (
      .clk_i  ( clk_i                      ),
      .rst_ni ( rst_ni                     ),
      .en_i   ( we_i                       ),
      .d_i    ( {mul_ax_ay_d, mul_bx_by_d} ),
      .q_o    ( {mul_ax_ay_q, mul_bx_by_q} )
    );

    // _D_y_z0 part: Cross-domain terms: d_x * _D_y_z0
    // Need to use registered version of input x.
    logic [NPower-1:0] mul_ax_byz0, mul_bx_ayz0;
    if (NPower == 4) begin : gen_cross_mul_gf2p4
      assign mul_ax_byz0 = aes_mul_gf2p4(a_x_q, b_yz0_q);
      assign mul_bx_ayz0 = aes_mul_gf2p4(b_x_q, a_yz0_q);

    end else begin : gen_cross_mul_gf2p2
      assign mul_ax_byz0 = aes_mul_gf2p2(a_x_q, b_yz0_q);
      assign mul_bx_ayz0 = aes_mul_gf2p2(b_x_q, a_yz0_q);
    end

    // Avoid aggressive synthesis optimizations.
    logic [NPower-1:0] mul_ax_byz0_buf, mul_bx_ayz0_buf;
    prim_buf #(
      .Width ( 2*NPower )
    ) u_prim_buf_mul_abx_bayz0 (
      .in_i  ( {mul_ax_byz0,     mul_bx_ayz0}     ),
      .out_o ( {mul_ax_byz0_buf, mul_bx_ayz0_buf} )
    );

    // Integration
    assign a_q = axz0_z1_q ^ mul_ax_ay_q ^ mul_ax_byz0_buf;
    assign b_q = bxz0_z1_q ^ mul_bx_by_q ^ mul_bx_ayz0_buf;

  end else begin : gen_not_pre_dom_indep
    // This DOM-dep multiplier is not directly followed by an un-pipelined DOM-indep multiplier. As
    // a result, the d_y and _D_y_z0 parts of d_b can be summed up prior to the multiplication
    // with input x which allows saving 2 GF multipliers.

    // Sum up d_y and _D_y_z0.
    logic [NPower-1:0] a_b, b_b;
    assign a_b = a_y_calc ^ b_yz0_q;
    assign b_b = b_y_calc ^ a_yz0_q;

    // Avoid aggressive synthesis optimizations.
    logic [NPower-1:0] a_b_buf, b_b_buf;
    prim_buf #(
      .Width ( 2*NPower )
    ) u_prim_buf_ab_b (
      .in_i  ( {a_b,     b_b}     ),
      .out_o ( {a_b_buf, b_b_buf} )
    );

    // GF multiplications
    logic [NPower-1:0] a_mul_ax_b, b_mul_bx_b;
    if (NPower == 4) begin : gen_mul_gf2p4
      assign a_mul_ax_b = aes_mul_gf2p4(a_x_calc, a_b_buf);
      assign b_mul_bx_b = aes_mul_gf2p4(b_x_calc, b_b_buf);
    end else begin : gen_mul_gf2p2
      assign a_mul_ax_b = aes_mul_gf2p2(a_x_calc, a_b_buf);
      assign b_mul_bx_b = aes_mul_gf2p2(b_x_calc, b_b_buf);
    end

    // Avoid aggressive synthesis optimizations.
    logic [NPower-1:0] a_mul_ax_b_buf, b_mul_bx_b_buf;
    prim_buf #(
      .Width ( 2*NPower )
    ) u_prim_buf_ab_mul_abx_b (
      .in_i  ( {a_mul_ax_b,     b_mul_bx_b}     ),
      .out_o ( {a_mul_ax_b_buf, b_mul_bx_b_buf} )
    );

    // Integration
    assign a_q = axz0_z1_q ^ a_mul_ax_b_buf;
    assign b_q = bxz0_z1_q ^ b_mul_bx_b_buf;
  end

  // Only GF(2^4) and GF(2^2) is supported.
  `ASSERT_INIT(AesDomDepMulPower, NPower == 4 || NPower == 2)

endmodule

// Inverse in GF(2^4) using first-order domain-oriented masking and normal basis [z^4, z].
// See Fig. 6 in [2] (grey block, Stages 2 and 3) and Formulas 6, 13, 14, 15, 16, 17 in [2].
module aes_dom_inverse_gf2p4 #(
  parameter bit PipelineMul = 1'b1
) (
  input  logic        clk_i,
  input  logic        rst_ni,
  input  logic  [1:0] we_i,
  input  logic  [3:0] a_gamma,
  input  logic  [3:0] b_gamma,
  input  logic  [3:0] prd_2_i,
  input  logic  [7:0] prd_3_i,
  output logic  [3:0] a_gamma_inv,
  output logic  [3:0] b_gamma_inv,
  output logic  [7:0] prd_2_o,
  output logic  [7:0] prd_3_o
);

  import aes_sbox_canright_pkg::*;

  /////////////
  // Stage 2 //
  /////////////
  // Formula 13 in [2].

  logic [1:0] a_gamma1, a_gamma0, b_gamma1, b_gamma0, a_gamma1_gamma0, b_gamma1_gamma0;
  assign a_gamma1 = a_gamma[3:2];
  assign a_gamma0 = a_gamma[1:0];
  assign b_gamma1 = b_gamma[3:2];
  assign b_gamma0 = b_gamma[1:0];

  logic [1:0] a_gamma_ss_d, b_gamma_ss_d;
  logic [1:0] a_gamma_ss_q, b_gamma_ss_q;
  assign a_gamma_ss_d = aes_scale_omega2_gf2p2(aes_square_gf2p2(a_gamma1 ^ a_gamma0));
  assign b_gamma_ss_d = aes_scale_omega2_gf2p2(aes_square_gf2p2(b_gamma1 ^ b_gamma0));
  prim_flop_en #(
    .Width      ( 4  ),
    .ResetValue ( '0 )
  ) u_prim_flop_ab_gamma_ss (
    .clk_i  ( clk_i                        ),
    .rst_ni ( rst_ni                       ),
    .en_i   ( we_i[0]                      ),
    .d_i    ( {a_gamma_ss_d, b_gamma_ss_d} ),
    .q_o    ( {a_gamma_ss_q, b_gamma_ss_q} )
  );

  logic [1:0] a_gamma1_q, a_gamma0_q, b_gamma1_q, b_gamma0_q;
  prim_flop_en #(
    .Width      ( 8  ),
    .ResetValue ( '0 )
  ) u_prim_flop_ab_gamma10 (
    .clk_i  ( clk_i                                            ),
    .rst_ni ( rst_ni                                           ),
    .en_i   ( we_i[0]                                          ),
    .d_i    ( {a_gamma1,   a_gamma0,   b_gamma1,   b_gamma0}   ),
    .q_o    ( {a_gamma1_q, a_gamma0_q, b_gamma1_q, b_gamma0_q} )
  );

  logic [3:0] b_gamma10_prd2;
  aes_dom_dep_mul_gf2pn #(
    .NPower      ( 2           ),
    .Pipeline    ( PipelineMul ),
    .PreDomIndep ( 1'b0        )
  ) u_aes_dom_mul_gamma1_gamma0 (
    .clk_i  ( clk_i           ),
    .rst_ni ( rst_ni          ),
    .we_i   ( we_i[0]         ),
    .a_x    ( a_gamma1        ), // Share a of x
    .a_y    ( a_gamma0        ), // Share a of y
    .b_x    ( b_gamma1        ), // Share b of x
    .b_y    ( b_gamma0        ), // Share b of y
    .a_x_q  ( a_gamma1_q      ), // Share a of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .a_y_q  ( a_gamma0_q      ), // Share a of y, pipelined (for Pipeline=1)
    .b_x_q  ( b_gamma1_q      ), // Share b of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .b_y_q  ( b_gamma0_q      ), // Share b of y, pipelined (for Pipeline=1)
    .z_0    ( prd_2_i[1:0]    ), // Randomness for blinding
    .z_1    ( prd_2_i[3:2]    ), // Randomness for resharing
    .a_q    ( a_gamma1_gamma0 ), // Share a of q
    .b_q    ( b_gamma1_gamma0 ), // Share b of q
    .prd_o  ( b_gamma10_prd2  )  // Randomness for use in another S-Box instance
  );

  // Use intermediate results for generating PRD for Stage 3 of another S-Box instance.
  // Use one share only. Directly use output of flops updating with we_i[0].
  // b_gamma10_prd2 is based on b_gamma1_q, b_gamma0_q but XORed with prd_2_i, thus uniformly
  // distributed and independent of b_gamma1/0_q (See Lemma 1 in [2]).
  //
  // In Stage 3 of another S-Box instance, the MSBs and LSBs of the term below are used:
  // 1. as randomness in the DOM-dep multipliers u_aes_dom_mul_omega_gamma1/0, and
  // 2. to generate randomness for the DOM-indep multipliers u_aes_dom_mul_theta_y1/0 in Stage 4 of
  //    yet another S-Box instance, respectively.
  // Without interleaving b_gamma1/0_q as well as the upper and lower halves of b_gamma10_prd2 here,
  // a glitch on the write-enable signal on the input pipeline register of these DOM-indep
  // multipliers may result in undesirable SCA leakage.
  assign prd_2_o = {b_gamma1_q, b_gamma10_prd2[3:2], b_gamma0_q, b_gamma10_prd2[1:0]};

  /////////////
  // Stage 3 //
  /////////////

  // Formulas 14 and 15 in [2].
  logic [1:0] a_omega, b_omega;
  assign a_omega = aes_square_gf2p2(a_gamma1_gamma0 ^ a_gamma_ss_q);
  assign b_omega = aes_square_gf2p2(b_gamma1_gamma0 ^ b_gamma_ss_q);

  // Avoid aggressive synthesis optimizations.
  logic [1:0] a_omega_buf, b_omega_buf;
  prim_buf #(
    .Width ( 4 )
  ) u_prim_buf_ab_omega (
    .in_i  ( {a_omega,     b_omega}     ),
    .out_o ( {a_omega_buf, b_omega_buf} )
  );

  // Pipeline registers
  logic [1:0] a_gamma1_qq, a_gamma0_qq, b_gamma1_qq, b_gamma0_qq, a_omega_buf_q, b_omega_buf_q;
  if (PipelineMul == 1'b1) begin: gen_prim_flop_omega_gamma10
    // We instantiate the input pipeline registers for the DOM-dep multiplier outside of the
    // multiplier to enable sharing of pipeline registers where applicable.

    prim_flop_en #(
      .Width      ( 8  ),
      .ResetValue ( '0 )
    ) u_prim_flop_ab_gamma10_q (
      .clk_i  ( clk_i                                                ),
      .rst_ni ( rst_ni                                               ),
      .en_i   ( we_i[1]                                              ),
      .d_i    ( {a_gamma1_q,  a_gamma0_q,  b_gamma1_q,  b_gamma0_q}  ),
      .q_o    ( {a_gamma1_qq, a_gamma0_qq, b_gamma1_qq, b_gamma0_qq} )
    );

    // These inputs are used by both DOM-dep multipliers below.
    prim_flop_en #(
      .Width      ( 4  ),
      .ResetValue ( '0 )
    ) u_prim_flop_ab_omega_buf (
      .clk_i  ( clk_i                          ),
      .rst_ni ( rst_ni                         ),
      .en_i   ( we_i[1]                        ),
      .d_i    ( {a_omega_buf,   b_omega_buf}   ),
      .q_o    ( {a_omega_buf_q, b_omega_buf_q} )
    );

  end else begin : gen_no_prim_flop_ab_y10
    // When using un-pipelined multipliers, there is no need to insert additional registers.
    // We drive the corresponding inputs to 0 to make sure the functionality isn't correct in case
    // the pipeliend inputs are erroneously used.

    assign a_gamma1_qq = '0;
    assign a_gamma0_qq = '0;
    assign b_gamma1_qq = '0;
    assign b_gamma0_qq = '0;
    assign a_omega_buf_q = '0;
    assign b_omega_buf_q = '0;
  end

  // Formulas 16 and 17 in [2].
  logic [3:0] b_gamma1_omega_prd3;
  aes_dom_dep_mul_gf2pn #(
    .NPower      ( 2           ),
    .Pipeline    ( PipelineMul ),
    .PreDomIndep ( 1'b0        )
  ) u_aes_dom_mul_omega_gamma1 (
    .clk_i  ( clk_i               ),
    .rst_ni ( rst_ni              ),
    .we_i   ( we_i[1]             ),
    .a_x    ( a_gamma1_q          ), // Share a of x
    .a_y    ( a_omega_buf         ), // Share a of y
    .b_x    ( b_gamma1_q          ), // Share b of x
    .b_y    ( b_omega_buf         ), // Share b of y
    .a_x_q  ( a_gamma1_qq         ), // Share a of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .a_y_q  ( a_omega_buf_q       ), // Share a of y, pipelined (for Pipeline=1)
    .b_x_q  ( b_gamma1_qq         ), // Share b of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .b_y_q  ( b_omega_buf_q       ), // Share b of y, pipelined (for Pipeline=1)
    .z_0    ( prd_3_i[5:4]        ), // Randomness for blinding
    .z_1    ( prd_3_i[7:6]        ), // Randomness for resharing
    .a_q    ( a_gamma_inv[1:0]    ), // Share a of q
    .b_q    ( b_gamma_inv[1:0]    ), // Share b of q
    .prd_o  ( b_gamma1_omega_prd3 )  // Randomness for use in another S-Box instance
  );

  logic [3:0] b_gamma0_omega_prd3;
  aes_dom_dep_mul_gf2pn #(
    .NPower      ( 2           ),
    .Pipeline    ( PipelineMul ),
    .PreDomIndep ( 1'b0        )
  ) u_aes_dom_mul_omega_gamma0 (
    .clk_i  ( clk_i               ),
    .rst_ni ( rst_ni              ),
    .we_i   ( we_i[1]             ),
    .a_x    ( a_omega_buf         ), // Share a of x
    .a_y    ( a_gamma0_q          ), // Share a of y
    .b_x    ( b_omega_buf         ), // Share b of x
    .b_y    ( b_gamma0_q          ), // Share b of y
    .a_x_q  ( a_omega_buf_q       ), // Share a of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .a_y_q  ( a_gamma0_qq         ), // Share a of y, pipelined (for Pipeline=1)
    .b_x_q  ( b_omega_buf_q       ), // Share b of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .b_y_q  ( b_gamma0_qq         ), // Share b of y, pipelined (for Pipeline=1)
    .z_0    ( prd_3_i[1:0]        ), // Randomness for blinding
    .z_1    ( prd_3_i[3:2]        ), // Randomness for resharing
    .a_q    ( a_gamma_inv[3:2]    ), // Share a of q
    .b_q    ( b_gamma_inv[3:2]    ), // Share b of q
    .prd_o  ( b_gamma0_omega_prd3 )  // Randomness for use in another S-Box instance
  );

  // Use intermediate results for generating PRD for Stage 4 of another S-Box instance.
  // Use one share only. Directly use output of flops updating with we_i[1].
  // b_gamma1/0_omega_prd3 are both based on b_omega but XORed with differend parts of prd_3_i,
  // thus uniformly distributed and independent of b_omega (see Lemma 1 in [2]).
  assign prd_3_o = {b_gamma1_omega_prd3, b_gamma0_omega_prd3};

endmodule

// Inverse in GF(2^8) using first-order domain-oriented masking and normal basis [y^16, y].
// See Fig. 6 in [1] and Formulas 3, 12, 18 and 19 in [2].
module aes_dom_inverse_gf2p8 #(
  parameter bit PipelineMul = 1'b1
) (
  input  logic        clk_i,
  input  logic        rst_ni,
  input  logic  [3:0] we_i,
  input  logic  [7:0] a_y,     // input data masked by b_y
  input  logic  [7:0] b_y,     // input mask
  input  prd_in_t     prd_i,   // pseudo-random data, e.g. for intermediate masks
  output logic  [7:0] a_y_inv, // output data masked by b_y_inv
  output logic  [7:0] b_y_inv, // output mask
  output prd_out_t    prd_o    // pseudo-random data, e.g. for use in another S-Box instance
);

  import aes_sbox_canright_pkg::*;

  /////////////
  // Stage 1 //
  /////////////
  // Formula 12 in [2].

  logic [3:0] a_y1, a_y0, b_y1, b_y0, a_y1_y0, b_y1_y0;
  assign a_y1 = a_y[7:4];
  assign a_y0 = a_y[3:0];
  assign b_y1 = b_y[7:4];
  assign b_y0 = b_y[3:0];

  logic [3:0] a_y_ss_d, b_y_ss_d;
  logic [3:0] a_y_ss_q, b_y_ss_q;
  assign a_y_ss_d = aes_square_scale_gf2p4_gf2p2(a_y1 ^ a_y0);
  assign b_y_ss_d = aes_square_scale_gf2p4_gf2p2(b_y1 ^ b_y0);
  prim_flop_en #(
    .Width      ( 8  ),
    .ResetValue ( '0 )
  ) u_prim_flop_ab_y_ss (
    .clk_i  ( clk_i                ),
    .rst_ni ( rst_ni               ),
    .en_i   ( we_i[0]              ),
    .d_i    ( {a_y_ss_d, b_y_ss_d} ),
    .q_o    ( {a_y_ss_q, b_y_ss_q} )
  );

  logic [3:0] a_y1_q, a_y0_q, b_y1_q, b_y0_q;
  if (PipelineMul == 1'b1) begin: gen_prim_flop_ab_y10
    // We instantiate the input pipeline registers for the DOM-dep multiplier outside of the
    // multiplier to enable sharing of pipeline registers where applicable.

    prim_flop_en #(
      .Width      ( 16  ),
      .ResetValue ( '0  )
    ) u_prim_flop_ab_y10 (
      .clk_i  ( clk_i                            ),
      .rst_ni ( rst_ni                           ),
      .en_i   ( we_i[0]                          ),
      .d_i    ( {a_y1,   a_y0,   b_y1,   b_y0}   ),
      .q_o    ( {a_y1_q, a_y0_q, b_y1_q, b_y0_q} )
    );

  end else begin : gen_no_prim_flop_ab_y10
    // When using un-pipelined multipliers, there is no need to insert additional registers.
    // We drive the corresponding inputs to 0 to make sure the functionality isn't correct in case
    // the pipeliend inputs are erroneously used.

    assign a_y1_q = '0;
    assign a_y0_q = '0;
    assign b_y1_q = '0;
    assign b_y0_q = '0;
  end

  logic [7:0] b_y10_prd1;
  aes_dom_dep_mul_gf2pn #(
    .NPower      ( 4           ),
    .Pipeline    ( PipelineMul ),
    .PreDomIndep ( 1'b0        )
  ) u_aes_dom_mul_y1_y0 (
    .clk_i  ( clk_i            ),
    .rst_ni ( rst_ni           ),
    .we_i   ( we_i[0]          ),
    .a_x    ( a_y1             ), // Share a of x
    .a_y    ( a_y0             ), // Share a of y
    .b_x    ( b_y1             ), // Share b of x
    .b_y    ( b_y0             ), // Share b of y
    .a_x_q  ( a_y1_q           ), // Share a of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .a_y_q  ( a_y0_q           ), // Share a of y, pipelined (for Pipeline=1)
    .b_x_q  ( b_y1_q           ), // Share b of x, pipelined (for Pipeline=1 or PreDomIndep=1)
    .b_y_q  ( b_y0_q           ), // Share b of y, pipelined (for Pipeline=1)
    .z_0    ( prd_i.prd_1[3:0] ), // Randomness for blinding
    .z_1    ( prd_i.prd_1[7:4] ), // Randomness for resharing
    .a_q    ( a_y1_y0          ), // Share a of q
    .b_q    ( b_y1_y0          ), // Share b of q
    .prd_o  ( b_y10_prd1       )  // Randomness for use in another S-Box instance
  );

  logic [3:0] a_gamma, b_gamma;
  assign a_gamma = a_y_ss_q ^ a_y1_y0;
  assign b_gamma = b_y_ss_q ^ b_y1_y0;

  // Avoid aggressive synthesis optimizations.
  logic [3:0] a_gamma_buf, b_gamma_buf;
  prim_buf #(
    .Width ( 8 )
  ) u_prim_buf_ab_gamma (
    .in_i  ( {a_gamma,     b_gamma}     ),
    .out_o ( {a_gamma_buf, b_gamma_buf} )
  );

  // Use intermediate results for generating PRD for Stage 2 of another S-Box instance.
  // Use one share only. Directly use output of flops updating with we_i[0].
  // b_y10_prd1 is based on b_y and XORed with prd_1. We just use the lower part involving a
  // non-linear element.
  assign prd_o.prd_1 = b_y10_prd1[3:0];
  logic [3:0] unused_prd;
  assign unused_prd  = b_y10_prd1[7:4];

  ////////////////////
  // Stages 2 and 3 //
  ////////////////////

  logic [3:0] a_theta, b_theta;

  // a_gamma is masked by b_gamma, a_gamma_inv is masked by b_gamma_inv.
  aes_dom_inverse_gf2p4 #(
    .PipelineMul ( PipelineMul )
  ) u_aes_dom_inverse_gf2p4 (
    .clk_i       ( clk_i       ),
    .rst_ni      ( rst_ni      ),
    .we_i        ( we_i[2:1]   ),
    .a_gamma     ( a_gamma_buf ),
    .b_gamma     ( b_gamma_buf ),
    .prd_2_i     ( prd_i.prd_2 ),
    .prd_3_i     ( prd_i.prd_3 ),
    .a_gamma_inv ( a_theta     ),
    .b_gamma_inv ( b_theta     ),
    .prd_2_o     ( prd_o.prd_2 ),
    .prd_3_o     ( prd_o.prd_3 )
  );

  /////////////
  // Stage 4 //
  /////////////
  // Formulas 18 and 19 in [2].

  logic [3:0] a_y1_qqq, a_y0_qqq, b_y1_qqq, b_y0_qqq;
  prim_flop_en #(
    .Width      ( 16 ),
    .ResetValue ( '0 )
  ) u_prim_flop_ab_y10_qqq (
    .clk_i  ( clk_i                                    ),
    .rst_ni ( rst_ni                                   ),
    .en_i   ( we_i[2]                                  ),
    .d_i    ( {a_y1,     a_y0,     b_y1,     b_y0}     ),
    .q_o    ( {a_y1_qqq, a_y0_qqq, b_y1_qqq, b_y0_qqq} )
  );

  aes_dom_indep_mul_gf2pn #(
    .NPower   ( 4           ),
    .Pipeline ( PipelineMul )
  ) u_aes_dom_mul_theta_y1 (
    .clk_i  ( clk_i            ),
    .rst_ni ( rst_ni           ),
    .we_i   ( we_i[3]          ),
    .a_x    ( a_y1_qqq         ), // Share a of x
    .a_y    ( a_theta          ), // Share a of y
    .b_x    ( b_y1_qqq         ), // Share b of x
    .b_y    ( b_theta          ), // Share b of y
    .z_0    ( prd_i.prd_4[7:4] ), // Randomness for resharing
    .a_q    ( a_y_inv[3:0]     ), // Share a of q
    .b_q    ( b_y_inv[3:0]     )  // Share b of q
  );

  aes_dom_indep_mul_gf2pn #(
    .NPower   ( 4           ),
    .Pipeline ( PipelineMul )
  ) u_aes_dom_mul_theta_y0 (
    .clk_i  ( clk_i            ),
    .rst_ni ( rst_ni           ),
    .we_i   ( we_i[3]          ),
    .a_x    ( a_theta          ), // Share a of x
    .a_y    ( a_y0_qqq         ), // Share a of y
    .b_x    ( b_theta          ), // Share b of x
    .b_y    ( b_y0_qqq         ), // Share b of y
    .z_0    ( prd_i.prd_4[3:0] ), // Randomness for resharing
    .a_q    ( a_y_inv[7:4]     ), // Share a of q
    .b_q    ( b_y_inv[7:4]     )  // Share b of q
  );

endmodule

// SEC_CM: KEY.MASKING
module aes_sbox_dom
#(
  parameter bit PipelineMul = 1'b1
) (
  input  logic              clk_i,
  input  logic              rst_ni,
  input  logic              en_i,
  input  logic              prd_we_i,
  output logic              out_req_o,
  input  logic              out_ack_i,
  input  aes_pkg::ciph_op_e op_i,
  input  logic        [7:0] data_i, // masked, the actual input data is data_i ^ mask_i
  input  logic        [7:0] mask_i, // input mask
  input  logic       [27:0] prd_i,  // pseudo-random data for remasking, in total we need 28 bits
                                    // of PRD per evaluation, but at most 8 bits per cycle
  output logic        [7:0] data_o, // masked, the actual output data is data_o ^ mask_o
  output logic        [7:0] mask_o, // output mask
  output logic       [19:0] prd_o   // PRD for usage in Stages 2 - 4 of other S-Box instances
);

  import aes_pkg::*;
  import aes_sbox_canright_pkg::*;

  logic [7:0] in_data_basis_x, out_data_basis_x;
  logic [7:0] in_mask_basis_x, out_mask_basis_x;
  logic [3:0] we;
  logic [7:0] prd1_d, prd1_q;
  prd_in_t    in_prd;
  prd_out_t   out_prd;

  // Convert data to normal basis X.
  assign in_data_basis_x = (op_i == CIPH_FWD) ? aes_mvm(data_i, A2X)         :
                           (op_i == CIPH_INV) ? aes_mvm(data_i ^ 8'h63, S2X) :
                                                aes_mvm(data_i, A2X);

  // Convert mask to normal basis X.
  // The addition of constant 8'h63 prior to the affine transformation is skipped.
  assign in_mask_basis_x = (op_i == CIPH_FWD) ? aes_mvm(mask_i, A2X) :
                           (op_i == CIPH_INV) ? aes_mvm(mask_i, S2X) :
                                                aes_mvm(mask_i, A2X);

  // Do the inversion in normal basis X.
  aes_dom_inverse_gf2p8 #(
    .PipelineMul ( PipelineMul )
  ) u_aes_dom_inverse_gf2p8 (
    .clk_i   ( clk_i            ),
    .rst_ni  ( rst_ni           ),
    .we_i    ( we               ),
    .a_y     ( in_data_basis_x  ), // input
    .b_y     ( in_mask_basis_x  ), // input
    .prd_i   ( in_prd           ), // input
    .a_y_inv ( out_data_basis_x ), // output
    .b_y_inv ( out_mask_basis_x ), // output
    .prd_o   ( out_prd          )  // output
  );

  // Convert data to basis S or A.
  assign data_o = (op_i == CIPH_FWD) ? (aes_mvm(out_data_basis_x, X2S) ^ 8'h63) :
                  (op_i == CIPH_INV) ? (aes_mvm(out_data_basis_x, X2A))         :
                                       (aes_mvm(out_data_basis_x, X2S) ^ 8'h63);

  // Convert mask to basis S or A.
  // The addition of constant 8'h63 following the affine transformation is skipped.
  assign mask_o = (op_i == CIPH_FWD) ? aes_mvm(out_mask_basis_x, X2S) :
                  (op_i == CIPH_INV) ? aes_mvm(out_mask_basis_x, X2A) :
                                       aes_mvm(out_mask_basis_x, X2S);

  // Counter register
  logic [2:0] count_d, count_q;
  assign count_d = (out_req_o && out_ack_i) ? '0             :
                   out_req_o                ? count_q        :
                   en_i                     ? count_q + 3'd1 : count_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_count
    if (!rst_ni) begin
      count_q <= '0;
    end else begin
      count_q <= count_d;
    end
  end
  assign out_req_o = en_i & count_q == 3'd4;

  // Write enable signals for internal registers
  assign we[0] = en_i & count_q == 3'd0;
  assign we[1] = en_i & count_q == 3'd1;
  assign we[2] = en_i & count_q == 3'd2;
  assign we[3] = en_i & count_q == 3'd3;

  // Buffer and forward PRD for the individual stages. We get 8 bits from the PRNG for usage in the
  // first cycle. Stages 2, 3 and 4 are driven by other S-Box instances.
  assign prd1_d = prd_we_i ? prd_i[7:0] : prd1_q;
  prim_flop #(
    .Width      ( 8  ),
    .ResetValue ( '0 )
  ) u_prim_flop_prd1_q (
    .clk_i  ( clk_i  ),
    .rst_ni ( rst_ni ),
    .d_i    ( prd1_d ),
    .q_o    ( prd1_q )
  );
  assign in_prd = '{prd_1: prd1_q,
                    prd_2: prd_i[11:8],
                    prd_3: prd_i[19:12],
                    prd_4: prd_i[27:20]};
  assign prd_o = {out_prd.prd_3, out_prd.prd_2, out_prd.prd_1};

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES ShiftRows

module aes_shift_rows (
  input  aes_pkg::ciph_op_e    op_i,
  input  logic [3:0][3:0][7:0] data_i,
  output logic [3:0][3:0][7:0] data_o
);

  import aes_pkg::*;

  // Row 0 is left untouched
  assign data_o[0] = data_i[0];

  // Row 2 does not depend on op_i
  assign data_o[2] = aes_circ_byte_shift(data_i[2], 2'h2);

  // Row 1
  assign data_o[1] = (op_i == CIPH_FWD) ? aes_circ_byte_shift(data_i[1], 2'h3) :
                     (op_i == CIPH_INV) ? aes_circ_byte_shift(data_i[1], 2'h1) :
                                          aes_circ_byte_shift(data_i[1], 2'h3);

  // Row 3
  assign data_o[3] = (op_i == CIPH_FWD) ? aes_circ_byte_shift(data_i[3], 2'h1) :
                     (op_i == CIPH_INV) ? aes_circ_byte_shift(data_i[3], 2'h3) :
                                          aes_circ_byte_shift(data_i[3], 2'h1);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES MixColumns

module aes_mix_columns (
  input  aes_pkg::ciph_op_e    op_i,
  input  logic [3:0][3:0][7:0] data_i,
  output logic [3:0][3:0][7:0] data_o
);

  import aes_pkg::*;

  // Transpose to operate on columns
  logic [3:0][3:0][7:0] data_i_transposed;
  logic [3:0][3:0][7:0] data_o_transposed;

  assign data_i_transposed = aes_transpose(data_i);

  // Individually mix columns
  for (genvar i = 0; i < 4; i++) begin : gen_mix_column
    aes_mix_single_column u_aes_mix_column_i (
      .op_i   ( op_i                 ),
      .data_i ( data_i_transposed[i] ),
      .data_o ( data_o_transposed[i] )
    );
  end

  assign data_o = aes_transpose(data_o_transposed);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES MixColumns for one single column of the state matrix
//
// For details, see Equations 4-7 of:
// Satoh et al., "A Compact Rijndael Hardware Architecture with S-Box Optimization"

module aes_mix_single_column (
  input  aes_pkg::ciph_op_e op_i,
  input  logic [3:0][7:0]   data_i,
  output logic [3:0][7:0]   data_o
);

  import aes_pkg::*;

  logic [3:0][7:0] x;
  logic [1:0][7:0] y;
  logic [1:0][7:0] z;

  logic [3:0][7:0] x_mul2;
  logic [1:0][7:0] y_pre_mul4;
  logic      [7:0] y2, y2_pre_mul2;

  logic [1:0][7:0] z_muxed;

  // Drive x
  assign x[0] = data_i[0] ^ data_i[3];
  assign x[1] = data_i[3] ^ data_i[2];
  assign x[2] = data_i[2] ^ data_i[1];
  assign x[3] = data_i[1] ^ data_i[0];

  // Mul2(x)
  for (genvar i = 0; i < 4; i++) begin : gen_x_mul2
    assign x_mul2[i] = aes_mul2(x[i]);
  end

  // Drive y_pre_mul4
  assign y_pre_mul4[0] = data_i[3] ^ data_i[1];
  assign y_pre_mul4[1] = data_i[2] ^ data_i[0];

  // Mul4(y_pre_mul4)
  for (genvar i = 0; i < 2; i++) begin : gen_mul4
    assign y[i] = aes_mul4(y_pre_mul4[i]);
  end

  // Drive y2_pre_mul2
  assign y2_pre_mul2 = y[0] ^ y[1];

  // Mul2(y)
  assign y2 = aes_mul2(y2_pre_mul2);

  // Drive z
  assign z[0] = y2 ^ y[0];
  assign z[1] = y2 ^ y[1];

  // Mux z
  assign z_muxed[0] = (op_i == CIPH_FWD) ? 8'b0 :
                      (op_i == CIPH_INV) ? z[0] : 8'b0;
  assign z_muxed[1] = (op_i == CIPH_FWD) ? 8'b0 :
                      (op_i == CIPH_INV) ? z[1] : 8'b0;

  // Drive outputs
  assign data_o[0] = data_i[1] ^ x_mul2[3] ^ x[1] ^ z_muxed[1];
  assign data_o[1] = data_i[0] ^ x_mul2[2] ^ x[1] ^ z_muxed[0];
  assign data_o[2] = data_i[3] ^ x_mul2[1] ^ x[3] ^ z_muxed[1];
  assign data_o[3] = data_i[2] ^ x_mul2[0] ^ x[3] ^ z_muxed[0];

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES KeyExpand

`include "prim_assert.sv"

module aes_key_expand import aes_pkg::*;
#(
  parameter bit         AES192Enable = 1,
  parameter bit         SecMasking   = 0,
  parameter sbox_impl_e SecSBoxImpl  = SBoxImplLut,

  localparam int        NumShares    = SecMasking ? 2 : 1 // derived parameter
) (
  input  logic                   clk_i,
  input  logic                   rst_ni,
  input  logic                   cfg_valid_i,
  input  ciph_op_e               op_i,
  input  sp2v_e                  en_i,
  input  logic                   prd_we_i,
  output sp2v_e                  out_req_o,
  input  sp2v_e                  out_ack_i,
  input  logic                   clear_i,
  input  logic             [3:0] round_i,
  input  key_len_e               key_len_i,
  input  logic       [7:0][31:0] key_i [NumShares],
  output logic       [7:0][31:0] key_o [NumShares],
  input  logic [WidthPRDKey-1:0] prd_i,
  output logic                   err_o
);

  sp2v_e            en;
  logic             en_err;
  sp2v_e            out_ack;
  logic             out_ack_err;

  logic       [7:0] rcon_d, rcon_q;
  logic             rcon_we;
  logic             use_rcon;

  logic       [3:0] rnd;
  logic       [3:0] rnd_type;

  logic      [31:0] spec_in_128 [NumShares];
  logic      [31:0] spec_in_192 [NumShares];
  logic      [31:0] rot_word_in [NumShares];
  logic      [31:0] rot_word_out [NumShares];
  logic             use_rot_word;
  logic             prd_we, prd_we_force, prd_we_inhibit;
  logic      [31:0] sub_word_in, sub_word_out;
  logic       [3:0] sub_word_out_req;
  logic      [31:0] sw_in_mask, sw_out_mask;
  logic       [7:0] rcon_add_in, rcon_add_out;
  logic      [31:0] rcon_added;

  logic      [31:0] irregular [NumShares];
  logic [7:0][31:0] regular [NumShares];

  // cfg_valid_i is used for gating assertions only.
  logic                     unused_cfg_valid;
  assign unused_cfg_valid = cfg_valid_i;

  // Get a shorter reference.
  assign rnd = round_i;

  // For AES-192, there are four different types of rounds.
  always_comb begin : get_rnd_type
    if (AES192Enable) begin
      rnd_type[0] = (rnd == 0);
      rnd_type[1] = (rnd == 1 || rnd == 4 || rnd == 7 || rnd == 10);
      rnd_type[2] = (rnd == 2 || rnd == 5 || rnd == 8 || rnd == 11);
      rnd_type[3] = (rnd == 3 || rnd == 6 || rnd == 9 || rnd == 12);
    end else begin
      rnd_type = '0;
    end
  end

  //////////////////////////////////////////////////////
  // Irregular part involving Rcon, RotWord & SubWord //
  //////////////////////////////////////////////////////

  // Depending on key length and round, RotWord may not be used.
  assign use_rot_word = (key_len_i == AES_256 && rnd[0] == 1'b0) ? 1'b0 : 1'b1;

  // Depending on operation, key length and round, Rcon may not be used thus must not be updated.
  always_comb begin : rcon_usage
    use_rcon = 1'b1;

    if (AES192Enable) begin
      if (key_len_i == AES_192 &&
          ((op_i == CIPH_FWD &&  rnd_type[1]) ||
           (op_i == CIPH_INV && (rnd_type[0] || rnd_type[3])))) begin
        use_rcon = 1'b0;
      end
    end

    if (key_len_i == AES_256 && rnd[0] == 1'b0) begin
      use_rcon = 1'b0;
    end
  end

  // Generate Rcon
  always_comb begin : rcon_update
    rcon_d = rcon_q;

    if (clear_i) begin
      rcon_d = (op_i == CIPH_FWD)                            ? 8'h01 :
              ((op_i == CIPH_INV) && (key_len_i == AES_128)) ? 8'h36 :
              ((op_i == CIPH_INV) && (key_len_i == AES_192)) ? 8'h80 :
              ((op_i == CIPH_INV) && (key_len_i == AES_256)) ? 8'h40 : 8'h01;
    end else begin
      rcon_d = (op_i == CIPH_FWD) ? aes_mul2(rcon_q) :
               (op_i == CIPH_INV) ? aes_div2(rcon_q) : 8'h01;
    end
  end

  // Advance.
  assign rcon_we = clear_i | use_rcon &
      (en == SP2V_HIGH) & (out_req_o == SP2V_HIGH) & (out_ack == SP2V_HIGH);

  // Rcon register
  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_rcon
    if (!rst_ni) begin
      rcon_q <= '0;
    end else if (rcon_we) begin
      rcon_q <= rcon_d;
    end
  end

  for (genvar s = 0; s < NumShares; s++) begin : gen_shares_rot_word_out
    // Special input, equivalent to key_o[3] in the used cases
    assign spec_in_128[s] = key_i[s][3] ^ key_i[s][2];
    assign spec_in_192[s] = AES192Enable ? key_i[s][5] ^ key_i[s][1] ^ key_i[s][0] : '0;

    // Select input
    always_comb begin : rot_word_in_mux
      unique case (key_len_i)

        /////////////
        // AES-128 //
        /////////////
        AES_128: begin
          unique case (op_i)
            CIPH_FWD: rot_word_in[s] = key_i[s][3];
            CIPH_INV: rot_word_in[s] = spec_in_128[s];
            default:  rot_word_in[s] = key_i[s][3];
          endcase
        end

        /////////////
        // AES-192 //
        /////////////
        AES_192: begin
          if (AES192Enable) begin
            unique case (op_i)
              CIPH_FWD: begin
                rot_word_in[s] = rnd_type[0] ? key_i[s][5]    :
                                 rnd_type[2] ? key_i[s][5]    :
                                 rnd_type[3] ? spec_in_192[s] : key_i[s][3];
              end
              CIPH_INV: begin
                rot_word_in[s] = rnd_type[1] ? key_i[s][3] :
                                 rnd_type[2] ? key_i[s][1] : key_i[s][3];
              end
              default: rot_word_in[s] = key_i[s][3];
            endcase
          end else begin
            rot_word_in[s] = key_i[s][3];
          end
        end

        /////////////
        // AES-256 //
        /////////////
        AES_256: begin
          unique case (op_i)
            CIPH_FWD: rot_word_in[s] = key_i[s][7];
            CIPH_INV: rot_word_in[s] = key_i[s][3];
            default:  rot_word_in[s] = key_i[s][7];
          endcase
        end

        default: rot_word_in[s] = key_i[s][3];
      endcase
    end

    // RotWord: cyclic byte shift
    assign rot_word_out[s] = aes_circ_byte_shift(rot_word_in[s], 2'h3);
  end

  // Mux input for SubWord
  assign sub_word_in = use_rot_word ? rot_word_out[0] : rot_word_in[0];

  // Masking
  if (!SecMasking) begin : gen_no_sw_in_mask
    // The mask share is ignored anyway, it can be 0.
    assign sw_in_mask  = '0;

    // Tie-off unused signals.
    logic [31:0] unused_sw_out_mask;
    assign unused_sw_out_mask = sw_out_mask;

  end else begin : gen_sw_in_mask
    // The input mask is the mask share of rot_word_in/out.
    assign sw_in_mask = use_rot_word ? rot_word_out[1] : rot_word_in[1];
  end

  // SubWord - individually substitute bytes.
  // Every DOM S-Box instance consumes 28 bits of randomness but itself produces 20 bits for use in
  // another S-Box instance. For other S-Box implementations, only the bits corresponding to prd_i
  // are used. Other bits are ignored and tied to 0.
  logic [3:0][WidthPRDSBox+19:0] in_prd;
  logic [3:0]             [19:0] out_prd;

  // Make sure that whenever the data/mask inputs of the S-Boxes update, the internally buffered
  // PRD is updated in sync. There are two special cases we need to handle here:
  // - For AES-256, the initial round is short (no round key computation). But the data/mask inputs
  //   are updated either way. Thus, we need to force a PRD update as well.
  // - For AES-192 in FWD mode, the data/mask inputs aren't updated in Round 1, 4, 7 and 10. Thus,
  //   we need to inhibit PRD updates triggred at the end of Round 0, 3, 6 and 9.
  assign prd_we_force = (key_len_i == AES_256) & (rnd == 0);
  assign prd_we_inhibit = (key_len_i == AES_192) & (op_i == CIPH_FWD) &
      (rnd == 0 || rnd == 3 || rnd == 6 || rnd == 9);
  assign prd_we = (prd_we_i & ~prd_we_inhibit) | prd_we_force;

  for (genvar i = 0; i < 4; i++) begin : gen_sbox
    // Rotate the randomness produced by the S-Boxes. The LSBs are taken from the masking PRNG
    // (prd_i) whereas the MSBs are produced by the other S-Box instances.
    assign in_prd[i] = {out_prd[aes_rot_int(i,4)], prd_i[WidthPRDSBox*i +: WidthPRDSBox]};

    aes_sbox #(
      .SecSBoxImpl ( SecSBoxImpl )
    ) u_aes_sbox_i (
      .clk_i     ( clk_i                  ),
      .rst_ni    ( rst_ni                 ),
      .en_i      ( en == SP2V_HIGH        ),
      .prd_we_i  ( prd_we                 ),
      .out_req_o ( sub_word_out_req[i]    ),
      .out_ack_i ( out_ack == SP2V_HIGH   ),
      .op_i      ( CIPH_FWD               ),
      .data_i    ( sub_word_in[8*i +: 8]  ),
      .mask_i    ( sw_in_mask[8*i +: 8]   ),
      .prd_i     ( in_prd[i]              ),
      .data_o    ( sub_word_out[8*i +: 8] ),
      .mask_o    ( sw_out_mask[8*i +: 8]  ),
      .prd_o     ( out_prd[i]             )
    );
  end

  // Add Rcon
  assign rcon_add_in  = sub_word_out[7:0];
  assign rcon_add_out = rcon_add_in ^ rcon_q;
  assign rcon_added   = {sub_word_out[31:8], rcon_add_out};

  // Mux output coming from Rcon & SubWord
  for (genvar s = 0; s < NumShares; s++) begin : gen_shares_irregular
    if (s == 0) begin : gen_irregular_rcon
      // The (masked) key share
      assign irregular[s] = use_rcon ? rcon_added : sub_word_out;
    end else begin : gen_irregular_no_rcon
      // The mask share
      assign irregular[s] = sw_out_mask;
    end
  end

  ///////////////////////////
  // The more regular part //
  ///////////////////////////

  // To reduce muxing resources, we re-use existing
  // connections for unused words and default cases.
  for (genvar s = 0; s < NumShares; s++) begin : gen_shares_regular
    always_comb begin : drive_regular
      unique case (key_len_i)

        /////////////
        // AES-128 //
        /////////////
        AES_128: begin
          // key_o[7:4] not used
          regular[s][7:4] = key_i[s][3:0];

          regular[s][0] = irregular[s] ^ key_i[s][0];
          unique case (op_i)
            CIPH_FWD: begin
              for (int i = 1; i < 4; i++) begin
                regular[s][i] = regular[s][i-1] ^ key_i[s][i];
              end
            end

            CIPH_INV: begin
              for (int i = 1; i < 4; i++) begin
                regular[s][i] = key_i[s][i-1] ^ key_i[s][i];
              end
            end

            default: regular[s] = {key_i[s][3:0], key_i[s][7:4]};
          endcase
        end

        /////////////
        // AES-192 //
        /////////////
        AES_192: begin
          // key_o[7:6] not used
          regular[s][7:6] = key_i[s][3:2];

          if (AES192Enable) begin
            unique case (op_i)
              CIPH_FWD: begin
                if (rnd_type[0]) begin
                  // Shift down four upper most words
                  regular[s][3:0] = key_i[s][5:2];
                  // Generate Words 6 and 7
                  regular[s][4]   = irregular[s]  ^ key_i[s][0];
                  regular[s][5]   = regular[s][4] ^ key_i[s][1];
                end else begin
                  // Shift down two upper most words
                  regular[s][1:0] = key_i[s][5:4];
                  // Generate new upper four words
                  for (int i = 0; i < 4; i++) begin
                    if ((i == 0 && rnd_type[2]) ||
                        (i == 2 && rnd_type[3])) begin
                      regular[s][i+2] = irregular[s]    ^ key_i[s][i];
                    end else begin
                      regular[s][i+2] = regular[s][i+1] ^ key_i[s][i];
                    end
                  end
                end // rnd_type[0]
              end

              CIPH_INV: begin
                if (rnd_type[0]) begin
                  // Shift up four lowest words
                  regular[s][5:2] = key_i[s][3:0];
                  // Generate Word 44 and 45
                  for (int i = 0; i < 2; i++) begin
                    regular[s][i] = key_i[s][3+i] ^ key_i[s][3+i+1];
                  end
                end else begin
                  // Shift up two lowest words
                  regular[s][5:4] = key_i[s][1:0];
                  // Generate new lower four words
                  for (int i = 0; i < 4; i++) begin
                    if ((i == 2 && rnd_type[1]) ||
                        (i == 0 && rnd_type[2])) begin
                      regular[s][i] = irregular[s]  ^ key_i[s][i+2];
                    end else begin
                      regular[s][i] = key_i[s][i+1] ^ key_i[s][i+2];
                    end
                  end
                end // rnd_type[0]
              end

              default: regular[s] = {key_i[s][3:0], key_i[s][7:4]};
            endcase

          end else begin
            regular[s] = {key_i[s][3:0], key_i[s][7:4]};
          end // AES192Enable
        end

        /////////////
        // AES-256 //
        /////////////
        AES_256: begin
          unique case (op_i)
            CIPH_FWD: begin
              if (rnd == 0) begin
                // Round 0: Nothing to be done
                // The Full Key registers are not updated
                regular[s] = {key_i[s][3:0], key_i[s][7:4]};
              end else begin
                // Shift down old upper half
                regular[s][3:0] = key_i[s][7:4];
                // Generate new upper half
                regular[s][4]   = irregular[s] ^ key_i[s][0];
                for (int i = 1; i < 4; i++) begin
                  regular[s][i+4] = regular[s][i+4-1] ^ key_i[s][i];
                end
              end // rnd == 0
            end

            CIPH_INV: begin
              if (rnd == 0) begin
                // Round 0: Nothing to be done
                // The Full Key registers are not updated
                regular[s] = {key_i[s][3:0], key_i[s][7:4]};
              end else begin
                // Shift up old lower half
                regular[s][7:4] = key_i[s][3:0];
                // Generate new lower half
                regular[s][0]   = irregular[s] ^ key_i[s][4];
                for (int i = 0; i < 3; i++) begin
                  regular[s][i+1] = key_i[s][4+i] ^ key_i[s][4+i+1];
                end
              end // rnd == 0
            end

            default: regular[s] = {key_i[s][3:0], key_i[s][7:4]};
          endcase
        end

        default: regular[s] = {key_i[s][3:0], key_i[s][7:4]};
      endcase // key_len_i
    end // drive_regular
  end // gen_shares_regular

  // Drive output
  assign key_o     = regular;
  assign out_req_o = &sub_word_out_req ? SP2V_HIGH : SP2V_LOW;

  //////////////////////////////
  // Sparsely Encoded Signals //
  //////////////////////////////

  logic [Sp2VWidth-1:0] en_raw;
  aes_sel_buf_chk #(
    .Num      ( Sp2VNum   ),
    .Width    ( Sp2VWidth ),
    .EnSecBuf ( 1'b1      )
  ) u_aes_key_expand_en_buf_chk (
    .clk_i  ( clk_i  ),
    .rst_ni ( rst_ni ),
    .sel_i  ( en_i   ),
    .sel_o  ( en_raw ),
    .err_o  ( en_err )
  );
  assign en = sp2v_e'(en_raw);

  logic [Sp2VWidth-1:0] out_ack_raw;
  aes_sel_buf_chk #(
    .Num      ( Sp2VNum   ),
    .Width    ( Sp2VWidth ),
    .EnSecBuf ( 1'b1      )
  ) u_aes_key_expand_out_ack_buf_chk (
    .clk_i  ( clk_i       ),
    .rst_ni ( rst_ni      ),
    .sel_i  ( out_ack_i   ),
    .sel_o  ( out_ack_raw ),
    .err_o  ( out_ack_err )
  );
  assign out_ack = sp2v_e'(out_ack_raw);

  // Collect encoding errors.
  assign err_o = en_err | out_ack_err;

  ////////////////
  // Assertions //
  ////////////////

  // Create a lint error to reduce the risk of accidentally disabling the masking.
  `ASSERT_STATIC_LINT_ERROR(AesKeyExpandSecMaskingNonDefault, SecMasking == 1)

  // Cipher core masking requires a masked SBox and vice versa.
  `ASSERT_INIT(AesMaskedCoreAndSBox,
      (SecMasking &&
      (SecSBoxImpl == SBoxImplCanrightMasked ||
       SecSBoxImpl == SBoxImplCanrightMaskedNoreuse ||
       SecSBoxImpl == SBoxImplDom)) ||
      (!SecMasking &&
      (SecSBoxImpl == SBoxImplLut ||
       SecSBoxImpl == SBoxImplCanright)))

  // Selectors must be known/valid
  `ASSERT(AesCiphOpValid, cfg_valid_i |-> op_i inside {
      CIPH_FWD,
      CIPH_INV
      })
  `ASSERT(AesKeyLenValid, cfg_valid_i |-> key_len_i inside {
      AES_128,
      AES_192,
      AES_256
      })

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES low-bandwidth pseudo-random number generator for register clearing
//
// This module uses an LFSR followed by an aligned permutation, a non-linear layer (PRINCE S-Boxes)
// and another permutation to generate pseudo-random data for the AES module for clearing
// registers (secure wipe). The LFSR can be reseeded using an external interface.

`include "prim_assert.sv"

module aes_prng_clearing import aes_pkg::*;
#(
  parameter int unsigned Width                = 64, // At the moment we just support a width of 64.
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,
  parameter bit          SecSkipPRNGReseeding = 0,  // The current SCA setup doesn't provide
                                                    // sufficient resources to implement the
                                                    // infrastructure required for PRNG reseeding.
                                                    // To enable SCA resistance evaluations, we
                                                    // need to skip reseeding requests.
  parameter clearing_lfsr_seed_t RndCnstLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstSharePerm = RndCnstClearingSharePermDefault
) (
  input  logic                    clk_i,
  input  logic                    rst_ni,

  // Connections to AES internals, PRNG consumers
  input  logic                    data_req_i,
  output logic                    data_ack_o,
  output logic        [Width-1:0] data_o [NumSharesKey],
  input  logic                    reseed_req_i,
  output logic                    reseed_ack_o,

  // Connections to outer world, LFSR re-seed
  output logic                    entropy_req_o,
  input  logic                    entropy_ack_i,
  input  logic [EntropyWidth-1:0] entropy_i
);

  logic             seed_valid;
  logic             seed_en;
  logic [Width-1:0] seed;
  logic             lfsr_en;
  logic [Width-1:0] lfsr_state;

  // In the current SCA setup, we don't have sufficient resources to implement the infrastructure
  // required for PRNG reseeding (CSRNG, EDN, etc.). Therefore, we skip any reseeding requests if
  // the SecSkipPRNGReseeding parameter is set. Performing the reseeding without proper entropy
  // provided from CSRNG would result in quickly repeating, fully deterministic PRNG output,
  // which prevents meaningful SCA resistance evaluations.

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(AesSecSkipPRNGReseedingNonDefault, SecSkipPRNGReseeding == 0)

  // LFSR control
  assign lfsr_en = data_req_i & data_ack_o;
  assign seed_en = SecSkipPRNGReseeding ? 1'b0 : seed_valid;

  // The data requests are fed from the LFSR, reseed requests have the highest priority.
  assign data_ack_o = reseed_req_i ? 1'b0 : data_req_i;

  // Width adaption for reseeding interface. We get EntropyWidth bits at a time.
  if (Width/2 == EntropyWidth) begin : gen_buffer
    // We buffer the first EntropyWidth bits.
    logic [EntropyWidth-1:0] buffer_d, buffer_q;
    logic                    buffer_valid_d, buffer_valid_q;

    // Stop requesting entropy once we have reseeded the LFSR.
    assign entropy_req_o = SecSkipPRNGReseeding ? 1'b0         : reseed_req_i;
    assign reseed_ack_o  = SecSkipPRNGReseeding ? reseed_req_i : seed_valid;

    // Buffer
    assign buffer_valid_d = entropy_req_o && entropy_ack_i ? ~buffer_valid_q : buffer_valid_q;

    // Only update the buffer upon receiving the first EntropyWidth bits.
    assign buffer_d = entropy_req_o && entropy_ack_i && !buffer_valid_q ? entropy_i : buffer_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin : reg_buffer
      if (!rst_ni) begin
        buffer_q       <= '0;
        buffer_valid_q <= 1'b0;
      end else begin
        buffer_q       <= buffer_d;
        buffer_valid_q <= buffer_valid_d;
      end
    end

    assign seed       = {buffer_q, entropy_i};
    assign seed_valid = buffer_valid_q & entropy_req_o & entropy_ack_i;

  end else begin : gen_packer
    // Upsizing of entropy input to correct width for LFSR reseeding.

    // Stop requesting entropy once the desired amount is available.
    assign entropy_req_o = SecSkipPRNGReseeding ? 1'b0         : reseed_req_i & ~seed_valid;
    assign reseed_ack_o  = SecSkipPRNGReseeding ? reseed_req_i : seed_valid;

    prim_packer_fifo #(
      .InW         ( EntropyWidth ),
      .OutW        ( Width        ),
      .ClearOnRead ( 1'b0         )
    ) u_prim_packer_fifo (
      .clk_i    ( clk_i         ),
      .rst_ni   ( rst_ni        ),
      .clr_i    ( 1'b0          ), // Not needed.
      .wvalid_i ( entropy_ack_i ),
      .wdata_i  ( entropy_i     ),
      .wready_o (               ), // Not needed, we're always ready to sink data at this point.
      .rvalid_o ( seed_valid    ),
      .rdata_o  ( seed          ),
      .rready_i ( 1'b1          ), // We're always ready to receive the packed output word.
      .depth_o  (               )  // Not needed.
    );
  end

  // LFSR instance
  prim_lfsr #(
    .LfsrType     ( "GAL_XOR"       ),
    .LfsrDw       ( Width           ),
    .StateOutDw   ( Width           ),
    .DefaultSeed  ( RndCnstLfsrSeed ),
    .StatePermEn  ( 1'b1            ),
    .StatePerm    ( RndCnstLfsrPerm ),
    .NonLinearOut ( 1'b1            )
  ) u_lfsr (
    .clk_i     ( clk_i      ),
    .rst_ni    ( rst_ni     ),
    .seed_en_i ( seed_en    ),
    .seed_i    ( seed       ),
    .lfsr_en_i ( lfsr_en    ),
    .entropy_i (         '0 ),
    .state_o   ( lfsr_state )
  );
  assign data_o[0] = lfsr_state;

  // A seperate permutation is applied to obtain the pseudo-random data for clearing the second
  // share of registers (e.g. key registers or state registers in case masking is enabled).
  for (genvar i = 0; i < Width; i++) begin : gen_share_perm
    assign data_o[1][i] = lfsr_state[RndCnstSharePerm[i]];
  end

  // Width must be 64.
  `ASSERT_INIT(AesPrngWidth, Width == 64)

// the code below is not meant to be synthesized,
// but it is intended to be used in simulation and FPV
`ifndef SYNTHESIS
  // Check that the supplied permutation is valid.
  logic [Width-1:0] share_perm_test, unused_share_perm_test;
  initial begin : p_share_perm_check
    share_perm_test = '0;
    for (int k = 0; k < Width; k++) begin
      share_perm_test[RndCnstSharePerm[k]] = 1'b1;
    end
    unused_share_perm_test = share_perm_test;
    // All bit positions must be marked with 1.
    `ASSERT_I(SharePermutationCheck_A, &share_perm_test)
  end
`endif

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES high-bandwidth pseudo-random number generator for masking
//
// This module uses multiple parallel LFSRs each one of them followed by an aligned permutation, a
// non-linear layer (PRINCE S-Boxes) and another permutation layer spanning across all LFSRs to
// generate pseudo-random data for masking the AES cipher core. The LFSRs can be reseeded using an
// external interface.

///////////////////////////////////////////////////////////////////////////////////////////////////
// IMPORTANT NOTE:                                                                               //
//                                   DO NOT USE THIS BLINDLY!                                    //
//                                                                                               //
// This implementation has been experimentally evaluated with / optimized for the masked AES     //
// cipher core using the S-Box implementation with first-order domain-oriented masking.          //
// Other masking schemes and S-Box implementations might have different requirements on the PRNG //
// in terms of uniformity and independence of the generated pseudo-random numbers. Upon changes  //
// to these parts of the design, it is thus recommended to again perform experimental            //
// evaluation. Use with care.                                                                    //
///////////////////////////////////////////////////////////////////////////////////////////////////

`include "prim_assert.sv"

module aes_prng_masking import aes_pkg::*;
#(
  parameter  int unsigned Width        = WidthPRDMasking,     // Must be divisble by ChunkSize and 8
  parameter  int unsigned ChunkSize    = ChunkSizePRDMasking, // Width of the LFSR primitives
  parameter  int unsigned EntropyWidth = edn_pkg::ENDPOINT_BUS_WIDTH,
  parameter  bit          SecAllowForcingMasks  = 0, // Allow forcing masks to constant values using
                                                     // force_masks_i. Useful for SCA only.
  parameter  bit          SecSkipPRNGReseeding  = 0, // The current SCA setup doesn't provide
                                                     // sufficient resources to implement the
                                                     // infrastructure required for PRNG reseeding.
                                                     // To enable SCA resistance evaluations, we
                                                     // need to skip reseeding requests.

  localparam int unsigned NumChunks = Width/ChunkSize, // derived parameter

  parameter masking_lfsr_seed_t RndCnstLfsrSeed = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t RndCnstLfsrPerm = RndCnstMaskingLfsrPermDefault
) (
  input  logic                    clk_i,
  input  logic                    rst_ni,

  input  logic                    force_masks_i,

  // Connections to AES internals, PRNG consumers
  input  logic                    data_update_i,
  output logic        [Width-1:0] data_o,
  input  logic                    reseed_req_i,
  output logic                    reseed_ack_o,

  // Connections to outer world, LFSR reseeding
  output logic                    entropy_req_o,
  input  logic                    entropy_ack_i,
  input  logic [EntropyWidth-1:0] entropy_i
);

  logic                [NumChunks-1:0] prng_seed_en;
  logic [NumChunks-1:0][ChunkSize-1:0] prng_seed;
  logic                                prng_en;
  logic [NumChunks-1:0][ChunkSize-1:0] prng_state, perm;
  logic                    [Width-1:0] prng_b, perm_b;
  logic                                phase_q;

  /////////////
  // Control //
  /////////////

  // The data requests are fed from the LFSRs. Reseed requests take precedence internally to the
  // LFSRs. If there is an outstanding reseed request, the PRNG can keep updating and providing
  // pseudo-random data (using the old seed). If the reseeding is taking place, the LFSRs will
  // provide fresh pseudo-random data (the new seed) in the next cycle anyway. This means the
  // PRNG is always ready to provide new pseudo-random data.

  // In the current SCA setup, we don't have sufficient resources to implement the infrastructure
  // required for PRNG reseeding (CSRNG, EDN, etc.). Therefore, we skip any reseeding requests if
  // the SecSkipPRNGReseeding parameter is set. Performing the reseeding without proper entropy
  // provided from CSRNG would result in quickly repeating, fully deterministic PRNG output,
  // which prevents meaningful SCA resistance evaluations.

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(AesSecAllowForcingMasksNonDefault, SecAllowForcingMasks == 0)

  if (SecAllowForcingMasks == 0) begin : gen_unused_force_masks
    logic unused_force_masks;
    assign unused_force_masks = force_masks_i;
  end

  // PRNG control
  assign prng_en = (SecAllowForcingMasks && force_masks_i) ? 1'b0 : data_update_i;

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(AesSecSkipPRNGReseedingNonDefault, SecSkipPRNGReseeding == 0)

  // Width adaption for reseeding interface. We get EntropyWidth bits at a time.
  if (ChunkSize == EntropyWidth) begin : gen_counter
    // We can reseed chunk by chunk as we get fresh entropy. Need to keep track of which chunk to
    // reseed next.
    localparam int unsigned ChunkIdxWidth = prim_util_pkg::vbits(NumChunks);
    logic [ChunkIdxWidth-1:0] chunk_idx_d, chunk_idx_q;
    logic                     prng_reseed_done;

    // Stop requesting entropy once every chunk got reseeded.
    assign entropy_req_o = SecSkipPRNGReseeding ? 1'b0         : reseed_req_i;
    assign reseed_ack_o  = SecSkipPRNGReseeding ? reseed_req_i : prng_reseed_done;

    // Counter
    assign prng_reseed_done =
        (chunk_idx_q == ChunkIdxWidth'(NumChunks - 1)) & entropy_req_o & entropy_ack_i;
    assign chunk_idx_d = prng_reseed_done ? '0                              :
        entropy_req_o && entropy_ack_i    ? chunk_idx_q + ChunkIdxWidth'(1) : chunk_idx_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin : reg_chunk_idx
      if (!rst_ni) begin
        chunk_idx_q <= '0;
      end else begin
        chunk_idx_q <= chunk_idx_d;
      end
    end

    // The entropy input is forwarded to all chunks, we just control the seed enable.
    for (genvar c = 0; c < NumChunks; c++) begin : gen_seeds
      assign prng_seed[c]    = entropy_i;
      assign prng_seed_en[c] = (c == chunk_idx_q) ? entropy_req_o & entropy_ack_i : 1'b0;
    end

  end else begin : gen_packer
    // Upsizing of entropy input to correct width for reseeding the full PRNG in one shot.
    logic [Width-1:0] seed;
    logic             seed_valid;

    // Stop requesting entropy once the desired amount is available.
    assign entropy_req_o = SecSkipPRNGReseeding ? 1'b0         : reseed_req_i & ~seed_valid;
    assign reseed_ack_o  = SecSkipPRNGReseeding ? reseed_req_i : seed_valid;

    prim_packer_fifo #(
      .InW         ( EntropyWidth ),
      .OutW        ( Width        ),
      .ClearOnRead ( 1'b0         )
    ) u_prim_packer_fifo (
      .clk_i    ( clk_i         ),
      .rst_ni   ( rst_ni        ),
      .clr_i    ( 1'b0          ), // Not needed.
      .wvalid_i ( entropy_ack_i ),
      .wdata_i  ( entropy_i     ),
      .wready_o (               ), // Not needed, we're always ready to sink data at this point.
      .rvalid_o ( seed_valid    ),
      .rdata_o  ( seed          ),
      .rready_i ( 1'b1          ), // We're always ready to receive the packed output word.
      .depth_o  (               )  // Not needed.
    );

    // Extract chunk seeds. All chunks get reseeded together.
    for (genvar c = 0; c < NumChunks; c++) begin : gen_seeds
      assign prng_seed[c]    = seed[c * ChunkSize +: ChunkSize];
      assign prng_seed_en[c] = SecSkipPRNGReseeding ? 1'b0 : seed_valid;
    end
  end

  ///////////
  // LFSRs //
  ///////////

  // We use multiple LFSR instances each having a width of ChunkSize.
  for (genvar c = 0; c < NumChunks; c++) begin : gen_lfsrs
    prim_lfsr #(
      .LfsrType     ( "GAL_XOR"                                   ),
      .LfsrDw       ( ChunkSize                                   ),
      .StateOutDw   ( ChunkSize                                   ),
      .DefaultSeed  ( RndCnstLfsrSeed[c * ChunkSize +: ChunkSize] ),
      .StatePermEn  ( 1'b0                                        ),
      .NonLinearOut ( 1'b1                                        )
    ) u_lfsr_chunk (
      .clk_i     ( clk_i           ),
      .rst_ni    ( rst_ni          ),
      .seed_en_i ( prng_seed_en[c] ),
      .seed_i    ( prng_seed[c]    ),
      .lfsr_en_i ( prng_en         ),
      .entropy_i ( '0              ),
      .state_o   ( prng_state[c]   )
    );
  end

  // Add a permutation layer spanning across all LFSRs to break linear shift patterns.
  assign prng_b = prng_state;
  for (genvar b = 0; b < Width; b++) begin : gen_perm
    assign perm_b[b] = prng_b[RndCnstLfsrPerm[b]];
  end
  assign perm = perm_b;

  /////////////
  // Outputs //
  /////////////

  // To achieve independence of input and output masks (the output mask of round X is the input
  // mask of round X+1), we assign the scrambled chunks to the output data in alternating fashion.
  assign data_o = phase_q ? {perm[0], perm[NumChunks-1:1]} : perm;

  always_ff @(posedge clk_i or negedge rst_ni) begin : reg_phase
    if (!rst_ni) begin
      phase_q <= '0;
    end else if (prng_en) begin
      phase_q <= ~phase_q;
    end
  end

  /////////////////
  // Asssertions //
  /////////////////

  // Width must be divisible by ChunkSize
  `ASSERT_INIT(AesPrngMaskingWidthByChunk, Width % ChunkSize == 0)
  // Width must be divisible by 8
  `ASSERT_INIT(AesPrngMaskingWidthBy8, Width % 8 == 0)

// the code below is not meant to be synthesized,
// but it is intended to be used in simulation and FPV
`ifndef SYNTHESIS
  // Check that the supplied permutation is valid.
  logic [Width-1:0] perm_test;
  initial begin : p_perm_check
    perm_test = '0;
    for (int k = 0; k < Width; k++) begin
      perm_test[RndCnstLfsrPerm[k]] = 1'b1;
    end
    // All bit positions must be marked with 1.
    `ASSERT_I(PermutationCheck_A, &perm_test)
  end
`endif

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES top-level wrapper

`include "prim_assert.sv"

module aes
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          AES192Enable          = 1, // Can be 0 (disable), or 1 (enable).
  parameter bit          SecMasking            = 1, // Can be 0 (no masking), or
                                                    // 1 (first-order masking) of the cipher
                                                    // core. Masking requires the use of a
                                                    // masked S-Box, see SecSBoxImpl parameter.
  parameter sbox_impl_e  SecSBoxImpl           = SBoxImplDom, // See aes_pkg.sv
  parameter int unsigned SecStartTriggerDelay  = 0, // Manual start trigger delay, useful for
                                                    // SCA measurements. A value of e.g. 40
                                                    // allows the processor to go into sleep
                                                    // before AES starts operation.
  parameter bit          SecAllowForcingMasks  = 0, // Allow forcing masks to constant values using
                                                    // FORCE_MASKS bit in Auxiliary Control
                                                    // Register. Useful for SCA only.
  parameter bit          SecSkipPRNGReseeding  = 0, // The current SCA setup doesn't provide enough
                                                    // resources to implement the infrastucture
                                                    // required for PRNG reseeding (CSRNG, EDN).
                                                    // To enable SCA resistance evaluations, we
                                                    // need to skip reseeding requests.
                                                    // Useful for SCA only.
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},
  parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingSharePerm = RndCnstClearingSharePermDefault,
  parameter masking_lfsr_seed_t  RndCnstMaskingLfsrSeed   = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t  RndCnstMaskingLfsrPerm   = RndCnstMaskingLfsrPermDefault
) (
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  input  logic                                      rst_shadowed_ni,

  // Idle indicator for clock manager
  output prim_mubi_pkg::mubi4_t                     idle_o,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t                       lc_escalate_en_i,

  // Entropy distribution network (EDN) interface
  input  logic                                      clk_edn_i,
  input  logic                                      rst_edn_ni,
  output edn_pkg::edn_req_t                         edn_o,
  input  edn_pkg::edn_rsp_t                         edn_i,

  // Key manager (keymgr) key sideload interface
  input  keymgr_pkg::hw_key_req_t                   keymgr_key_i,

  // Bus interface
  input  tlul_pkg::tl_h2d_t                         tl_i,
  output tlul_pkg::tl_d2h_t                         tl_o,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o
);

  localparam int unsigned EntropyWidth = edn_pkg::ENDPOINT_BUS_WIDTH;

  // Signals
  aes_reg2hw_t               reg2hw;
  aes_hw2reg_t               hw2reg;

  logic      [NumAlerts-1:0] alert;
  lc_ctrl_pkg::lc_tx_t       lc_escalate_en;

  logic                      edn_req_int;
  logic                      edn_req_hold_d, edn_req_hold_q;
  logic                      edn_req;
  logic                      edn_ack;
  logic   [EntropyWidth-1:0] edn_data;
  logic                      unused_edn_fips;
  logic                      entropy_clearing_req, entropy_masking_req;
  logic                      entropy_clearing_ack, entropy_masking_ack;

  ////////////
  // Inputs //
  ////////////

  // SEC_CM: BUS.INTEGRITY
  // SEC_CM: AUX.CONFIG.SHADOW
  // SEC_CM: AUX.CONFIG.REGWEN
  // SEC_CM: KEY.SW_UNREADABLE
  // SEC_CM: DATA_REG.SW_UNREADABLE
  // Register interface
  logic intg_err_alert;
  logic shadowed_storage_err, shadowed_update_err;
  aes_reg_top u_reg (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .tl_i,
    .tl_o,
    .reg2hw,
    .hw2reg,
    .shadowed_storage_err_o(shadowed_storage_err),
    .shadowed_update_err_o(shadowed_update_err),
    .intg_err_o(intg_err_alert),
    .devmode_i(1'b1)
  );

  // SEC_CM: LC_ESCALATE_EN.INTERSIG.MUBI
  // Synchronize life cycle input
  prim_lc_sync #(
    .NumCopies (1)
  ) u_prim_lc_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i ( lc_escalate_en_i ),
    .lc_en_o ( {lc_escalate_en} )
  );

  ///////////////////
  // EDN Interface //
  ///////////////////

  // Internally, we have up to two PRNGs that share the EDN interface for reseeding. Here, we just
  // arbitrate the requests. Upsizing of the entropy to the correct width is performed inside the
  // PRNGs.
  // Reseed operations for the clearing PRNG are initiated by software. Reseed operations for the
  // masking PRNG can also be automatically initiated.
  assign edn_req_int          = entropy_clearing_req | entropy_masking_req;
  // Only forward ACK to PRNG currently requesting entropy. Give higher priority to clearing PRNG.
  assign entropy_clearing_ack =  entropy_clearing_req & edn_ack;
  assign entropy_masking_ack  = ~entropy_clearing_req & entropy_masking_req & edn_ack;

  // Upon escalation or detection of a fatal alert, an EDN request signal can be dropped before
  // getting acknowledged. This is okay with respect to AES as the module will need to be reset
  // anyway. However, to not leave EDN in a strange state, we hold the request until it's actually
  // acknowledged.
  assign edn_req        = edn_req_int | edn_req_hold_q;
  assign edn_req_hold_d = (edn_req_hold_q | edn_req) & ~edn_ack;
  always_ff @(posedge clk_i or negedge rst_ni) begin : edn_req_reg
    if (!rst_ni) begin
      edn_req_hold_q <= '0;
    end else begin
      edn_req_hold_q <= edn_req_hold_d;
    end
  end

  // Synchronize EDN interface
  prim_sync_reqack_data #(
    .Width(EntropyWidth),
    .DataSrc2Dst(1'b0),
    .DataReg(1'b0)
  ) u_prim_sync_reqack_data (
    .clk_src_i  ( clk_i         ),
    .rst_src_ni ( rst_ni        ),
    .clk_dst_i  ( clk_edn_i     ),
    .rst_dst_ni ( rst_edn_ni    ),
    .req_chk_i  ( 1'b1          ),
    .src_req_i  ( edn_req       ),
    .src_ack_o  ( edn_ack       ),
    .dst_req_o  ( edn_o.edn_req ),
    .dst_ack_i  ( edn_i.edn_ack ),
    .data_i     ( edn_i.edn_bus ),
    .data_o     ( edn_data      )
  );
  // We don't track whether the entropy is pre-FIPS or not inside AES.
  assign unused_edn_fips = edn_i.edn_fips;

  //////////
  // Core //
  //////////

  // AES core
  aes_core #(
    .AES192Enable             ( AES192Enable             ),
    .SecMasking               ( SecMasking               ),
    .SecSBoxImpl              ( SecSBoxImpl              ),
    .SecStartTriggerDelay     ( SecStartTriggerDelay     ),
    .SecAllowForcingMasks     ( SecAllowForcingMasks     ),
    .SecSkipPRNGReseeding     ( SecSkipPRNGReseeding     ),
    .EntropyWidth             ( EntropyWidth             ),
    .RndCnstClearingLfsrSeed  ( RndCnstClearingLfsrSeed  ),
    .RndCnstClearingLfsrPerm  ( RndCnstClearingLfsrPerm  ),
    .RndCnstClearingSharePerm ( RndCnstClearingSharePerm ),
    .RndCnstMaskingLfsrSeed   ( RndCnstMaskingLfsrSeed   ),
    .RndCnstMaskingLfsrPerm   ( RndCnstMaskingLfsrPerm   )
  ) u_aes_core (
    .clk_i                  ( clk_i                ),
    .rst_ni                 ( rst_ni               ),
    .rst_shadowed_ni        ( rst_shadowed_ni      ),
    .entropy_clearing_req_o ( entropy_clearing_req ),
    .entropy_clearing_ack_i ( entropy_clearing_ack ),
    .entropy_clearing_i     ( edn_data             ),
    .entropy_masking_req_o  ( entropy_masking_req  ),
    .entropy_masking_ack_i  ( entropy_masking_ack  ),
    .entropy_masking_i      ( edn_data             ),

    .keymgr_key_i           ( keymgr_key_i         ),

    .lc_escalate_en_i       ( lc_escalate_en       ),

    .shadowed_storage_err_i ( shadowed_storage_err ),
    .shadowed_update_err_i  ( shadowed_update_err  ),
    .intg_err_alert_i       ( intg_err_alert       ),
    .alert_recov_o          ( alert[0]             ),
    .alert_fatal_o          ( alert[1]             ),

    .reg2hw                 ( reg2hw               ),
    .hw2reg                 ( hw2reg               )
  );

  assign idle_o = prim_mubi_pkg::mubi4_bool_to_mubi(reg2hw.status.idle.q);

  ////////////
  // Alerts //
  ////////////

  logic [NumAlerts-1:0] alert_test;
  assign alert_test = {
    reg2hw.alert_test.fatal_fault.q &
    reg2hw.alert_test.fatal_fault.qe,
    reg2hw.alert_test.recov_ctrl_update_err.q &
    reg2hw.alert_test.recov_ctrl_update_err.qe
  };

  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i)
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i] ),
      .alert_req_i   ( alert[i]      ),
      .alert_ack_o   (               ),
      .alert_state_o (               ),
      .alert_rx_i    ( alert_rx_i[i] ),
      .alert_tx_o    ( alert_tx_o[i] )
    );
  end

  ////////////////
  // Assertions //
  ////////////////

  // All outputs should have a known value after reset
  `ASSERT_KNOWN(TlODValidKnown, tl_o.d_valid)
  `ASSERT_KNOWN(TlOAReadyKnown, tl_o.a_ready)
  `ASSERT_KNOWN(IdleKnown, idle_o)
  `ASSERT_KNOWN(EdnReqKnown, edn_o)
  `ASSERT_KNOWN(AlertTxKnown, alert_tx_o)

  // Alert assertions for sparse FSMs.
  for (genvar i = 0; i < Sp2VWidth; i++) begin : gen_control_fsm_svas
    if (SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_control_fsm_svas_p
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesControlFsmCheck_A,
          u_aes_core.u_aes_control.gen_fsm[i].gen_fsm_p.
              u_aes_control_fsm_i.u_aes_control_fsm.u_state_regs,
          alert_tx_o[1])
    end else begin : gen_control_fsm_svas_n
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesControlFsmCheck_A,
          u_aes_core.u_aes_control.gen_fsm[i].gen_fsm_n.
              u_aes_control_fsm_i.u_aes_control_fsm.u_state_regs,
          alert_tx_o[1])
    end
  end

  for (genvar i = 0; i < Sp2VWidth; i++) begin : gen_ctr_fsm_svas
    if (SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_ctr_fsm_svas_p
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCtrFsmCheck_A,
          u_aes_core.u_aes_ctr.gen_fsm[i].gen_fsm_p.
              u_aes_ctr_fsm_i.u_aes_ctr_fsm.u_state_regs,
          alert_tx_o[1])
    end else begin : gen_ctr_fsm_svas_n
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCtrFsmCheck_A,
          u_aes_core.u_aes_ctr.gen_fsm[i].gen_fsm_n.
              u_aes_ctr_fsm_i.u_aes_ctr_fsm.u_state_regs,
          alert_tx_o[1])
    end
  end

  for (genvar i = 0; i < Sp2VWidth; i++) begin : gen_cipher_control_fsm_svas
    if (SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_cipher_control_fsm_svas_p
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCipherControlFsmCheck_A,
          u_aes_core.u_aes_cipher_core.u_aes_cipher_control.gen_fsm[i].gen_fsm_p.
              u_aes_cipher_control_fsm_i.u_aes_cipher_control_fsm.u_state_regs,
          alert_tx_o[1])
    end else begin : gen_cipher_control_fsm_svas_n
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCipherControlFsmCheck_A,
          u_aes_core.u_aes_cipher_core.u_aes_cipher_control.gen_fsm[i].gen_fsm_n.
              u_aes_cipher_control_fsm_i.u_aes_cipher_control_fsm.u_state_regs,
          alert_tx_o[1])
    end
  end

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module edn_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output edn_reg_pkg::edn_reg2hw_t reg2hw, // Write
  input  edn_reg_pkg::edn_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import edn_reg_pkg::* ;

  localparam int AW = 7;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [16:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(17)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_edn_cmd_req_done_qs;
  logic intr_state_edn_cmd_req_done_wd;
  logic intr_state_edn_fatal_err_qs;
  logic intr_state_edn_fatal_err_wd;
  logic intr_enable_we;
  logic intr_enable_edn_cmd_req_done_qs;
  logic intr_enable_edn_cmd_req_done_wd;
  logic intr_enable_edn_fatal_err_qs;
  logic intr_enable_edn_fatal_err_wd;
  logic intr_test_we;
  logic intr_test_edn_cmd_req_done_wd;
  logic intr_test_edn_fatal_err_wd;
  logic alert_test_we;
  logic alert_test_recov_alert_wd;
  logic alert_test_fatal_alert_wd;
  logic regwen_we;
  logic regwen_qs;
  logic regwen_wd;
  logic ctrl_we;
  logic [3:0] ctrl_edn_enable_qs;
  logic [3:0] ctrl_edn_enable_wd;
  logic [3:0] ctrl_boot_req_mode_qs;
  logic [3:0] ctrl_boot_req_mode_wd;
  logic [3:0] ctrl_auto_req_mode_qs;
  logic [3:0] ctrl_auto_req_mode_wd;
  logic [3:0] ctrl_cmd_fifo_rst_qs;
  logic [3:0] ctrl_cmd_fifo_rst_wd;
  logic boot_ins_cmd_we;
  logic [31:0] boot_ins_cmd_qs;
  logic [31:0] boot_ins_cmd_wd;
  logic boot_gen_cmd_we;
  logic [31:0] boot_gen_cmd_qs;
  logic [31:0] boot_gen_cmd_wd;
  logic sw_cmd_req_we;
  logic [31:0] sw_cmd_req_wd;
  logic sw_cmd_sts_cmd_rdy_qs;
  logic sw_cmd_sts_cmd_sts_qs;
  logic reseed_cmd_we;
  logic [31:0] reseed_cmd_wd;
  logic generate_cmd_we;
  logic [31:0] generate_cmd_wd;
  logic max_num_reqs_between_reseeds_we;
  logic [31:0] max_num_reqs_between_reseeds_qs;
  logic [31:0] max_num_reqs_between_reseeds_wd;
  logic recov_alert_sts_we;
  logic recov_alert_sts_edn_enable_field_alert_qs;
  logic recov_alert_sts_edn_enable_field_alert_wd;
  logic recov_alert_sts_boot_req_mode_field_alert_qs;
  logic recov_alert_sts_boot_req_mode_field_alert_wd;
  logic recov_alert_sts_auto_req_mode_field_alert_qs;
  logic recov_alert_sts_auto_req_mode_field_alert_wd;
  logic recov_alert_sts_cmd_fifo_rst_field_alert_qs;
  logic recov_alert_sts_cmd_fifo_rst_field_alert_wd;
  logic recov_alert_sts_edn_bus_cmp_alert_qs;
  logic recov_alert_sts_edn_bus_cmp_alert_wd;
  logic err_code_sfifo_rescmd_err_qs;
  logic err_code_sfifo_gencmd_err_qs;
  logic err_code_sfifo_output_err_qs;
  logic err_code_edn_ack_sm_err_qs;
  logic err_code_edn_main_sm_err_qs;
  logic err_code_edn_cntr_err_qs;
  logic err_code_fifo_write_err_qs;
  logic err_code_fifo_read_err_qs;
  logic err_code_fifo_state_err_qs;
  logic err_code_test_we;
  logic [4:0] err_code_test_qs;
  logic [4:0] err_code_test_wd;
  logic [8:0] main_sm_state_qs;

  // Register instances
  // R[intr_state]: V(False)
  //   F[edn_cmd_req_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_edn_cmd_req_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_edn_cmd_req_done_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.edn_cmd_req_done.de),
    .d      (hw2reg.intr_state.edn_cmd_req_done.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.edn_cmd_req_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_edn_cmd_req_done_qs)
  );

  //   F[edn_fatal_err]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_edn_fatal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_edn_fatal_err_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.edn_fatal_err.de),
    .d      (hw2reg.intr_state.edn_fatal_err.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.edn_fatal_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_edn_fatal_err_qs)
  );


  // R[intr_enable]: V(False)
  //   F[edn_cmd_req_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_edn_cmd_req_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_edn_cmd_req_done_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.edn_cmd_req_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_edn_cmd_req_done_qs)
  );

  //   F[edn_fatal_err]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_edn_fatal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_edn_fatal_err_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.edn_fatal_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_edn_fatal_err_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [1:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  //   F[edn_cmd_req_done]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_edn_cmd_req_done (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_edn_cmd_req_done_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.edn_cmd_req_done.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.edn_cmd_req_done.qe = intr_test_qe;

  //   F[edn_fatal_err]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_edn_fatal_err (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_edn_fatal_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[1]),
    .q      (reg2hw.intr_test.edn_fatal_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.edn_fatal_err.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[recov_alert]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov_alert (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_alert_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.recov_alert.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov_alert.qe = alert_test_qe;

  //   F[fatal_alert]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal_alert (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_alert_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.fatal_alert.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal_alert.qe = alert_test_qe;


  // R[regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (regwen_we),
    .wd     (regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (regwen_qs)
  );


  // R[ctrl]: V(False)
  // Create REGWEN-gated WE signal
  logic ctrl_gated_we;
  assign ctrl_gated_we = ctrl_we & regwen_qs;
  //   F[edn_enable]: 3:0
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_edn_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_edn_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.edn_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_edn_enable_qs)
  );

  //   F[boot_req_mode]: 7:4
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_boot_req_mode (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_boot_req_mode_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.boot_req_mode.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_boot_req_mode_qs)
  );

  //   F[auto_req_mode]: 11:8
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_auto_req_mode (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_auto_req_mode_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.auto_req_mode.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_auto_req_mode_qs)
  );

  //   F[cmd_fifo_rst]: 15:12
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_cmd_fifo_rst (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_cmd_fifo_rst_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.cmd_fifo_rst.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_cmd_fifo_rst_qs)
  );


  // R[boot_ins_cmd]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h901)
  ) u_boot_ins_cmd (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (boot_ins_cmd_we),
    .wd     (boot_ins_cmd_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.boot_ins_cmd.q),
    .ds     (),

    // to register interface (read)
    .qs     (boot_ins_cmd_qs)
  );


  // R[boot_gen_cmd]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'hfff003)
  ) u_boot_gen_cmd (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (boot_gen_cmd_we),
    .wd     (boot_gen_cmd_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.boot_gen_cmd.q),
    .ds     (),

    // to register interface (read)
    .qs     (boot_gen_cmd_qs)
  );


  // R[sw_cmd_req]: V(True)
  logic sw_cmd_req_qe;
  logic [0:0] sw_cmd_req_flds_we;
  assign sw_cmd_req_qe = &sw_cmd_req_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_sw_cmd_req (
    .re     (1'b0),
    .we     (sw_cmd_req_we),
    .wd     (sw_cmd_req_wd),
    .d      ('0),
    .qre    (),
    .qe     (sw_cmd_req_flds_we[0]),
    .q      (reg2hw.sw_cmd_req.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.sw_cmd_req.qe = sw_cmd_req_qe;


  // R[sw_cmd_sts]: V(False)
  //   F[cmd_rdy]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_sw_cmd_sts_cmd_rdy (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.sw_cmd_sts.cmd_rdy.de),
    .d      (hw2reg.sw_cmd_sts.cmd_rdy.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_cmd_sts_cmd_rdy_qs)
  );

  //   F[cmd_sts]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_sw_cmd_sts_cmd_sts (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.sw_cmd_sts.cmd_sts.de),
    .d      (hw2reg.sw_cmd_sts.cmd_sts.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_cmd_sts_cmd_sts_qs)
  );


  // R[reseed_cmd]: V(True)
  logic reseed_cmd_qe;
  logic [0:0] reseed_cmd_flds_we;
  assign reseed_cmd_qe = &reseed_cmd_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_reseed_cmd (
    .re     (1'b0),
    .we     (reseed_cmd_we),
    .wd     (reseed_cmd_wd),
    .d      ('0),
    .qre    (),
    .qe     (reseed_cmd_flds_we[0]),
    .q      (reg2hw.reseed_cmd.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.reseed_cmd.qe = reseed_cmd_qe;


  // R[generate_cmd]: V(True)
  logic generate_cmd_qe;
  logic [0:0] generate_cmd_flds_we;
  assign generate_cmd_qe = &generate_cmd_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_generate_cmd (
    .re     (1'b0),
    .we     (generate_cmd_we),
    .wd     (generate_cmd_wd),
    .d      ('0),
    .qre    (),
    .qe     (generate_cmd_flds_we[0]),
    .q      (reg2hw.generate_cmd.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.generate_cmd.qe = generate_cmd_qe;


  // R[max_num_reqs_between_reseeds]: V(False)
  logic max_num_reqs_between_reseeds_qe;
  logic [0:0] max_num_reqs_between_reseeds_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_max_num_reqs_between_reseeds0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&max_num_reqs_between_reseeds_flds_we),
    .q_o(max_num_reqs_between_reseeds_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_max_num_reqs_between_reseeds (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (max_num_reqs_between_reseeds_we),
    .wd     (max_num_reqs_between_reseeds_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (max_num_reqs_between_reseeds_flds_we[0]),
    .q      (reg2hw.max_num_reqs_between_reseeds.q),
    .ds     (),

    // to register interface (read)
    .qs     (max_num_reqs_between_reseeds_qs)
  );
  assign reg2hw.max_num_reqs_between_reseeds.qe = max_num_reqs_between_reseeds_qe;


  // R[recov_alert_sts]: V(False)
  //   F[edn_enable_field_alert]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_edn_enable_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_edn_enable_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.edn_enable_field_alert.de),
    .d      (hw2reg.recov_alert_sts.edn_enable_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_edn_enable_field_alert_qs)
  );

  //   F[boot_req_mode_field_alert]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_boot_req_mode_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_boot_req_mode_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.boot_req_mode_field_alert.de),
    .d      (hw2reg.recov_alert_sts.boot_req_mode_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_boot_req_mode_field_alert_qs)
  );

  //   F[auto_req_mode_field_alert]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_auto_req_mode_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_auto_req_mode_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.auto_req_mode_field_alert.de),
    .d      (hw2reg.recov_alert_sts.auto_req_mode_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_auto_req_mode_field_alert_qs)
  );

  //   F[cmd_fifo_rst_field_alert]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_cmd_fifo_rst_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_cmd_fifo_rst_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.cmd_fifo_rst_field_alert.de),
    .d      (hw2reg.recov_alert_sts.cmd_fifo_rst_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_cmd_fifo_rst_field_alert_qs)
  );

  //   F[edn_bus_cmp_alert]: 12:12
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_edn_bus_cmp_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_edn_bus_cmp_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.edn_bus_cmp_alert.de),
    .d      (hw2reg.recov_alert_sts.edn_bus_cmp_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_edn_bus_cmp_alert_qs)
  );


  // R[err_code]: V(False)
  //   F[sfifo_rescmd_err]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_rescmd_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_rescmd_err.de),
    .d      (hw2reg.err_code.sfifo_rescmd_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_rescmd_err_qs)
  );

  //   F[sfifo_gencmd_err]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_gencmd_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_gencmd_err.de),
    .d      (hw2reg.err_code.sfifo_gencmd_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_gencmd_err_qs)
  );

  //   F[sfifo_output_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_output_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_output_err.de),
    .d      (hw2reg.err_code.sfifo_output_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_output_err_qs)
  );

  //   F[edn_ack_sm_err]: 20:20
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_edn_ack_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.edn_ack_sm_err.de),
    .d      (hw2reg.err_code.edn_ack_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_edn_ack_sm_err_qs)
  );

  //   F[edn_main_sm_err]: 21:21
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_edn_main_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.edn_main_sm_err.de),
    .d      (hw2reg.err_code.edn_main_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_edn_main_sm_err_qs)
  );

  //   F[edn_cntr_err]: 22:22
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_edn_cntr_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.edn_cntr_err.de),
    .d      (hw2reg.err_code.edn_cntr_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_edn_cntr_err_qs)
  );

  //   F[fifo_write_err]: 28:28
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_write_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_write_err.de),
    .d      (hw2reg.err_code.fifo_write_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_write_err_qs)
  );

  //   F[fifo_read_err]: 29:29
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_read_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_read_err.de),
    .d      (hw2reg.err_code.fifo_read_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_read_err_qs)
  );

  //   F[fifo_state_err]: 30:30
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_state_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_state_err.de),
    .d      (hw2reg.err_code.fifo_state_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_state_err_qs)
  );


  // R[err_code_test]: V(False)
  logic err_code_test_qe;
  logic [0:0] err_code_test_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_err_code_test0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&err_code_test_flds_we),
    .q_o(err_code_test_qe)
  );
  prim_subreg #(
    .DW      (5),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (5'h0)
  ) u_err_code_test (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (err_code_test_we),
    .wd     (err_code_test_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (err_code_test_flds_we[0]),
    .q      (reg2hw.err_code_test.q),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_test_qs)
  );
  assign reg2hw.err_code_test.qe = err_code_test_qe;


  // R[main_sm_state]: V(False)
  prim_subreg #(
    .DW      (9),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (9'h185)
  ) u_main_sm_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.main_sm_state.de),
    .d      (hw2reg.main_sm_state.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (main_sm_state_qs)
  );



  logic [16:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == EDN_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == EDN_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == EDN_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == EDN_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == EDN_REGWEN_OFFSET);
    addr_hit[ 5] = (reg_addr == EDN_CTRL_OFFSET);
    addr_hit[ 6] = (reg_addr == EDN_BOOT_INS_CMD_OFFSET);
    addr_hit[ 7] = (reg_addr == EDN_BOOT_GEN_CMD_OFFSET);
    addr_hit[ 8] = (reg_addr == EDN_SW_CMD_REQ_OFFSET);
    addr_hit[ 9] = (reg_addr == EDN_SW_CMD_STS_OFFSET);
    addr_hit[10] = (reg_addr == EDN_RESEED_CMD_OFFSET);
    addr_hit[11] = (reg_addr == EDN_GENERATE_CMD_OFFSET);
    addr_hit[12] = (reg_addr == EDN_MAX_NUM_REQS_BETWEEN_RESEEDS_OFFSET);
    addr_hit[13] = (reg_addr == EDN_RECOV_ALERT_STS_OFFSET);
    addr_hit[14] = (reg_addr == EDN_ERR_CODE_OFFSET);
    addr_hit[15] = (reg_addr == EDN_ERR_CODE_TEST_OFFSET);
    addr_hit[16] = (reg_addr == EDN_MAIN_SM_STATE_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(EDN_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(EDN_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(EDN_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(EDN_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(EDN_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(EDN_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(EDN_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(EDN_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(EDN_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(EDN_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(EDN_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(EDN_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(EDN_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(EDN_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(EDN_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(EDN_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(EDN_PERMIT[16] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_edn_cmd_req_done_wd = reg_wdata[0];

  assign intr_state_edn_fatal_err_wd = reg_wdata[1];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_edn_cmd_req_done_wd = reg_wdata[0];

  assign intr_enable_edn_fatal_err_wd = reg_wdata[1];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_edn_cmd_req_done_wd = reg_wdata[0];

  assign intr_test_edn_fatal_err_wd = reg_wdata[1];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_recov_alert_wd = reg_wdata[0];

  assign alert_test_fatal_alert_wd = reg_wdata[1];
  assign regwen_we = addr_hit[4] & reg_we & !reg_error;

  assign regwen_wd = reg_wdata[0];
  assign ctrl_we = addr_hit[5] & reg_we & !reg_error;

  assign ctrl_edn_enable_wd = reg_wdata[3:0];

  assign ctrl_boot_req_mode_wd = reg_wdata[7:4];

  assign ctrl_auto_req_mode_wd = reg_wdata[11:8];

  assign ctrl_cmd_fifo_rst_wd = reg_wdata[15:12];
  assign boot_ins_cmd_we = addr_hit[6] & reg_we & !reg_error;

  assign boot_ins_cmd_wd = reg_wdata[31:0];
  assign boot_gen_cmd_we = addr_hit[7] & reg_we & !reg_error;

  assign boot_gen_cmd_wd = reg_wdata[31:0];
  assign sw_cmd_req_we = addr_hit[8] & reg_we & !reg_error;

  assign sw_cmd_req_wd = reg_wdata[31:0];
  assign reseed_cmd_we = addr_hit[10] & reg_we & !reg_error;

  assign reseed_cmd_wd = reg_wdata[31:0];
  assign generate_cmd_we = addr_hit[11] & reg_we & !reg_error;

  assign generate_cmd_wd = reg_wdata[31:0];
  assign max_num_reqs_between_reseeds_we = addr_hit[12] & reg_we & !reg_error;

  assign max_num_reqs_between_reseeds_wd = reg_wdata[31:0];
  assign recov_alert_sts_we = addr_hit[13] & reg_we & !reg_error;

  assign recov_alert_sts_edn_enable_field_alert_wd = reg_wdata[0];

  assign recov_alert_sts_boot_req_mode_field_alert_wd = reg_wdata[1];

  assign recov_alert_sts_auto_req_mode_field_alert_wd = reg_wdata[2];

  assign recov_alert_sts_cmd_fifo_rst_field_alert_wd = reg_wdata[3];

  assign recov_alert_sts_edn_bus_cmp_alert_wd = reg_wdata[12];
  assign err_code_test_we = addr_hit[15] & reg_we & !reg_error;

  assign err_code_test_wd = reg_wdata[4:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = regwen_we;
    reg_we_check[5] = ctrl_gated_we;
    reg_we_check[6] = boot_ins_cmd_we;
    reg_we_check[7] = boot_gen_cmd_we;
    reg_we_check[8] = sw_cmd_req_we;
    reg_we_check[9] = 1'b0;
    reg_we_check[10] = reseed_cmd_we;
    reg_we_check[11] = generate_cmd_we;
    reg_we_check[12] = max_num_reqs_between_reseeds_we;
    reg_we_check[13] = recov_alert_sts_we;
    reg_we_check[14] = 1'b0;
    reg_we_check[15] = err_code_test_we;
    reg_we_check[16] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_edn_cmd_req_done_qs;
        reg_rdata_next[1] = intr_state_edn_fatal_err_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_edn_cmd_req_done_qs;
        reg_rdata_next[1] = intr_enable_edn_fatal_err_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[0] = regwen_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[3:0] = ctrl_edn_enable_qs;
        reg_rdata_next[7:4] = ctrl_boot_req_mode_qs;
        reg_rdata_next[11:8] = ctrl_auto_req_mode_qs;
        reg_rdata_next[15:12] = ctrl_cmd_fifo_rst_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = boot_ins_cmd_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = boot_gen_cmd_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[9]: begin
        reg_rdata_next[0] = sw_cmd_sts_cmd_rdy_qs;
        reg_rdata_next[1] = sw_cmd_sts_cmd_sts_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = max_num_reqs_between_reseeds_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[0] = recov_alert_sts_edn_enable_field_alert_qs;
        reg_rdata_next[1] = recov_alert_sts_boot_req_mode_field_alert_qs;
        reg_rdata_next[2] = recov_alert_sts_auto_req_mode_field_alert_qs;
        reg_rdata_next[3] = recov_alert_sts_cmd_fifo_rst_field_alert_qs;
        reg_rdata_next[12] = recov_alert_sts_edn_bus_cmp_alert_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[0] = err_code_sfifo_rescmd_err_qs;
        reg_rdata_next[1] = err_code_sfifo_gencmd_err_qs;
        reg_rdata_next[2] = err_code_sfifo_output_err_qs;
        reg_rdata_next[20] = err_code_edn_ack_sm_err_qs;
        reg_rdata_next[21] = err_code_edn_main_sm_err_qs;
        reg_rdata_next[22] = err_code_edn_cntr_err_qs;
        reg_rdata_next[28] = err_code_fifo_write_err_qs;
        reg_rdata_next[29] = err_code_fifo_read_err_qs;
        reg_rdata_next[30] = err_code_fifo_state_err_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[4:0] = err_code_test_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[8:0] = main_sm_state_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: interface between a req/ack interface and a fifo
//

module edn_ack_sm (
  input logic                clk_i,
  input logic                rst_ni,

  input logic                enable_i,
  input logic                req_i,
  output logic               ack_o,
  input logic                local_escalate_i,
  input logic                fifo_not_empty_i,
  output logic               fifo_pop_o,
  output logic               fifo_clr_o,
  output logic               ack_sm_err_o
);

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 6 \
  //      -s 2299232677 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (50.00%)
  //  4: ||||||||||||| (33.33%)
  //  5: |||||| (16.67%)
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 5
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4
  //
  localparam int StateWidth = 9;
  typedef enum logic [StateWidth-1:0] {
    Disabled      = 9'b100110010, // Disabled
    EndPointClear = 9'b110001110, // Clear out end point before beginning
    Idle          = 9'b001011100, // idle (hamming distance = 3)
    DataWait      = 9'b011101011, // wait for data to return
    AckPls        = 9'b000100101, // signal ack to endpoint
    Error         = 9'b111010001  // illegal state reached and hang
  } state_e;
  state_e state_d, state_q;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, Disabled)

  always_comb begin
    state_d      = state_q;
    ack_o        = 1'b0;
    fifo_clr_o   = 1'b0;
    fifo_pop_o   = 1'b0;
    ack_sm_err_o = 1'b0;
    unique case (state_q)
      Disabled: begin
        if (enable_i) begin
          state_d = EndPointClear;
          fifo_clr_o = 1'b1;
        end
      end
      EndPointClear: begin
        state_d = Idle;
      end
      Idle: begin
        if (req_i) begin
          if (fifo_not_empty_i) begin
            fifo_pop_o = 1'b1;
          end
          state_d = DataWait;
        end
      end
      DataWait: begin
        if (fifo_not_empty_i) begin
          state_d = AckPls;
        end
      end
      AckPls: begin
        ack_o = 1'b1;
        state_d = Idle;
      end
      Error: begin
        ack_sm_err_o = 1'b1;
      end
      default: begin
        ack_sm_err_o = 1'b1;
        state_d = Error;
      end
    endcase // unique case (state_q)

    // If local escalation is seen, transition directly to
    // error state.
    if (local_escalate_i) begin
      state_d = Error;
      // Tie off outputs, except for ack_sm_err_o.
      ack_o      = 1'b0;
      fifo_clr_o = 1'b0;
      fifo_pop_o = 1'b0;
    end else if (!enable_i && state_q inside {EndPointClear, Idle, DataWait, AckPls}) begin
      // Only disable if state is legal and not Disabled or Error.
      // Even when disabled, illegal states must result in a transition to Error.
      state_d = Disabled;
      // Tie off all outputs, except for ack_sm_err_o.
      ack_o        = 1'b0;
      fifo_pop_o   = 1'b0;
      fifo_clr_o   = 1'b0;
    end
  end

  // The `local_escalate_i` includes `ack_sm_err_o`.
  // The following assertion ensures the Error state is stable until reset.
  // With `FpvSecCm` prefix, this assertion will added to weekly FPV sec_cm regression.
  `ASSERT(FpvSecCmErrorStEscalate_A, state_q == Error |-> local_escalate_i)

  // This assertion does not have `FpvSecCm` prefix because the sec_cm FPV environment will
  // blackbox the `prim_sparse_fsm` `state_q` output.
  `ASSERT(AckSmErrorStStable_A,   state_q == Error |=> $stable(state_q))

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: edn csrng application request state machine module
//
//   does hardware-based csrng app interface command requests

module edn_main_sm import edn_pkg::*; #(
  localparam int StateWidth = 9
) (
  input logic                   clk_i,
  input logic                   rst_ni,

  input logic                   edn_enable_i,
  input logic                   boot_req_mode_i,
  input logic                   auto_req_mode_i,
  input logic                   sw_cmd_req_load_i,
  output logic                  sw_cmd_valid_o,
  output logic                  boot_wr_cmd_reg_o,
  output logic                  boot_wr_cmd_genfifo_o,
  output logic                  auto_set_intr_gate_o,
  output logic                  auto_clr_intr_gate_o,
  output logic                  auto_first_ack_wait_o,
  output logic                  main_sm_done_pulse_o,
  input logic                   csrng_cmd_ack_i,
  output logic                  capt_gencmd_fifo_cnt_o,
  output logic                  boot_send_gencmd_o,
  output logic                  send_gencmd_o,
  input logic                   max_reqs_cnt_zero_i,
  output logic                  capt_rescmd_fifo_cnt_o,
  output logic                  send_rescmd_o,
  input logic                   cmd_sent_i,
  input logic                   local_escalate_i,
  output logic                  auto_req_mode_busy_o,
  output logic                  main_sm_busy_o,
  output logic [StateWidth-1:0] main_sm_state_o,
  output logic                  main_sm_err_o
);
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: ||||||||||| (17.54%)
//  4: |||||||||||||||||||| (29.82%)
//  5: ||||||||||||||||| (26.32%)
//  6: ||||||||||| (17.54%)
//  7: ||||| (7.60%)
//  8:  (1.17%)
//  9: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 8
// Minimum Hamming weight: 2
// Maximum Hamming weight: 7
//

  state_e state_d, state_q;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, Idle)

  assign main_sm_state_o = state_q;

  assign main_sm_busy_o = (state_q != Idle) && (state_q != BootPulse) &&
         (state_q != BootDone) && (state_q != SWPortMode);

  always_comb begin
    state_d                = state_q;
    boot_wr_cmd_reg_o      = 1'b0;
    boot_wr_cmd_genfifo_o  = 1'b0;
    boot_send_gencmd_o     = 1'b0;
    auto_set_intr_gate_o   = 1'b0;
    auto_clr_intr_gate_o   = 1'b0;
    auto_first_ack_wait_o  = 1'b0;
    auto_req_mode_busy_o   = 1'b0;
    capt_gencmd_fifo_cnt_o = 1'b0;
    send_gencmd_o          = 1'b0;
    capt_rescmd_fifo_cnt_o = 1'b0;
    send_rescmd_o          = 1'b0;
    main_sm_done_pulse_o   = 1'b0;
    main_sm_err_o          = 1'b0;
    sw_cmd_valid_o         = 1'b1;
    unique case (state_q)
      Idle: begin
        if (boot_req_mode_i && edn_enable_i) begin
          state_d = BootLoadIns;
        end else if (auto_req_mode_i && edn_enable_i) begin
          state_d = AutoLoadIns;
        end else if (edn_enable_i) begin
          main_sm_done_pulse_o = 1'b1;
          state_d = SWPortMode;
        end
      end
      BootLoadIns: begin
        boot_wr_cmd_reg_o = 1'b1;
        state_d = BootLoadGen;
      end
      BootLoadGen: begin
        boot_wr_cmd_genfifo_o = 1'b1;
        state_d = BootInsAckWait;
      end
      BootInsAckWait: begin
        if (csrng_cmd_ack_i) begin
          state_d = BootCaptGenCnt;
        end
      end
      BootCaptGenCnt: begin
        capt_gencmd_fifo_cnt_o = 1'b1;
        state_d = BootSendGenCmd;
      end
      BootSendGenCmd: begin
        boot_send_gencmd_o = 1'b1;
        if (cmd_sent_i) begin
          state_d = BootGenAckWait;
        end
      end
      BootGenAckWait: begin
        if (csrng_cmd_ack_i) begin
          state_d = BootPulse;
        end
      end
      BootPulse: begin
        main_sm_done_pulse_o = 1'b1;
        state_d = BootDone;
      end
      BootDone: begin
      end
      //-----------------------------------
      AutoLoadIns: begin
        auto_set_intr_gate_o = 1'b1;
        auto_first_ack_wait_o = 1'b1;
        if (sw_cmd_req_load_i) begin
          state_d = AutoFirstAckWait;
        end
      end
      AutoFirstAckWait: begin
        auto_first_ack_wait_o = 1'b1;
        if (csrng_cmd_ack_i) begin
          auto_clr_intr_gate_o = 1'b1;
          state_d = AutoDispatch;
        end
      end
      AutoAckWait: begin
        sw_cmd_valid_o = 1'b0;
        auto_req_mode_busy_o = 1'b1;
        if (csrng_cmd_ack_i) begin
          state_d = AutoDispatch;
        end
      end
      AutoDispatch: begin
        auto_req_mode_busy_o = 1'b1;
        sw_cmd_valid_o = 1'b0;
        if (!auto_req_mode_i) begin
          main_sm_done_pulse_o = 1'b1;
          state_d = Idle;
        end else begin
          if (max_reqs_cnt_zero_i) begin
            state_d = AutoCaptReseedCnt;
          end else begin
            state_d = AutoCaptGenCnt;
          end
        end
      end
      AutoCaptGenCnt: begin
        sw_cmd_valid_o = 1'b0;
        auto_req_mode_busy_o = 1'b1;
        capt_gencmd_fifo_cnt_o = 1'b1;
        state_d = AutoSendGenCmd;
      end
      AutoSendGenCmd: begin
        sw_cmd_valid_o = 1'b0;
        auto_req_mode_busy_o = 1'b1;
        send_gencmd_o = 1'b1;
        if (cmd_sent_i) begin
          state_d = AutoAckWait;
        end
      end
      AutoCaptReseedCnt: begin
        sw_cmd_valid_o = 1'b0;
        auto_req_mode_busy_o = 1'b1;
        capt_rescmd_fifo_cnt_o = 1'b1;
        state_d = AutoSendReseedCmd;
      end
      AutoSendReseedCmd: begin
        sw_cmd_valid_o = 1'b0;
        auto_req_mode_busy_o = 1'b1;
        send_rescmd_o = 1'b1;
        if (cmd_sent_i) begin
          state_d = AutoAckWait;
        end
      end
      SWPortMode: begin
      end
      Error: begin
        main_sm_err_o = 1'b1;
      end
      default: begin
        state_d = Error;
        main_sm_err_o = 1'b1;
      end
    endcase

    if (local_escalate_i) begin
      state_d = Error;
      // Tie off outputs, except for main_sm_err_o.
      boot_wr_cmd_reg_o      = 1'b0;
      boot_wr_cmd_genfifo_o  = 1'b0;
      boot_send_gencmd_o     = 1'b0;
      auto_set_intr_gate_o   = 1'b0;
      auto_clr_intr_gate_o   = 1'b0;
      auto_first_ack_wait_o  = 1'b0;
      auto_req_mode_busy_o   = 1'b0;
      capt_gencmd_fifo_cnt_o = 1'b0;
      send_gencmd_o          = 1'b0;
      capt_rescmd_fifo_cnt_o = 1'b0;
      send_rescmd_o          = 1'b0;
      main_sm_done_pulse_o   = 1'b0;
    end else if (!edn_enable_i && state_q inside {BootLoadIns, BootLoadGen, BootInsAckWait,
                                                  BootCaptGenCnt, BootSendGenCmd, BootGenAckWait,
                                                  BootPulse, BootDone, AutoLoadIns,
                                                  AutoFirstAckWait, AutoAckWait, AutoDispatch,
                                                  AutoCaptGenCnt, AutoSendGenCmd,
                                                  AutoCaptReseedCnt, AutoSendReseedCmd, SWPortMode
                                                 }) begin
      // Only go to idle if the state is legal and not Idle or Error.
      // Even when disabled, illegal states must result in a transition to Error.
      state_d = Idle;
      // Tie off outputs, except for main_sm_err_o.
      boot_wr_cmd_reg_o      = 1'b0;
      boot_wr_cmd_genfifo_o  = 1'b0;
      boot_send_gencmd_o     = 1'b0;
      auto_set_intr_gate_o   = 1'b0;
      auto_clr_intr_gate_o   = 1'b0;
      auto_first_ack_wait_o  = 1'b0;
      auto_req_mode_busy_o   = 1'b0;
      capt_gencmd_fifo_cnt_o = 1'b0;
      send_gencmd_o          = 1'b0;
      capt_rescmd_fifo_cnt_o = 1'b0;
      send_rescmd_o          = 1'b0;
      main_sm_done_pulse_o   = 1'b0;
    end
  end

  // The `local_escalate_i` includes `main_sm_err_o`.
  // The following assertion ensures the Error state is stable until reset.
  // With `FpvSecCm` prefix, this assertion will added to weekly FPV sec_cm regression.
  `ASSERT(FpvSecCmErrorStEscalate_A, state_q == Error |-> local_escalate_i)

  // This assertion does not have `FpvSecCm` prefix because the sec_cm FPV environment will
  // blackbox the `prim_sparse_fsm` `state_q` output.
  `ASSERT(ErrorStStable_A, state_q == Error |=> $stable(state_q))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy distrubution network core module
//  - this module will make requests to the CSRNG module
//    and return the genbits back to up four requesting
//    end points.
//

module edn_core import edn_pkg::*;
#(
  parameter int NumEndPoints = 4
) (
  input logic clk_i,
  input logic rst_ni,

  input  edn_reg_pkg::edn_reg2hw_t reg2hw,
  output edn_reg_pkg::edn_hw2reg_t hw2reg,

  // EDN interfaces
  input  edn_req_t [NumEndPoints-1:0] edn_i,
  output edn_rsp_t [NumEndPoints-1:0] edn_o,

  // CSRNG Application Interface
  output  csrng_pkg::csrng_req_t  csrng_cmd_o,
  input   csrng_pkg::csrng_rsp_t  csrng_cmd_i,

  // Alerts
  output logic        recov_alert_test_o,
  output logic        fatal_alert_test_o,
  output logic        recov_alert_o,
  output logic        fatal_alert_o,

  // Interrupts
  output logic        intr_edn_cmd_req_done_o,
  output logic        intr_edn_fatal_err_o
);

  import edn_reg_pkg::*;

  localparam int RegWidth = 32;
  localparam int RescmdFifoWidth = 32;
  localparam int RescmdFifoDepth = 13;
  localparam int GencmdFifoWidth = 32;
  localparam int GencmdFifoDepth = 13;
  localparam int OutputFifoWidth = 32;
  localparam int OutputFifoDepth = 13;
  localparam int CSGenBitsWidth = 128;
  localparam int EndPointBusWidth = 32;
  localparam int RescmdFifoIdxWidth = $clog2(RescmdFifoDepth);
  localparam int FifoRstCopies = 4;
  localparam int BootReqCopies = 2;

  typedef enum logic [4:0] {
    MuBiCheck,
    FatalErr,
    ReseedCmdErr,
    GenCmdErr,
    OutputErr,
    FifoWrErr,
    FifoRdErr,
    FifoStErr,
    CsrngCmdReq,
    CsrngCmdReqValid,
    CsrngCmdReqOut,
    CsrngCmdReqValidOut,
    EnDelay,
    IntrStatus,
    SendReseedCmd,
    SendGenCmd,
    OutputClr,
    MainFsmEn,
    CmdFifoCnt,
    CsrngPackerClr,
    CsrngFipsEn,
    CsrngDataVld,
    AckFsmEn,
    LastEdnEntry
  } edn_enable_e;
  localparam int EdnEnableCopies = int'(LastEdnEntry);

  // signals
  logic event_edn_cmd_req_done;
  logic event_edn_fatal_err;
  logic [EdnEnableCopies-1:FatalErr] edn_enable_fo;
  logic [FifoRstCopies-1:1] cmd_fifo_rst_fo;
  logic [BootReqCopies-1:1] boot_req_mode_fo;
  logic edn_enable_pfa;
  logic cmd_fifo_rst_pfa;
  logic packer_arb_valid;
  logic packer_arb_ready;
  logic [NumEndPoints-1:0] packer_arb_req;
  logic [NumEndPoints-1:0] packer_arb_gnt;
  logic                    auto_req_mode_pfe;
  logic                    auto_req_mode_pfa;
  logic                    main_sm_done_pulse;
  logic                    main_sm_busy;
  logic                    capt_gencmd_fifo_cnt;
  logic                    capt_rescmd_fifo_cnt;
  logic                    max_reqs_cnt_zero;
  logic                    max_reqs_cnt_load;
  logic                    max_reqs_between_reseed_load;
  logic [31:0]             max_reqs_between_reseed_bus;
  logic                    csrng_cmd_ack;
  logic                    csrng_cmd_ack_gated;
  logic                    send_rescmd;
  logic                    cmd_sent;
  logic                    send_gencmd;
  logic                    boot_send_gencmd;
  logic                    sw_cmd_req_load;
  logic                    sw_cmd_valid;
  logic [31:0]             sw_cmd_req_bus;
  logic                    reseed_cmd_load;
  logic [31:0]             reseed_cmd_bus;
  logic                    generate_cmd_load;
  logic [31:0]             generate_cmd_bus;
  logic                    packer_cs_clr;
  logic                    packer_cs_push;
  logic [CSGenBitsWidth-1:0] packer_cs_wdata;
  logic                      packer_cs_wready;
  logic                      packer_cs_rvalid;
  logic                      packer_cs_rready;
  logic [CSGenBitsWidth-1:0] packer_cs_rdata;
  logic                      boot_req_mode_pfa;
  logic                      boot_wr_cmd_reg;
  logic                      boot_wr_cmd_genfifo;
  logic                      auto_first_ack_wait;
  logic                      auto_req_mode_busy;
  logic                      auto_set_intr_gate;
  logic                      auto_clr_intr_gate;

  logic [NumEndPoints-1:0]   packer_ep_clr;
  logic [NumEndPoints-1:0]   packer_ep_ack;
  logic [NumEndPoints-1:0]   packer_ep_push;
  logic [CSGenBitsWidth-1:0] packer_ep_wdata [NumEndPoints];
  logic [NumEndPoints-1:0]   packer_ep_wready;
  logic [NumEndPoints-1:0]   packer_ep_rvalid;
  logic [NumEndPoints-1:0]   packer_ep_rready;
  logic                      edn_ack_sm_err_sum;
  logic [NumEndPoints-1:0]   edn_ack_sm_err;
  logic [EndPointBusWidth-1:0] packer_ep_rdata [NumEndPoints];

  // rescmd fifo
  logic [RescmdFifoIdxWidth-1:0]      sfifo_rescmd_depth;
  logic [RescmdFifoWidth-1:0]         sfifo_rescmd_rdata;
  logic                               sfifo_rescmd_clr;
  logic                               sfifo_rescmd_push;
  logic [RescmdFifoWidth-1:0]         sfifo_rescmd_wdata;
  logic                               sfifo_rescmd_pop;
  logic                               sfifo_rescmd_err_sum;
  logic [2:0]                         sfifo_rescmd_err;
  logic                               sfifo_rescmd_full;
  logic                               sfifo_rescmd_not_empty;

  // gencmd fifo
  logic [GencmdFifoWidth-1:0]         sfifo_gencmd_rdata;
  logic [$clog2(GencmdFifoDepth)-1:0] sfifo_gencmd_depth;
  logic                               sfifo_gencmd_clr;
  logic                               sfifo_gencmd_push;
  logic [GencmdFifoWidth-1:0]         sfifo_gencmd_wdata;
  logic                               sfifo_gencmd_pop;
  logic                               sfifo_gencmd_err_sum;
  logic [2:0]                         sfifo_gencmd_err;
  logic                               sfifo_gencmd_full;
  logic                               sfifo_gencmd_not_empty;

  // output fifo
  logic [OutputFifoWidth-1:0]         sfifo_output_rdata;
  logic                               sfifo_output_clr;
  logic                               sfifo_output_push;
  logic [OutputFifoWidth-1:0]         sfifo_output_wdata;
  logic                               sfifo_output_pop;
  logic                               sfifo_output_full;
  logic                               sfifo_output_err_sum;
  logic [2:0]                         sfifo_output_err;
  logic                               sfifo_output_not_empty;

  logic                               edn_main_sm_err_sum;
  logic [8:0]                         edn_main_sm_state;
  logic                               edn_main_sm_err;
  logic [30:0]                        err_code_test_bit;
  logic                               fifo_write_err_sum;
  logic                               fifo_read_err_sum;
  logic                               fifo_status_err_sum;
  logic                               cs_rdata_capt_vld;
  logic                               edn_bus_cmp_alert;
  logic                               edn_cntr_err_sum;
  logic                               edn_cntr_err;
  logic [RegWidth-1:0]                max_reqs_cnt;
  logic                               max_reqs_cnt_err;
  logic                               cmd_rdy;
  logic [31:0]                        boot_ins_cmd;
  logic [31:0]                        boot_gen_cmd;

  // unused
  logic                               unused_err_code_test_bit;

  import prim_mubi_pkg::mubi4_t;
  import prim_mubi_pkg::mubi4_test_true_strict;
  import prim_mubi_pkg::mubi4_test_invalid;

  prim_mubi_pkg::mubi4_t [EdnEnableCopies-1:0] mubi_edn_enable_fanout;
  prim_mubi_pkg::mubi4_t [FifoRstCopies-1:0] mubi_cmd_fifo_rst_fanout;
  prim_mubi_pkg::mubi4_t [BootReqCopies-1:0] mubi_boot_req_mode_fanout;
  prim_mubi_pkg::mubi4_t [1:0] mubi_auto_req_mode_fanout;

  // flops
  logic [31:0]                        cs_cmd_req_q, cs_cmd_req_d;
  logic                               cs_cmd_req_vld_q, cs_cmd_req_vld_d;
  logic [31:0]                        cs_cmd_req_out_q, cs_cmd_req_out_d;
  logic                               cs_cmd_req_vld_out_q, cs_cmd_req_vld_out_d;
  logic [RescmdFifoIdxWidth-1:0]      cmd_fifo_cnt_q, cmd_fifo_cnt_d;
  logic                               send_rescmd_q, send_rescmd_d;
  logic                               send_gencmd_q, send_gencmd_d;
  logic                               csrng_fips_q, csrng_fips_d;
  logic [NumEndPoints-1:0]            edn_fips_q, edn_fips_d;
  logic [63:0]                        cs_rdata_capt_q, cs_rdata_capt_d;
  logic                               cs_rdata_capt_vld_q, cs_rdata_capt_vld_d;
  logic                               sw_rdy_sts_q, sw_rdy_sts_d;
  logic                               intr_sts_gate_q, intr_sts_gate_d;
  logic                               edn_enable_q, edn_enable_d;

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      cs_cmd_req_q  <= '0;
      cs_cmd_req_vld_q  <= '0;
      cs_cmd_req_out_q  <= '0;
      cs_cmd_req_vld_out_q  <= '0;
      cmd_fifo_cnt_q <= '0;
      send_rescmd_q <= '0;
      send_gencmd_q <= '0;
      csrng_fips_q <= '0;
      edn_fips_q <= '0;
      cs_rdata_capt_q <= '0;
      cs_rdata_capt_vld_q <= '0;
      sw_rdy_sts_q   <= '0;
      intr_sts_gate_q   <= '0;
      edn_enable_q  <= '0;
    end else begin
      cs_cmd_req_q  <= cs_cmd_req_d;
      cs_cmd_req_vld_q  <= cs_cmd_req_vld_d;
      cs_cmd_req_out_q <= cs_cmd_req_out_d;
      cs_cmd_req_vld_out_q <= cs_cmd_req_vld_out_d;
      cmd_fifo_cnt_q <= cmd_fifo_cnt_d;
      send_rescmd_q <= send_rescmd_d;
      send_gencmd_q <= send_gencmd_d;
      csrng_fips_q <= csrng_fips_d;
      edn_fips_q <= edn_fips_d;
      cs_rdata_capt_q <= cs_rdata_capt_d;
      cs_rdata_capt_vld_q <= cs_rdata_capt_vld_d;
      sw_rdy_sts_q   <= sw_rdy_sts_d;
      intr_sts_gate_q   <= intr_sts_gate_d;
      edn_enable_q  <= edn_enable_d;
    end

  //--------------------------------------------
  // instantiate interrupt hardware primitives
  //--------------------------------------------

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_edn_cmd_req_done (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_edn_cmd_req_done),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.edn_cmd_req_done.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.edn_cmd_req_done.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.edn_cmd_req_done.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.edn_cmd_req_done.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.edn_cmd_req_done.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.edn_cmd_req_done.d),
    .intr_o                 (intr_edn_cmd_req_done_o)
  );


  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_edn_fatal_err (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_edn_fatal_err),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.edn_fatal_err.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.edn_fatal_err.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.edn_fatal_err.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.edn_fatal_err.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.edn_fatal_err.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.edn_fatal_err.d),
    .intr_o                 (intr_edn_fatal_err_o)
  );

  // interrupt for sw app interface only
  assign event_edn_cmd_req_done = csrng_cmd_ack_gated;

  // Counter and fsm errors are structural errors and are always
  // active regardless of the functional state.
  logic fatal_loc_events;
  assign fatal_loc_events =  edn_cntr_err_sum ||
                             edn_main_sm_err_sum ||
                             edn_ack_sm_err_sum;

  // set the interrupt sources
  assign event_edn_fatal_err = (edn_enable_fo[FatalErr] && (
         sfifo_rescmd_err_sum ||
         sfifo_gencmd_err_sum ||
         sfifo_output_err_sum )) ||
         fatal_loc_events;

  // set fifo errors that are single instances of source
  assign sfifo_rescmd_err_sum = (|sfifo_rescmd_err) ||
         err_code_test_bit[0];
  assign sfifo_gencmd_err_sum = (|sfifo_gencmd_err) ||
         err_code_test_bit[1];
  assign sfifo_output_err_sum = (|sfifo_output_err) ||
         err_code_test_bit[2];
  assign edn_ack_sm_err_sum = (|edn_ack_sm_err) ||
         err_code_test_bit[20];
  assign edn_main_sm_err_sum = edn_main_sm_err ||
         err_code_test_bit[21];
  assign edn_cntr_err_sum = edn_cntr_err ||
         err_code_test_bit[22];

  assign fifo_write_err_sum =
         sfifo_rescmd_err[2] ||
         sfifo_gencmd_err[2] ||
         sfifo_output_err[2] ||
         err_code_test_bit[28];
  assign fifo_read_err_sum =
         sfifo_rescmd_err[1] ||
         sfifo_gencmd_err[1] ||
         sfifo_output_err[1] ||
         err_code_test_bit[29];
  assign fifo_status_err_sum =
         sfifo_rescmd_err[0] ||
         sfifo_gencmd_err[0] ||
         sfifo_output_err[0] ||
         err_code_test_bit[30];


  // set the err code source bits
  assign hw2reg.err_code.sfifo_rescmd_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_rescmd_err.de = edn_enable_fo[ReseedCmdErr] && sfifo_rescmd_err_sum;

  assign hw2reg.err_code.sfifo_gencmd_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_gencmd_err.de = edn_enable_fo[GenCmdErr] && sfifo_gencmd_err_sum;

  assign hw2reg.err_code.sfifo_output_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_output_err.de = edn_enable_fo[OutputErr] && sfifo_output_err_sum;

  assign hw2reg.err_code.edn_ack_sm_err.d = 1'b1;
  assign hw2reg.err_code.edn_ack_sm_err.de = edn_ack_sm_err_sum;

  assign hw2reg.err_code.edn_main_sm_err.d = 1'b1;
  assign hw2reg.err_code.edn_main_sm_err.de = edn_main_sm_err_sum;

  assign hw2reg.err_code.edn_cntr_err.d = 1'b1;
  assign hw2reg.err_code.edn_cntr_err.de = edn_cntr_err_sum;

  assign boot_ins_cmd = reg2hw.boot_ins_cmd.q;
  assign boot_gen_cmd = reg2hw.boot_gen_cmd.q;


 // set the err code type bits
  assign hw2reg.err_code.fifo_write_err.d = 1'b1;
  assign hw2reg.err_code.fifo_write_err.de = edn_enable_fo[FifoWrErr] && fifo_write_err_sum;

  assign hw2reg.err_code.fifo_read_err.d = 1'b1;
  assign hw2reg.err_code.fifo_read_err.de = edn_enable_fo[FifoRdErr] && fifo_read_err_sum;

  assign hw2reg.err_code.fifo_state_err.d = 1'b1;
  assign hw2reg.err_code.fifo_state_err.de = edn_enable_fo[FifoStErr] && fifo_status_err_sum;


  // Error forcing
  for (genvar i = 0; i < 31; i = i+1) begin : gen_err_code_test_bit
    assign err_code_test_bit[i] = (reg2hw.err_code_test.q == i) && reg2hw.err_code_test.qe;
  end : gen_err_code_test_bit


  // alert - send all interrupt sources to the alert for the fatal case
  assign fatal_alert_o = event_edn_fatal_err;

  // alert test
  assign recov_alert_test_o = {
    reg2hw.alert_test.recov_alert.q &&
    reg2hw.alert_test.recov_alert.qe
  };
  assign fatal_alert_test_o = {
    reg2hw.alert_test.fatal_alert.q &&
    reg2hw.alert_test.fatal_alert.qe
  };

  // check for illegal enable field states, and set alert if detected

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_edn_enable;
  assign mubi_edn_enable = mubi4_t'(reg2hw.ctrl.edn_enable.q);
  assign edn_enable_pfa = mubi4_test_invalid(mubi_edn_enable_fanout[MuBiCheck]);
  assign hw2reg.recov_alert_sts.edn_enable_field_alert.de = edn_enable_pfa;
  assign hw2reg.recov_alert_sts.edn_enable_field_alert.d  = edn_enable_pfa;

  for (genvar i = int'(FatalErr); i < LastEdnEntry; i = i+1) begin : gen_mubi_en_copies
    assign edn_enable_fo[i] = mubi4_test_true_strict(mubi_edn_enable_fanout[i]);
  end : gen_mubi_en_copies

  prim_mubi4_sync #(
    .NumCopies(EdnEnableCopies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_edn_enable (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_edn_enable),
    .mubi_o(mubi_edn_enable_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_cmd_fifo_rst;
  assign mubi_cmd_fifo_rst = mubi4_t'(reg2hw.ctrl.cmd_fifo_rst.q);
  assign cmd_fifo_rst_pfa = mubi4_test_invalid(mubi_cmd_fifo_rst_fanout[0]);
  assign hw2reg.recov_alert_sts.cmd_fifo_rst_field_alert.de = cmd_fifo_rst_pfa;
  assign hw2reg.recov_alert_sts.cmd_fifo_rst_field_alert.d  = cmd_fifo_rst_pfa;

  for (genvar i = 1; i < FifoRstCopies; i = i+1) begin : gen_mubi_rst_copies
    assign cmd_fifo_rst_fo[i] = mubi4_test_true_strict(mubi_cmd_fifo_rst_fanout[i]);
  end : gen_mubi_rst_copies

  prim_mubi4_sync #(
    .NumCopies(FifoRstCopies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_cmd_fifo_rst (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_cmd_fifo_rst),
    .mubi_o(mubi_cmd_fifo_rst_fanout)
  );

  // counter errors
  assign edn_cntr_err = max_reqs_cnt_err;

  //--------------------------------------------
  // sw register interface
  //--------------------------------------------
  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_auto_req_mode;
  assign mubi_auto_req_mode = mubi4_t'(reg2hw.ctrl.auto_req_mode.q);
  assign auto_req_mode_pfe = mubi4_test_true_strict(mubi_auto_req_mode_fanout[0]);
  assign auto_req_mode_pfa = mubi4_test_invalid(mubi_auto_req_mode_fanout[1]);
  assign hw2reg.recov_alert_sts.auto_req_mode_field_alert.de = auto_req_mode_pfa;
  assign hw2reg.recov_alert_sts.auto_req_mode_field_alert.d  = auto_req_mode_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_auto_req_mode (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_auto_req_mode),
    .mubi_o(mubi_auto_req_mode_fanout)
  );


  // SW interface connection
  // cmd req
  assign sw_cmd_req_load = reg2hw.sw_cmd_req.qe & sw_cmd_valid;
  assign sw_cmd_req_bus = reg2hw.sw_cmd_req.q;

  assign max_reqs_between_reseed_load = reg2hw.max_num_reqs_between_reseeds.qe;
  assign max_reqs_between_reseed_bus = reg2hw.max_num_reqs_between_reseeds.q;

  assign reseed_cmd_load = reg2hw.reseed_cmd.qe;
  assign reseed_cmd_bus = reg2hw.reseed_cmd.q;

  assign generate_cmd_load = reg2hw.generate_cmd.qe;
  assign generate_cmd_bus = reg2hw.generate_cmd.q;

  assign cs_cmd_req_d =
         (!edn_enable_fo[CsrngCmdReq]) ? '0 :
         boot_wr_cmd_reg ? boot_ins_cmd :
         sw_cmd_req_load ? sw_cmd_req_bus :
         cs_cmd_req_q;

  assign cs_cmd_req_vld_d =
         (!edn_enable_fo[CsrngCmdReqValid]) ? '0 :
         (sw_cmd_req_load || boot_wr_cmd_reg); // cmd reg write

  assign cs_cmd_req_out_d =
         (!edn_enable_fo[CsrngCmdReqOut]) ? '0 :
         send_rescmd ? sfifo_rescmd_rdata :
         (send_gencmd || boot_send_gencmd) ? sfifo_gencmd_rdata :
         cs_cmd_req_q;

  assign cs_cmd_req_vld_out_d =
         (!edn_enable_fo[CsrngCmdReqValidOut]) ? '0 :
         (send_rescmd || send_gencmd || (boot_send_gencmd && cmd_sent)) ? 1'b1 :
         cs_cmd_req_vld_q;


  // receive rdy
  assign hw2reg.sw_cmd_sts.cmd_rdy.de = 1'b1;
  assign hw2reg.sw_cmd_sts.cmd_rdy.d = cmd_rdy;
  assign cmd_rdy = !sw_cmd_req_load && sw_rdy_sts_q;
  assign sw_rdy_sts_d =
         !edn_enable_q ? 1'b0 :
         sw_cmd_req_load ? 1'b0 :
         auto_first_ack_wait ? 1'b1 :
         main_sm_busy ? 1'b0 :
         csrng_cmd_i.csrng_req_ready ? 1'b1 :
         sw_rdy_sts_q;

  assign edn_enable_d = edn_enable_fo[EnDelay];

  // receive cmd ack
  assign csrng_cmd_ack = csrng_cmd_i.csrng_rsp_ack;
  assign csrng_cmd_ack_gated = csrng_cmd_ack && intr_sts_gate_q;
  assign hw2reg.sw_cmd_sts.cmd_sts.de = csrng_cmd_ack_gated;
  assign hw2reg.sw_cmd_sts.cmd_sts.d = csrng_cmd_i.csrng_rsp_sts;

  assign intr_sts_gate_d =
         !edn_enable_fo[IntrStatus] ? 1'b0 :
         main_sm_done_pulse ? 1'b1 :
         auto_set_intr_gate ? 1'b1 :
         auto_clr_intr_gate ? 1'b0 :
         intr_sts_gate_q;

  // rescmd fifo
  prim_fifo_sync #(
    .Width(RescmdFifoWidth),
    .Pass(0),
    .Depth(RescmdFifoDepth)
  ) u_prim_fifo_sync_rescmd (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (sfifo_rescmd_clr),
    .wvalid_i (sfifo_rescmd_push),
    .wready_o (),
    .wdata_i  (sfifo_rescmd_wdata),
    .rvalid_o (sfifo_rescmd_not_empty),
    .rready_i (sfifo_rescmd_pop),
    .rdata_o  (sfifo_rescmd_rdata),
    .full_o   (sfifo_rescmd_full),
    .depth_o  (sfifo_rescmd_depth),
    .err_o    ()
  );

  // feedback cmd back into rescmd fifo
  assign send_rescmd_d = send_rescmd;

  assign sfifo_rescmd_push =
         (send_rescmd_q & edn_enable_fo[SendReseedCmd]) ? 1'b1  :
         reseed_cmd_load;

  assign sfifo_rescmd_wdata =
         auto_req_mode_busy ? cs_cmd_req_out_q :
         reseed_cmd_bus;

  assign sfifo_rescmd_pop = send_rescmd;

  assign sfifo_rescmd_clr = (cmd_fifo_rst_fo[1] || main_sm_done_pulse);

  assign sfifo_rescmd_err =
         {(sfifo_rescmd_push && sfifo_rescmd_full),
          (sfifo_rescmd_pop && !sfifo_rescmd_not_empty),
          (sfifo_rescmd_full && !sfifo_rescmd_not_empty)};

  // gencmd fifo
  prim_fifo_sync #(
    .Width(GencmdFifoWidth),
    .Pass(0),
    .Depth(GencmdFifoDepth)
  ) u_prim_fifo_sync_gencmd (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (sfifo_gencmd_clr),
    .wvalid_i (sfifo_gencmd_push),
    .wready_o (),
    .wdata_i  (sfifo_gencmd_wdata),
    .rvalid_o (sfifo_gencmd_not_empty),
    .rready_i (sfifo_gencmd_pop),
    .rdata_o  (sfifo_gencmd_rdata),
    .full_o   (sfifo_gencmd_full),
    .depth_o  (sfifo_gencmd_depth),
    .err_o    ()
  );

  // feedback cmd back into gencmd fifo
  assign send_gencmd_d = send_gencmd;

  assign sfifo_gencmd_push =
         (boot_wr_cmd_genfifo & edn_enable_fo[SendGenCmd]) ? 1'b1 :
         (send_gencmd_q & edn_enable_fo[SendGenCmd]) ? 1'b1  :
         generate_cmd_load;

  assign sfifo_gencmd_wdata =
         boot_wr_cmd_genfifo ? boot_gen_cmd :
         auto_req_mode_busy ? cs_cmd_req_out_q :
         generate_cmd_bus;

  assign sfifo_gencmd_pop = send_gencmd || boot_send_gencmd;

  assign sfifo_gencmd_clr = (cmd_fifo_rst_fo[2] || main_sm_done_pulse);

  assign sfifo_gencmd_err =
         {(sfifo_gencmd_push && sfifo_gencmd_full),
          (sfifo_gencmd_pop && !sfifo_gencmd_not_empty),
          (sfifo_gencmd_full && !sfifo_gencmd_not_empty)};

  // output fifo
  prim_fifo_sync #(
    .Width(OutputFifoWidth),
    .Pass(0),
    .Depth(OutputFifoDepth)
  ) u_prim_fifo_sync_output (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (sfifo_output_clr),
    .wvalid_i (sfifo_output_push),
    .wready_o (),
    .wdata_i  (sfifo_output_wdata),
    .rvalid_o (sfifo_output_not_empty),
    .rready_i (sfifo_output_pop),
    .rdata_o  (sfifo_output_rdata),
    .full_o   (sfifo_output_full),
    .depth_o  (),
    .err_o    ()
  );

  // drive outputs
  assign csrng_cmd_o.csrng_req_valid = sfifo_output_not_empty;
  assign csrng_cmd_o.csrng_req_bus = sfifo_output_rdata;

  assign sfifo_output_clr = !edn_enable_fo[OutputClr];
  assign sfifo_output_push = cs_cmd_req_vld_out_q;
  assign sfifo_output_wdata = cs_cmd_req_out_q;
  assign sfifo_output_pop = sfifo_output_not_empty && csrng_cmd_i.csrng_req_ready;

  assign sfifo_output_err =
         {(sfifo_output_push && sfifo_output_full),
          (sfifo_output_pop && !sfifo_output_not_empty),
          (sfifo_output_full && !sfifo_output_not_empty)};

  // sm to process csrng commands
  // SEC_CM: MAIN_SM.FSM.SPARSE
  // SEC_CM: MAIN_SM.CTR.LOCAL_ESC
  edn_main_sm u_edn_main_sm (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .edn_enable_i           (edn_enable_fo[MainFsmEn]),
    .boot_req_mode_i        (boot_req_mode_fo[1]),
    .auto_req_mode_i        (auto_req_mode_pfe),
    .sw_cmd_req_load_i      (sw_cmd_req_load),
    .sw_cmd_valid_o         (sw_cmd_valid),
    .boot_wr_cmd_reg_o      (boot_wr_cmd_reg),
    .boot_wr_cmd_genfifo_o  (boot_wr_cmd_genfifo),
    .auto_set_intr_gate_o   (auto_set_intr_gate),
    .auto_clr_intr_gate_o   (auto_clr_intr_gate),
    .auto_first_ack_wait_o  (auto_first_ack_wait),
    .main_sm_done_pulse_o   (main_sm_done_pulse),
    .csrng_cmd_ack_i        (csrng_cmd_ack),
    .capt_gencmd_fifo_cnt_o (capt_gencmd_fifo_cnt),
    .boot_send_gencmd_o     (boot_send_gencmd),
    .send_gencmd_o          (send_gencmd),
    .max_reqs_cnt_zero_i    (max_reqs_cnt_zero),
    .capt_rescmd_fifo_cnt_o (capt_rescmd_fifo_cnt),
    .send_rescmd_o          (send_rescmd),
    .cmd_sent_i             (cmd_sent),
    .local_escalate_i       (fatal_loc_events),
    .auto_req_mode_busy_o   (auto_req_mode_busy),
    .main_sm_busy_o         (main_sm_busy),
    .main_sm_state_o        (edn_main_sm_state),
    .main_sm_err_o          (edn_main_sm_err)
  );


  // Maximum requests counter for a generate command

  // SEC_CM: CTR.REDUN
  prim_count #(
    .Width(RegWidth),
    .ResetValue({RegWidth{1'b1}})
  ) u_prim_count_max_reqs_cntr (
    .clk_i,
    .rst_ni,
    .clr_i(1'b0),
    .set_i(max_reqs_cnt_load),
    .set_cnt_i(max_reqs_between_reseed_bus),
    .incr_en_i(1'b0),
    .decr_en_i(send_gencmd && cmd_sent), // count down
    .step_i(RegWidth'(1)),
    .cnt_o(max_reqs_cnt),
    .cnt_next_o(),
    .err_o(max_reqs_cnt_err)
  );


  assign max_reqs_cnt_load = (max_reqs_between_reseed_load || // sw initial load
                              send_rescmd && cmd_sent ||      // runtime decrement
                              main_sm_done_pulse);            // restore when auto mode done

  assign max_reqs_cnt_zero = (max_reqs_cnt == '0);


  assign cmd_fifo_cnt_d =
         (!edn_enable_fo[CmdFifoCnt]) ? '0 :
         (cmd_fifo_rst_fo[3] || main_sm_done_pulse) ? '0 :
         capt_gencmd_fifo_cnt ? (sfifo_gencmd_depth) :
         capt_rescmd_fifo_cnt ? (sfifo_rescmd_depth) :
         (send_gencmd || boot_send_gencmd || send_rescmd)? (cmd_fifo_cnt_q-1) :
         cmd_fifo_cnt_q;

  assign cmd_sent = (cmd_fifo_cnt_q == RescmdFifoIdxWidth'(1));

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_boot_req_mode;
  assign mubi_boot_req_mode = mubi4_t'(reg2hw.ctrl.boot_req_mode.q);
  assign boot_req_mode_pfa = mubi4_test_invalid(mubi_boot_req_mode_fanout[0]);
  assign hw2reg.recov_alert_sts.boot_req_mode_field_alert.de = boot_req_mode_pfa;
  assign hw2reg.recov_alert_sts.boot_req_mode_field_alert.d  = boot_req_mode_pfa;

  for (genvar i = 1; i < BootReqCopies; i = i+1) begin : gen_mubi_boot_copies
    assign boot_req_mode_fo[i] = mubi4_test_true_strict(mubi_boot_req_mode_fanout[i]);
  end : gen_mubi_boot_copies

  prim_mubi4_sync #(
    .NumCopies(BootReqCopies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_boot_req_mode (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_boot_req_mode),
    .mubi_o(mubi_boot_req_mode_fanout)
  );


  //--------------------------------------------
  // packer arbitration
  //--------------------------------------------

  prim_arbiter_ppc #(
    .EnDataPort(0),    // Ignore data port
    .N(NumEndPoints),  // Number of request ports
    .DW(1)  // Data width
  ) u_prim_arbiter_ppc_packer_arb (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .req_chk_i(1'b1),
    .req_i(packer_arb_req), // N number of reqs
    .data_i('{default: 1'b0}),
    .gnt_o(packer_arb_gnt), // N number of gnts
    .idx_o(), //NC
    .valid_o(packer_arb_valid),
    .data_o(), // NC
    .ready_i(packer_arb_ready)
  );

  for (genvar i = 0; i < NumEndPoints; i=i+1) begin : gen_arb
    assign packer_arb_req[i] = !packer_ep_rvalid[i] && edn_i[i].edn_req;
  end

  //--------------------------------------------
  // csrng interface packer
  //--------------------------------------------

  prim_packer_fifo #(
     .InW(CSGenBitsWidth),
     .OutW(CSGenBitsWidth),
     .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_cs (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (packer_cs_clr),
    .wvalid_i   (packer_cs_push),
    .wdata_i    (packer_cs_wdata),
    .wready_o   (packer_cs_wready),
    .rvalid_o   (packer_cs_rvalid),
    .rdata_o    (packer_cs_rdata),
    .rready_i   (packer_cs_rready),
    .depth_o    ()
  );

  assign packer_cs_clr = !edn_enable_fo[CsrngPackerClr];
  assign packer_cs_push = csrng_cmd_i.genbits_valid;
  assign packer_cs_wdata = csrng_cmd_i.genbits_bus;
  assign csrng_cmd_o.genbits_ready = packer_cs_wready;
  assign packer_cs_rready = packer_arb_valid;
  assign packer_arb_ready = packer_cs_rvalid;

  assign csrng_fips_d =
         !edn_enable_fo[CsrngFipsEn] ? 1'b0 :
         (packer_cs_push && packer_cs_wready) ? csrng_cmd_i.genbits_fips :
         csrng_fips_q;

  //--------------------------------------------
  // data path integrity check
  // - a counter measure to software genbits bus tampering
  // - checks to make sure repeated data sets off
  //   an alert for sw to handle
  //--------------------------------------------

  // SEC_CM: CS_RDATA.BUS.CONSISTENCY

  // capture a copy of the entropy data
  assign cs_rdata_capt_vld = (packer_cs_rvalid && packer_cs_rready);

  assign cs_rdata_capt_d = cs_rdata_capt_vld ? packer_cs_rdata[63:0] : cs_rdata_capt_q;

  assign cs_rdata_capt_vld_d =
         !edn_enable_fo[CsrngDataVld] ? 1'b0 :
         cs_rdata_capt_vld ? 1'b1 :
         cs_rdata_capt_vld_q;

  // continuous compare of the entropy data
  assign edn_bus_cmp_alert = cs_rdata_capt_vld && cs_rdata_capt_vld_q &&
         (cs_rdata_capt_q == packer_cs_rdata[63:0]);



  prim_edge_detector #(
    .Width(1),
    .ResetValue(0),
    .EnSync(0)
  ) u_prim_edge_detector_recov_alert (
    .clk_i,
    .rst_ni,
    .d_i(edn_bus_cmp_alert),
    .q_sync_o(),
    .q_posedge_pulse_o(recov_alert_o),
    .q_negedge_pulse_o()
  );

  assign hw2reg.recov_alert_sts.edn_bus_cmp_alert.de = edn_bus_cmp_alert;
  assign hw2reg.recov_alert_sts.edn_bus_cmp_alert.d  = edn_bus_cmp_alert;

  //--------------------------------------------
  // end point interface packers generation
  //--------------------------------------------

  for (genvar i = 0; i < NumEndPoints; i=i+1) begin : gen_ep_blk
    prim_packer_fifo #(
      .InW(CSGenBitsWidth),
      .OutW(EndPointBusWidth),
      .ClearOnRead(1'b0)
    ) u_prim_packer_fifo_ep (
      .clk_i      (clk_i),
      .rst_ni     (rst_ni),
      .clr_i      (packer_ep_clr[i]),
      .wvalid_i   (packer_ep_push[i]),
      .wdata_i    (packer_ep_wdata[i]),
      .wready_o   (packer_ep_wready[i]),
      .rvalid_o   (packer_ep_rvalid[i]),
      .rdata_o    (packer_ep_rdata[i]),
      .rready_i   (packer_ep_rready[i]),
      .depth_o    ()
    );

    assign packer_ep_push[i] = packer_arb_valid && packer_ep_wready[i] && packer_arb_gnt[i];
    assign packer_ep_wdata[i] = packer_cs_rdata;

    // fips indication
    assign edn_fips_d[i] = packer_ep_clr[i] ? 1'b0 :
           (packer_ep_push[i] && packer_ep_wready[i]) ?  csrng_fips_q :
           edn_fips_q[i];
    assign edn_o[i].edn_fips = edn_fips_q[i];

    // gate returned data
    assign edn_o[i].edn_ack = packer_ep_ack[i];
    assign edn_o[i].edn_bus = packer_ep_rdata[i];

  // SEC_CM: ACK_SM.FSM.SPARSE
    edn_ack_sm u_edn_ack_sm_ep (
      .clk_i            (clk_i),
      .rst_ni           (rst_ni),
      .enable_i         (edn_enable_fo[AckFsmEn]),
      .req_i            (edn_i[i].edn_req),
      .ack_o            (packer_ep_ack[i]),
      .fifo_not_empty_i (packer_ep_rvalid[i]),
      .fifo_pop_o       (packer_ep_rready[i]),
      .fifo_clr_o       (packer_ep_clr[i]),
      .local_escalate_i (fatal_loc_events),
      .ack_sm_err_o     (edn_ack_sm_err[i])
    );

  end

  // state machine status
  assign hw2reg.main_sm_state.de = 1'b1;
  assign hw2reg.main_sm_state.d = edn_main_sm_state;

  //--------------------------------------------
  // unused signals
  //--------------------------------------------

  assign unused_err_code_test_bit = (|err_code_test_bit[19:3]) || (|err_code_test_bit[27:22]);


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: edn top level wrapper file

`include "prim_assert.sv"

module edn
  import edn_pkg::*;
  import edn_reg_pkg::*;
#(
  parameter int NumEndPoints = 8,
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}}
) (
  input logic clk_i,
  input logic rst_ni,

  // Tilelink Bus registers
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // EDN interfaces
  input  edn_req_t [NumEndPoints-1:0] edn_i,
  output edn_rsp_t [NumEndPoints-1:0] edn_o,

  // CSRNG Application Interface
  output  csrng_pkg::csrng_req_t  csrng_cmd_o,
  input   csrng_pkg::csrng_rsp_t  csrng_cmd_i,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // Interrupts
  output logic      intr_edn_cmd_req_done_o,
  output logic      intr_edn_fatal_err_o
);

  edn_reg2hw_t reg2hw;
  edn_hw2reg_t hw2reg;

  logic [NumAlerts-1:0] alert_test;
  logic [NumAlerts-1:0] alert;

  logic [NumAlerts-1:0] intg_err_alert;
  assign intg_err_alert[0] = 1'b0;


  // SEC_CM: CONFIG.REGWEN
  // SEC_CM: TILE_LINK.BUS.INTEGRITY

  edn_reg_top u_reg (
    .clk_i,
    .rst_ni,
    .tl_i,
    .tl_o,
    .reg2hw,
    .hw2reg,
    .intg_err_o(intg_err_alert[1]), // Assign this alert to the fatal alert index.
    .devmode_i(1'b1)
  );

  edn_core #(
    .NumEndPoints(NumEndPoints)
  ) u_edn_core (
    .clk_i,
    .rst_ni,
    .reg2hw,
    .hw2reg,

    .edn_i,
    .edn_o,

    .csrng_cmd_o,
    .csrng_cmd_i,

    // Alerts

    .recov_alert_o(alert[0]),
    .fatal_alert_o(alert[1]),

    .recov_alert_test_o(alert_test[0]),
    .fatal_alert_test_o(alert_test[1]),

    .intr_edn_cmd_req_done_o,
    .intr_edn_fatal_err_o
  );



  ///////////////////////////
  // Alert generation
  ///////////////////////////
  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i)
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i]                 ),
      .alert_req_i   ( alert[i] || intg_err_alert[i] ),
      .alert_ack_o   (                               ),
      .alert_state_o (                               ),
      .alert_rx_i    ( alert_rx_i[i]                 ),
      .alert_tx_o    ( alert_tx_o[i]                 )
    );
  end


  // Assertions

  `ASSERT_KNOWN(TlDValidKnownO_A, tl_o.d_valid)
  `ASSERT_KNOWN(TlAReadyKnownO_A, tl_o.a_ready)

  // Endpoint Asserts
  for (genvar i = 0; i < NumEndPoints; i = i+1) begin : gen_edn_if_asserts
    `ASSERT_KNOWN(EdnEndPointOut_A, edn_o[i])

    // These assertions check that EDN data will be stable from edn_ack until the next EDN request
    // or until next EDN enablement.
    `ASSERT(EdnDataStable_A, $rose(edn_o[i].edn_ack) |=>
            $stable(edn_o[i].edn_bus) throughout edn_i[i].edn_req[->1],
            clk_i, !rst_ni || !u_edn_core.edn_enable_q)

    `ASSERT(EdnDataStableDisable_A, u_edn_core.edn_enable_q == 0 |=> $stable(edn_o[i].edn_bus))

    `ASSERT(EdnFatalAlertNoRsp_A, alert[1] |-> edn_o[i].edn_ack == 0)
  end : gen_edn_if_asserts

  // CSRNG Asserts
  `ASSERT_KNOWN(CsrngAppIfOut_A, csrng_cmd_o)

  // Alerts
  `ASSERT_KNOWN(AlertTxKnownO_A, alert_tx_o)

  // Interrupt Asserts
  `ASSERT_KNOWN(IntrEdnCmdReqDoneKnownO_A, intr_edn_cmd_req_done_o)

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck_A,
    u_edn_core.u_prim_count_max_reqs_cntr,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(MainFsmCheck_A,
    u_edn_core.u_edn_main_sm.u_state_regs,
    alert_tx_o[1])

  for (genvar i = 0; i < NumEndPoints; i = i+1) begin : gen_edn_fsm_asserts
    `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AckFsmCheck_A,
      u_edn_core.gen_ep_blk[i].u_edn_ack_sm_ep.u_state_regs,
      alert_tx_o[1])
  end

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//

package hmac_pkg;

  localparam int MsgFifoDepth = 16;

  localparam int NumRound = 64;   // SHA-224, SHA-256

  typedef logic [31:0] sha_word_t;
  localparam int WordByte = $bits(sha_word_t)/8;

  typedef struct packed {
    sha_word_t           data;
    logic [WordByte-1:0] mask;
  } sha_fifo_t;


  localparam sha_word_t InitHash [8]= '{
    32'h 6a09_e667, 32'h bb67_ae85, 32'h 3c6e_f372, 32'h a54f_f53a,
    32'h 510e_527f, 32'h 9b05_688c, 32'h 1f83_d9ab, 32'h 5be0_cd19
  };

  localparam sha_word_t CubicRootPrime [64] = '{
    32'h 428a_2f98, 32'h 7137_4491, 32'h b5c0_fbcf, 32'h e9b5_dba5,
    32'h 3956_c25b, 32'h 59f1_11f1, 32'h 923f_82a4, 32'h ab1c_5ed5,
    32'h d807_aa98, 32'h 1283_5b01, 32'h 2431_85be, 32'h 550c_7dc3,
    32'h 72be_5d74, 32'h 80de_b1fe, 32'h 9bdc_06a7, 32'h c19b_f174,
    32'h e49b_69c1, 32'h efbe_4786, 32'h 0fc1_9dc6, 32'h 240c_a1cc,
    32'h 2de9_2c6f, 32'h 4a74_84aa, 32'h 5cb0_a9dc, 32'h 76f9_88da,
    32'h 983e_5152, 32'h a831_c66d, 32'h b003_27c8, 32'h bf59_7fc7,
    32'h c6e0_0bf3, 32'h d5a7_9147, 32'h 06ca_6351, 32'h 1429_2967,
    32'h 27b7_0a85, 32'h 2e1b_2138, 32'h 4d2c_6dfc, 32'h 5338_0d13,
    32'h 650a_7354, 32'h 766a_0abb, 32'h 81c2_c92e, 32'h 9272_2c85,
    32'h a2bf_e8a1, 32'h a81a_664b, 32'h c24b_8b70, 32'h c76c_51a3,
    32'h d192_e819, 32'h d699_0624, 32'h f40e_3585, 32'h 106a_a070,
    32'h 19a4_c116, 32'h 1e37_6c08, 32'h 2748_774c, 32'h 34b0_bcb5,
    32'h 391c_0cb3, 32'h 4ed8_aa4a, 32'h 5b9c_ca4f, 32'h 682e_6ff3,
    32'h 748f_82ee, 32'h 78a5_636f, 32'h 84c8_7814, 32'h 8cc7_0208,
    32'h 90be_fffa, 32'h a450_6ceb, 32'h bef9_a3f7, 32'h c671_78f2
  };

  function automatic sha_word_t conv_endian( input logic [31:0] v, input logic swap);
    logic [31:0] conv_data = {<<8{v}};
    // sha_word_t conv_data = {v[7:0], v[15:8], v[23:16], v[31:24]};
    conv_endian = (swap) ? conv_data : v ;
  endfunction : conv_endian

  function automatic sha_word_t rotr( input sha_word_t v , input int amt );
    rotr = (v >> amt) | (v << (32-amt));
  endfunction : rotr

  function automatic sha_word_t shiftr( input sha_word_t v, input int amt );
    shiftr = (v >> amt);
  endfunction : shiftr

  function automatic sha_word_t [7:0] compress( input sha_word_t w, input sha_word_t k,
                                                input sha_word_t [7:0] h_i);
    automatic sha_word_t sigma_0, sigma_1, ch, maj, temp1, temp2;

    sigma_1 = rotr(h_i[4], 6) ^ rotr(h_i[4], 11) ^ rotr(h_i[4], 25);
    ch = (h_i[4] & h_i[5]) ^ (~h_i[4] & h_i[6]);
    temp1 = (h_i[7] + sigma_1 + ch + k + w);
    sigma_0 = rotr(h_i[0], 2) ^ rotr(h_i[0], 13) ^ rotr(h_i[0], 22);
    maj = (h_i[0] & h_i[1]) ^ (h_i[0] & h_i[2]) ^ (h_i[1] & h_i[2]);
    temp2 = (sigma_0 + maj);

    compress[7] = h_i[6];          // h = g
    compress[6] = h_i[5];          // g = f
    compress[5] = h_i[4];          // f = e
    compress[4] = h_i[3] + temp1;  // e = (d + temp1)
    compress[3] = h_i[2];          // d = c
    compress[2] = h_i[1];          // c = b
    compress[1] = h_i[0];          // b = a
    compress[0] = (temp1 + temp2); // a = (temp1 + temp2)
  endfunction : compress

  function automatic sha_word_t calc_w(input sha_word_t w_0,
                                       input sha_word_t w_1,
                                       input sha_word_t w_9,
                                       input sha_word_t w_14);
    automatic sha_word_t sum0, sum1;
    sum0 = rotr(w_1,   7) ^ rotr(w_1,  18) ^ shiftr(w_1,   3);
    sum1 = rotr(w_14, 17) ^ rotr(w_14, 19) ^ shiftr(w_14, 10);
    calc_w = w_0 + sum0 + w_9 + sum1;
  endfunction : calc_w

  typedef enum logic [31:0] {
    NoError                    = 32'h 0000_0000,
    // SwPushMsgWhenShaDisabled is not used in this version. The error code is
    // guarded by the HW. HW drops the message write request if `sha_en` is
    // off. eunchan@ left the error code to not corrupt the code sequence.
    // Need to rename to DeprecatedSwPush...
    //
    // Issue #3022
    SwPushMsgWhenShaDisabled   = 32'h 0000_0001,
    SwHashStartWhenShaDisabled = 32'h 0000_0002,
    SwUpdateSecretKeyInProcess = 32'h 0000_0003,
    SwHashStartWhenActive      = 32'h 0000_0004,
    SwPushMsgWhenDisallowed    = 32'h 0000_0005
  } err_code_e;

endpackage : hmac_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SHA-256 algorithm
//

module sha2 import hmac_pkg::*; (
  input clk_i,
  input rst_ni,

  input            wipe_secret,
  input sha_word_t wipe_v,

  // FIFO read signal
  input             fifo_rvalid,
  input  sha_fifo_t fifo_rdata,
  output logic      fifo_rready,

  // Control signals
  input        sha_en,   // If disabled, it clears internal content.
  input        hash_start,
  input        hash_process,
  output logic hash_done,

  input        [63:0] message_length,   // bits but byte based
  output sha_word_t [7:0] digest,

  output logic idle
);

  localparam int unsigned RoundWidth = $clog2(NumRound);

  logic msg_feed_complete;

  logic      shaf_rready;
  sha_word_t shaf_rdata;
  logic      shaf_rvalid;

  logic [RoundWidth-1:0] round;

  logic      [3:0]  w_index;
  sha_word_t [15:0] w;

  localparam sha_word_t ZeroWord = '0;

  // w, hash, digest update logic control signals
  logic update_w_from_fifo, calculate_next_w;
  logic init_hash, run_hash, complete_one_chunk;
  logic update_digest, clear_digest;

  logic hash_done_next; // to meet the phase with digest value.

  sha_word_t [7:0] hash;    // a,b,c,d,e,f,g,h

  // Fill up w
  always_ff @(posedge clk_i or negedge rst_ni) begin : fill_w
    if (!rst_ni) begin
      w <= '0;
    end else if (wipe_secret) begin
      w <= w ^ {16{wipe_v}};
    end else if (!sha_en) begin
      w <= '0;
    end else if (!run_hash && update_w_from_fifo) begin
      // this logic runs at the first stage of SHA.
      w <= {shaf_rdata, w[15:1]};
    end else if (calculate_next_w) begin
      w <= {calc_w(w[0], w[1], w[9], w[14]), w[15:1]};
    //end else if (run_hash && update_w_from_fifo) begin
    //  // This code runs when round is in [48, 63]. At this time, it reads from the fifo
    //  // to fill the register if available. If FIFO goes to empty, w_index doesn't increase
    //  // and it cannot reach 15. Then the sha engine doesn't start, which introduces latency.
    //  //
    //  // But in this case, still w should be shifted to feed SHA compress engine. Then
    //  // fifo_rdata should be inserted in the middle of w index.
    //  // w[64-round + w_index] <= fifo_rdata;
    //  for (int i = 0 ; i < 16 ; i++) begin
    //    if (i == (64 - round + w_index)) begin
    //      w[i] <= shaf_rdata;
    //    end else if (i == 15) begin
    //      w[i] <= '0;
    //    end else begin
    //      w[i] <= w[i+1];
    //    end
    //  end
    end else if (run_hash) begin
      // Just shift-out. There's no incoming data
      w <= {ZeroWord, w[15:1]};
    end
  end : fill_w

  // Update engine
  always_ff @(posedge clk_i or negedge rst_ni) begin : compress_round
    if (!rst_ni) begin
      hash <= '{default:'0};
    end else if (wipe_secret) begin
      for (int i = 0 ; i < 8 ; i++) begin
        hash[i] <= hash[i] ^ wipe_v;
      end
    end else if (init_hash) begin
      hash <= digest;
    end else if (run_hash) begin
      hash <= compress( w[0], CubicRootPrime[round], hash);
    end
  end : compress_round

  // Digest
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      digest <= '{default: '0};
    end else if (wipe_secret) begin
      for (int i = 0 ; i < 8 ; i++) begin
        digest[i] <= digest[i] ^ wipe_v;
      end
    end else if (hash_start) begin
      for (int i = 0 ; i < 8 ; i++) begin
        digest[i] <= InitHash[i];
      end
    end else if (!sha_en || clear_digest) begin
      digest <= '0;
    end else if (update_digest) begin
      for (int i = 0 ; i < 8 ; i++) begin
        digest[i] <= digest[i] + hash[i];
      end
    end
  end

  // round
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      round <= '0;
    end else if (!sha_en) begin
      round <= '0;
    end else if (run_hash) begin
      if (round == RoundWidth'(unsigned'(NumRound-1))) begin
        round <= '0;
      end else begin
        round <= round + 1;
      end
    end
  end

  // w_index
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      w_index <= '0;
    end else if (!sha_en) begin
      w_index <= '0;
    end else if (update_w_from_fifo) begin
      w_index <= w_index + 1;
    end
  end

  assign shaf_rready = update_w_from_fifo;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) hash_done <= 1'b0;
    else         hash_done <= hash_done_next;
  end

  typedef enum logic [1:0] {
    FifoIdle,
    FifoLoadFromFifo,
    FifoWait
  } fifoctl_state_e;

  fifoctl_state_e fifo_st_q, fifo_st_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      fifo_st_q <= FifoIdle;
    end else begin
      fifo_st_q <= fifo_st_d;
    end
  end

  always_comb begin
    fifo_st_d = FifoIdle;
    update_w_from_fifo = 1'b0;
    hash_done_next = 1'b0;

    unique case (fifo_st_q)
      FifoIdle: begin
        if (hash_start) begin
          fifo_st_d = FifoLoadFromFifo;
        end else begin
          fifo_st_d = FifoIdle;
        end
      end

      FifoLoadFromFifo: begin
        if (!sha_en) begin
          fifo_st_d = FifoIdle;
          update_w_from_fifo = 1'b0;
        end else if (!shaf_rvalid) begin
          // Wait until it is filled
          fifo_st_d = FifoLoadFromFifo;
          update_w_from_fifo = 1'b0;
        end else if (w_index == 4'd 15) begin
          fifo_st_d = FifoWait;
          update_w_from_fifo = 1'b1;
        end else begin
          fifo_st_d = FifoLoadFromFifo;
          update_w_from_fifo = 1'b1;
        end
      end

      FifoWait: begin
        // Wait until next fetch begins (begin at round == 48)a
        if (msg_feed_complete && complete_one_chunk) begin
          fifo_st_d = FifoIdle;

          hash_done_next = 1'b1;
        end else if (complete_one_chunk) begin
          fifo_st_d = FifoLoadFromFifo;
        end else begin
          fifo_st_d = FifoWait;
        end
      end

      default: begin
        fifo_st_d = FifoIdle;
      end
    endcase
  end

  // SHA control
  typedef enum logic [1:0] {
    ShaIdle,
    ShaCompress,
    ShaUpdateDigest
  } sha_st_t;

  sha_st_t sha_st_q, sha_st_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      sha_st_q <= ShaIdle;
    end else begin
      sha_st_q <= sha_st_d;
    end
  end

  assign clear_digest = hash_start;

  always_comb begin
    update_digest    = 1'b0;
    calculate_next_w = 1'b0;

    init_hash        = 1'b0;
    run_hash         = 1'b0;

    unique case (sha_st_q)
      ShaIdle: begin
        if (fifo_st_q == FifoWait) begin
          init_hash = 1'b1;
          sha_st_d = ShaCompress;
        end else begin
          sha_st_d = ShaIdle;
        end
      end

      ShaCompress: begin
        run_hash = 1'b1;

        if (round < 48) begin
          calculate_next_w = 1'b1;
        end

        if (complete_one_chunk) begin
          sha_st_d = ShaUpdateDigest;
        end else begin
          sha_st_d = ShaCompress;
        end
      end

      ShaUpdateDigest: begin
        update_digest = 1'b1;
        if (fifo_st_q == FifoWait) begin
          init_hash = 1'b1;
          sha_st_d = ShaCompress;
        end else begin
          sha_st_d = ShaIdle;
        end
      end

      default: begin
        sha_st_d = ShaIdle;
      end
    endcase
  end

  // complete_one_chunk
  assign complete_one_chunk = (round == 6'd63);

  sha2_pad u_pad (
    .clk_i,
    .rst_ni,

    .wipe_secret,
    .wipe_v,

    .fifo_rvalid,
    .fifo_rdata,
    .fifo_rready,

    .shaf_rvalid,
    .shaf_rdata,
    .shaf_rready,

    .sha_en,
    .hash_start,
    .hash_process,
    .hash_done,

    .message_length,
    .msg_feed_complete
  );

  // Idle
  assign idle = (fifo_st_q == FifoIdle) && (sha_st_q == ShaIdle) && !hash_start;

endmodule : sha2


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SHA-256 Padding logic
//

`include "prim_assert.sv"

module sha2_pad import hmac_pkg::*; (
  input clk_i,
  input rst_ni,

  input            wipe_secret,
  input sha_word_t wipe_v,

  // To actual FIFO
  input                 fifo_rvalid,
  input  sha_fifo_t     fifo_rdata,
  output logic          fifo_rready,

  // from SHA2 compress engine
  output logic          shaf_rvalid,
  output sha_word_t     shaf_rdata,
  input                 shaf_rready,

  input sha_en,
  input hash_start,
  input hash_process,
  input hash_done,

  input        [63:0] message_length, // # of bytes in bits (8 bits granularity)
  output logic        msg_feed_complete // Indicates, all message is feeded
);

  //logic [8:0] length_added;

  logic [63:0] tx_count;    // fin received data count.

  logic inc_txcount;
  logic fifo_partial;
  logic txcnt_eq_1a0;
  logic hash_process_flag; // Set by hash_process, clear by hash_done

  assign fifo_partial = ~&fifo_rdata.mask;

  // tx_count[8:0] == 'h1c0 --> should send LenHi
  assign txcnt_eq_1a0 = (tx_count[8:0] == 9'h1a0);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      hash_process_flag <= 1'b0;
    end else if (hash_process) begin
      hash_process_flag <= 1'b1;
    end else if (hash_done || hash_start) begin
      hash_process_flag <= 1'b0;
    end
  end

  // Data path: fout_wdata
  typedef enum logic [2:0] {
    FifoIn,         // fin_wdata, fin_wstrb
    Pad80,          // {8'h80, 8'h00} , strb (calc based on len[4:3])
    Pad00,          // 32'h0, full strb
    LenHi,          // len[63:32], full strb
    LenLo           // len[31:0], full strb
  } sel_data_e;
  sel_data_e sel_data;

  always_comb begin
    unique case (sel_data)
      FifoIn: begin
        shaf_rdata = fifo_rdata.data;
      end

      Pad80: begin
        // {a[7:0], b[7:0], c[7:0], d[7:0]}
        // msglen[4:3] == 00 |-> {'h80, 'h00, 'h00, 'h00}
        // msglen[4:3] == 01 |-> {msg,  'h80, 'h00, 'h00}
        // msglen[4:3] == 10 |-> {msg[15:0],  'h80, 'h00}
        // msglen[4:3] == 11 |-> {msg[23:0],        'h80}
        unique case (message_length[4:3])
          2'b 00: shaf_rdata = 32'h 8000_0000;
          2'b 01: shaf_rdata = {fifo_rdata.data[31:24], 24'h 8000_00};
          2'b 10: shaf_rdata = {fifo_rdata.data[31:16], 16'h 8000};
          2'b 11: shaf_rdata = {fifo_rdata.data[31: 8],  8'h 80};
          default: shaf_rdata = 32'h0;
        endcase
      end

      Pad00: begin
        shaf_rdata = '0;
      end

      LenHi: begin
        shaf_rdata = message_length[63:32];
      end

      LenLo: begin
        shaf_rdata = message_length[31:0];
      end

      default: begin
        shaf_rdata = '0;
      end
    endcase
  end

  // Padded length
  // $ceil(message_length + 8 + 64, 512) -> message_length [8:0] + 440 and ignore carry
  //assign length_added = (message_length[8:0] + 9'h1b8) ;

  // fifo control
  // add 8'h 80 , N 8'h00, 64'h message_length

  // Steps
  // 1. `hash_start` from CPU (or DMA?)
  // 2. calculate `padded_length` from `message_length`
  // 3. Check if tx_count == message_length, then go to 5
  // 4. Receiving FIFO input (hand over to fifo output)
  // 5. Padding bit 1 (8'h80) followed by 8'h00 if needed
  // 6. Padding with length (high -> low)

  // State Machine
  typedef enum logic [2:0] {
    StIdle,        // fin_full to prevent unwanted FIFO write
    StFifoReceive, // Check tx_count == message_length
    StPad80,       // 8'h 80 + 8'h 00 X N
    StPad00,
    StLenHi,
    StLenLo
  } pad_st_e;

  pad_st_e st_q, st_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      st_q <= StIdle;
    end else begin
      st_q <= st_d;
    end
  end

  // Next state
  always_comb begin
    shaf_rvalid = 1'b0;
    inc_txcount = 1'b0;
    sel_data = FifoIn;
    fifo_rready = 1'b0;

    st_d = StIdle;

    unique case (st_q)
      StIdle: begin
        sel_data = FifoIn;
        shaf_rvalid = 1'b0;

        if (sha_en && hash_start) begin
          inc_txcount = 1'b0;

          st_d = StFifoReceive;
        end else begin
          st_d = StIdle;
        end
      end

      StFifoReceive: begin
        sel_data = FifoIn;

        if (fifo_partial && fifo_rvalid) begin
          // End of the message, assume hash_process_flag is set
          shaf_rvalid  = 1'b0; // Update entry at StPad80
          inc_txcount = 1'b0;
          fifo_rready = 1'b0;

          st_d = StPad80;
        end else if (!hash_process_flag) begin
          fifo_rready = shaf_rready;
          shaf_rvalid  = fifo_rvalid;
          inc_txcount = shaf_rready;

          st_d = StFifoReceive;
        end else if (tx_count == message_length) begin
          // already received all msg and was waiting process flag
          shaf_rvalid  = 1'b0;
          inc_txcount = 1'b0;
          fifo_rready = 1'b0;

          st_d = StPad80;
        end else begin
          shaf_rvalid  = fifo_rvalid;
          fifo_rready = shaf_rready; // 0 always
          inc_txcount = shaf_rready; // 0 always

          st_d = StFifoReceive;
        end
      end

      StPad80: begin
        sel_data = Pad80;

        shaf_rvalid = 1'b1;
        fifo_rready = shaf_rready && |message_length[4:3]; // Only when partial

        // exactly 96 bits left, do not need to pad00's
        if (shaf_rready && txcnt_eq_1a0) begin
          st_d = StLenHi;
          inc_txcount = 1'b1;
        // it does not matter if value is < or > than 416 bits.  If it's the former, 00 pad until
        // length field.  If >, then the next chunk will contain the length field with appropriate
        // 0 padding.
        end else if (shaf_rready && !txcnt_eq_1a0) begin
          st_d = StPad00;
          inc_txcount = 1'b1;
        end else begin
          st_d = StPad80;
          inc_txcount = 1'b0;
        end

        // # Below part is temporal code to speed up the SHA by 16 clocks per chunk
        // # (80 clk --> 64 clk)
        // # leaving this as a reference but needs to verify it.
        //if (shaf_rready && !txcnt_eq_1a0) begin
        //  st_d = StPad00;
        //
        //  inc_txcount = 1'b1;
        //  shaf_rvalid = (msg_word_aligned) ? 1'b1 : fifo_rvalid;
        //  fifo_rready = (msg_word_aligned) ? 1'b0 : 1'b1;
        //end else if (!shaf_rready && !txcnt_eq_1a0) begin
        //  st_d = StPad80;
        //
        //  inc_txcount = 1'b0;
        //  shaf_rvalid = (msg_word_aligned) ? 1'b1 : fifo_rvalid;
        //
        //end else if (shaf_rready && txcnt_eq_1a0) begin
        //  st_d = StLenHi;
        //  inc_txcount = 1'b1;
        //end else begin
        //  // !shaf_rready && txcnt_eq_1a0 , just wait until fifo_rready asserted
        //  st_d = StPad80;
        //  inc_txcount = 1'b0;
        //end
      end

      StPad00: begin
        sel_data = Pad00;
        shaf_rvalid = 1'b1;

        if (shaf_rready) begin
          inc_txcount = 1'b1;

          if (txcnt_eq_1a0) begin
            st_d = StLenHi;
          end else begin
            st_d = StPad00;
          end
        end else begin
          st_d = StPad00;
        end
      end

      StLenHi: begin
        sel_data = LenHi;
        shaf_rvalid = 1'b1;

        if (shaf_rready) begin
          st_d = StLenLo;

          inc_txcount = 1'b1;
        end else begin
          st_d = StLenHi;

          inc_txcount = 1'b0;
        end
      end

      StLenLo: begin
        sel_data = LenLo;
        shaf_rvalid = 1'b1;

        if (shaf_rready) begin
          st_d = StIdle;

          inc_txcount = 1'b1;
        end else begin
          st_d = StLenLo;

          inc_txcount = 1'b0;
        end
      end

      default: begin
        st_d = StIdle;
      end
    endcase
  end

  // tx_count
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      tx_count <= '0;
    end else if (hash_start) begin
      tx_count <= '0;
    end else if (inc_txcount) begin
      tx_count[63:5] <= tx_count[63:5] + 1'b1;
    end
  end

  // State machine is in Idle only when it meets tx_count == message length
  assign msg_feed_complete = hash_process_flag && (st_q == StIdle);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package hmac_reg_pkg;

  // Param list
  parameter int NumWords = 8;
  parameter int NumAlerts = 1;

  // Address widths within the block
  parameter int BlockAw = 12;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } hmac_done;
    struct packed {
      logic        q;
    } fifo_empty;
    struct packed {
      logic        q;
    } hmac_err;
  } hmac_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } hmac_done;
    struct packed {
      logic        q;
    } fifo_empty;
    struct packed {
      logic        q;
    } hmac_err;
  } hmac_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } hmac_done;
    struct packed {
      logic        q;
      logic        qe;
    } fifo_empty;
    struct packed {
      logic        q;
      logic        qe;
    } hmac_err;
  } hmac_reg2hw_intr_test_reg_t;

  typedef struct packed {
    logic        q;
    logic        qe;
  } hmac_reg2hw_alert_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } hmac_en;
    struct packed {
      logic        q;
      logic        qe;
    } sha_en;
    struct packed {
      logic        q;
      logic        qe;
    } endian_swap;
    struct packed {
      logic        q;
      logic        qe;
    } digest_swap;
  } hmac_reg2hw_cfg_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } hash_start;
    struct packed {
      logic        q;
      logic        qe;
    } hash_process;
  } hmac_reg2hw_cmd_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } hmac_reg2hw_wipe_secret_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } hmac_reg2hw_key_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } hmac_done;
    struct packed {
      logic        d;
      logic        de;
    } fifo_empty;
    struct packed {
      logic        d;
      logic        de;
    } hmac_err;
  } hmac_hw2reg_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } hmac_en;
    struct packed {
      logic        d;
    } sha_en;
    struct packed {
      logic        d;
    } endian_swap;
    struct packed {
      logic        d;
    } digest_swap;
  } hmac_hw2reg_cfg_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } fifo_empty;
    struct packed {
      logic        d;
    } fifo_full;
    struct packed {
      logic [4:0]  d;
    } fifo_depth;
  } hmac_hw2reg_status_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } hmac_hw2reg_err_code_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } hmac_hw2reg_key_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } hmac_hw2reg_digest_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } hmac_hw2reg_msg_length_lower_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } hmac_hw2reg_msg_length_upper_reg_t;

  // Register -> HW type
  typedef struct packed {
    hmac_reg2hw_intr_state_reg_t intr_state; // [322:320]
    hmac_reg2hw_intr_enable_reg_t intr_enable; // [319:317]
    hmac_reg2hw_intr_test_reg_t intr_test; // [316:311]
    hmac_reg2hw_alert_test_reg_t alert_test; // [310:309]
    hmac_reg2hw_cfg_reg_t cfg; // [308:301]
    hmac_reg2hw_cmd_reg_t cmd; // [300:297]
    hmac_reg2hw_wipe_secret_reg_t wipe_secret; // [296:264]
    hmac_reg2hw_key_mreg_t [7:0] key; // [263:0]
  } hmac_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    hmac_hw2reg_intr_state_reg_t intr_state; // [627:622]
    hmac_hw2reg_cfg_reg_t cfg; // [621:618]
    hmac_hw2reg_status_reg_t status; // [617:611]
    hmac_hw2reg_err_code_reg_t err_code; // [610:578]
    hmac_hw2reg_key_mreg_t [7:0] key; // [577:322]
    hmac_hw2reg_digest_mreg_t [7:0] digest; // [321:66]
    hmac_hw2reg_msg_length_lower_reg_t msg_length_lower; // [65:33]
    hmac_hw2reg_msg_length_upper_reg_t msg_length_upper; // [32:0]
  } hmac_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] HMAC_INTR_STATE_OFFSET = 12'h 0;
  parameter logic [BlockAw-1:0] HMAC_INTR_ENABLE_OFFSET = 12'h 4;
  parameter logic [BlockAw-1:0] HMAC_INTR_TEST_OFFSET = 12'h 8;
  parameter logic [BlockAw-1:0] HMAC_ALERT_TEST_OFFSET = 12'h c;
  parameter logic [BlockAw-1:0] HMAC_CFG_OFFSET = 12'h 10;
  parameter logic [BlockAw-1:0] HMAC_CMD_OFFSET = 12'h 14;
  parameter logic [BlockAw-1:0] HMAC_STATUS_OFFSET = 12'h 18;
  parameter logic [BlockAw-1:0] HMAC_ERR_CODE_OFFSET = 12'h 1c;
  parameter logic [BlockAw-1:0] HMAC_WIPE_SECRET_OFFSET = 12'h 20;
  parameter logic [BlockAw-1:0] HMAC_KEY_0_OFFSET = 12'h 24;
  parameter logic [BlockAw-1:0] HMAC_KEY_1_OFFSET = 12'h 28;
  parameter logic [BlockAw-1:0] HMAC_KEY_2_OFFSET = 12'h 2c;
  parameter logic [BlockAw-1:0] HMAC_KEY_3_OFFSET = 12'h 30;
  parameter logic [BlockAw-1:0] HMAC_KEY_4_OFFSET = 12'h 34;
  parameter logic [BlockAw-1:0] HMAC_KEY_5_OFFSET = 12'h 38;
  parameter logic [BlockAw-1:0] HMAC_KEY_6_OFFSET = 12'h 3c;
  parameter logic [BlockAw-1:0] HMAC_KEY_7_OFFSET = 12'h 40;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_0_OFFSET = 12'h 44;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_1_OFFSET = 12'h 48;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_2_OFFSET = 12'h 4c;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_3_OFFSET = 12'h 50;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_4_OFFSET = 12'h 54;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_5_OFFSET = 12'h 58;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_6_OFFSET = 12'h 5c;
  parameter logic [BlockAw-1:0] HMAC_DIGEST_7_OFFSET = 12'h 60;
  parameter logic [BlockAw-1:0] HMAC_MSG_LENGTH_LOWER_OFFSET = 12'h 64;
  parameter logic [BlockAw-1:0] HMAC_MSG_LENGTH_UPPER_OFFSET = 12'h 68;

  // Reset values for hwext registers and their fields
  parameter logic [2:0] HMAC_INTR_TEST_RESVAL = 3'h 0;
  parameter logic [0:0] HMAC_INTR_TEST_HMAC_DONE_RESVAL = 1'h 0;
  parameter logic [0:0] HMAC_INTR_TEST_FIFO_EMPTY_RESVAL = 1'h 0;
  parameter logic [0:0] HMAC_INTR_TEST_HMAC_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] HMAC_ALERT_TEST_RESVAL = 1'h 0;
  parameter logic [0:0] HMAC_ALERT_TEST_FATAL_FAULT_RESVAL = 1'h 0;
  parameter logic [3:0] HMAC_CFG_RESVAL = 4'h 0;
  parameter logic [0:0] HMAC_CFG_ENDIAN_SWAP_RESVAL = 1'h 0;
  parameter logic [0:0] HMAC_CFG_DIGEST_SWAP_RESVAL = 1'h 0;
  parameter logic [1:0] HMAC_CMD_RESVAL = 2'h 0;
  parameter logic [8:0] HMAC_STATUS_RESVAL = 9'h 1;
  parameter logic [0:0] HMAC_STATUS_FIFO_EMPTY_RESVAL = 1'h 1;
  parameter logic [31:0] HMAC_WIPE_SECRET_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_0_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_1_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_2_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_3_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_4_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_5_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_6_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_KEY_7_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_0_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_1_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_2_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_3_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_4_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_5_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_6_RESVAL = 32'h 0;
  parameter logic [31:0] HMAC_DIGEST_7_RESVAL = 32'h 0;

  // Window parameters
  parameter logic [BlockAw-1:0] HMAC_MSG_FIFO_OFFSET = 12'h 800;
  parameter int unsigned        HMAC_MSG_FIFO_SIZE   = 'h 800;

  // Register index
  typedef enum int {
    HMAC_INTR_STATE,
    HMAC_INTR_ENABLE,
    HMAC_INTR_TEST,
    HMAC_ALERT_TEST,
    HMAC_CFG,
    HMAC_CMD,
    HMAC_STATUS,
    HMAC_ERR_CODE,
    HMAC_WIPE_SECRET,
    HMAC_KEY_0,
    HMAC_KEY_1,
    HMAC_KEY_2,
    HMAC_KEY_3,
    HMAC_KEY_4,
    HMAC_KEY_5,
    HMAC_KEY_6,
    HMAC_KEY_7,
    HMAC_DIGEST_0,
    HMAC_DIGEST_1,
    HMAC_DIGEST_2,
    HMAC_DIGEST_3,
    HMAC_DIGEST_4,
    HMAC_DIGEST_5,
    HMAC_DIGEST_6,
    HMAC_DIGEST_7,
    HMAC_MSG_LENGTH_LOWER,
    HMAC_MSG_LENGTH_UPPER
  } hmac_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] HMAC_PERMIT [27] = '{
    4'b 0001, // index[ 0] HMAC_INTR_STATE
    4'b 0001, // index[ 1] HMAC_INTR_ENABLE
    4'b 0001, // index[ 2] HMAC_INTR_TEST
    4'b 0001, // index[ 3] HMAC_ALERT_TEST
    4'b 0001, // index[ 4] HMAC_CFG
    4'b 0001, // index[ 5] HMAC_CMD
    4'b 0011, // index[ 6] HMAC_STATUS
    4'b 1111, // index[ 7] HMAC_ERR_CODE
    4'b 1111, // index[ 8] HMAC_WIPE_SECRET
    4'b 1111, // index[ 9] HMAC_KEY_0
    4'b 1111, // index[10] HMAC_KEY_1
    4'b 1111, // index[11] HMAC_KEY_2
    4'b 1111, // index[12] HMAC_KEY_3
    4'b 1111, // index[13] HMAC_KEY_4
    4'b 1111, // index[14] HMAC_KEY_5
    4'b 1111, // index[15] HMAC_KEY_6
    4'b 1111, // index[16] HMAC_KEY_7
    4'b 1111, // index[17] HMAC_DIGEST_0
    4'b 1111, // index[18] HMAC_DIGEST_1
    4'b 1111, // index[19] HMAC_DIGEST_2
    4'b 1111, // index[20] HMAC_DIGEST_3
    4'b 1111, // index[21] HMAC_DIGEST_4
    4'b 1111, // index[22] HMAC_DIGEST_5
    4'b 1111, // index[23] HMAC_DIGEST_6
    4'b 1111, // index[24] HMAC_DIGEST_7
    4'b 1111, // index[25] HMAC_MSG_LENGTH_LOWER
    4'b 1111  // index[26] HMAC_MSG_LENGTH_UPPER
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module hmac_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // Output port for window
  output tlul_pkg::tl_h2d_t tl_win_o,
  input  tlul_pkg::tl_d2h_t tl_win_i,

  // To HW
  output hmac_reg_pkg::hmac_reg2hw_t reg2hw, // Write
  input  hmac_reg_pkg::hmac_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import hmac_reg_pkg::* ;

  localparam int AW = 12;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [26:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(27)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  tlul_pkg::tl_h2d_t tl_socket_h2d [2];
  tlul_pkg::tl_d2h_t tl_socket_d2h [2];

  logic [0:0] reg_steer;

  // socket_1n connection
  assign tl_reg_h2d = tl_socket_h2d[1];
  assign tl_socket_d2h[1] = tl_reg_d2h;

  assign tl_win_o = tl_socket_h2d[0];
  assign tl_socket_d2h[0] = tl_win_i;

  // Create Socket_1n
  tlul_socket_1n #(
    .N            (2),
    .HReqPass     (1'b1),
    .HRspPass     (1'b1),
    .DReqPass     ({2{1'b1}}),
    .DRspPass     ({2{1'b1}}),
    .HReqDepth    (4'h0),
    .HRspDepth    (4'h0),
    .DReqDepth    ({2{4'h0}}),
    .DRspDepth    ({2{4'h0}}),
    .ExplicitErrs (1'b0)
  ) u_socket (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),
    .tl_h_i (tl_i),
    .tl_h_o (tl_o_pre),
    .tl_d_o (tl_socket_h2d),
    .tl_d_i (tl_socket_d2h),
    .dev_select_i (reg_steer)
  );

  // Create steering logic
  always_comb begin
    reg_steer =
        tl_i.a_address[AW-1:0] inside {[2048:4095]} ? 1'd0 :
        // Default set to register
        1'd1;

    // Override this in case of an integrity error
    if (intg_err) begin
      reg_steer = 1'd1;
    end
  end

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_hmac_done_qs;
  logic intr_state_hmac_done_wd;
  logic intr_state_fifo_empty_qs;
  logic intr_state_fifo_empty_wd;
  logic intr_state_hmac_err_qs;
  logic intr_state_hmac_err_wd;
  logic intr_enable_we;
  logic intr_enable_hmac_done_qs;
  logic intr_enable_hmac_done_wd;
  logic intr_enable_fifo_empty_qs;
  logic intr_enable_fifo_empty_wd;
  logic intr_enable_hmac_err_qs;
  logic intr_enable_hmac_err_wd;
  logic intr_test_we;
  logic intr_test_hmac_done_wd;
  logic intr_test_fifo_empty_wd;
  logic intr_test_hmac_err_wd;
  logic alert_test_we;
  logic alert_test_wd;
  logic cfg_re;
  logic cfg_we;
  logic cfg_hmac_en_qs;
  logic cfg_hmac_en_wd;
  logic cfg_sha_en_qs;
  logic cfg_sha_en_wd;
  logic cfg_endian_swap_qs;
  logic cfg_endian_swap_wd;
  logic cfg_digest_swap_qs;
  logic cfg_digest_swap_wd;
  logic cmd_we;
  logic cmd_hash_start_wd;
  logic cmd_hash_process_wd;
  logic status_re;
  logic status_fifo_empty_qs;
  logic status_fifo_full_qs;
  logic [4:0] status_fifo_depth_qs;
  logic [31:0] err_code_qs;
  logic wipe_secret_we;
  logic [31:0] wipe_secret_wd;
  logic key_0_we;
  logic [31:0] key_0_wd;
  logic key_1_we;
  logic [31:0] key_1_wd;
  logic key_2_we;
  logic [31:0] key_2_wd;
  logic key_3_we;
  logic [31:0] key_3_wd;
  logic key_4_we;
  logic [31:0] key_4_wd;
  logic key_5_we;
  logic [31:0] key_5_wd;
  logic key_6_we;
  logic [31:0] key_6_wd;
  logic key_7_we;
  logic [31:0] key_7_wd;
  logic digest_0_re;
  logic [31:0] digest_0_qs;
  logic digest_1_re;
  logic [31:0] digest_1_qs;
  logic digest_2_re;
  logic [31:0] digest_2_qs;
  logic digest_3_re;
  logic [31:0] digest_3_qs;
  logic digest_4_re;
  logic [31:0] digest_4_qs;
  logic digest_5_re;
  logic [31:0] digest_5_qs;
  logic digest_6_re;
  logic [31:0] digest_6_qs;
  logic digest_7_re;
  logic [31:0] digest_7_qs;
  logic [31:0] msg_length_lower_qs;
  logic [31:0] msg_length_upper_qs;

  // Register instances
  // R[intr_state]: V(False)
  //   F[hmac_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_hmac_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_hmac_done_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.hmac_done.de),
    .d      (hw2reg.intr_state.hmac_done.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.hmac_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_hmac_done_qs)
  );

  //   F[fifo_empty]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_fifo_empty (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_fifo_empty_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.fifo_empty.de),
    .d      (hw2reg.intr_state.fifo_empty.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.fifo_empty.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_fifo_empty_qs)
  );

  //   F[hmac_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_hmac_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_hmac_err_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.hmac_err.de),
    .d      (hw2reg.intr_state.hmac_err.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.hmac_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_hmac_err_qs)
  );


  // R[intr_enable]: V(False)
  //   F[hmac_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_hmac_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_hmac_done_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.hmac_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_hmac_done_qs)
  );

  //   F[fifo_empty]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_fifo_empty (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_fifo_empty_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.fifo_empty.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_fifo_empty_qs)
  );

  //   F[hmac_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_hmac_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_hmac_err_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.hmac_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_hmac_err_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [2:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  //   F[hmac_done]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_hmac_done (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_hmac_done_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.hmac_done.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.hmac_done.qe = intr_test_qe;

  //   F[fifo_empty]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_fifo_empty (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_fifo_empty_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[1]),
    .q      (reg2hw.intr_test.fifo_empty.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.fifo_empty.qe = intr_test_qe;

  //   F[hmac_err]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_hmac_err (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_hmac_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[2]),
    .q      (reg2hw.intr_test.hmac_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.hmac_err.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [0:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.qe = alert_test_qe;


  // R[cfg]: V(True)
  logic cfg_qe;
  logic [3:0] cfg_flds_we;
  assign cfg_qe = &cfg_flds_we;
  //   F[hmac_en]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_cfg_hmac_en (
    .re     (cfg_re),
    .we     (cfg_we),
    .wd     (cfg_hmac_en_wd),
    .d      (hw2reg.cfg.hmac_en.d),
    .qre    (),
    .qe     (cfg_flds_we[0]),
    .q      (reg2hw.cfg.hmac_en.q),
    .ds     (),
    .qs     (cfg_hmac_en_qs)
  );
  assign reg2hw.cfg.hmac_en.qe = cfg_qe;

  //   F[sha_en]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_cfg_sha_en (
    .re     (cfg_re),
    .we     (cfg_we),
    .wd     (cfg_sha_en_wd),
    .d      (hw2reg.cfg.sha_en.d),
    .qre    (),
    .qe     (cfg_flds_we[1]),
    .q      (reg2hw.cfg.sha_en.q),
    .ds     (),
    .qs     (cfg_sha_en_qs)
  );
  assign reg2hw.cfg.sha_en.qe = cfg_qe;

  //   F[endian_swap]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_cfg_endian_swap (
    .re     (cfg_re),
    .we     (cfg_we),
    .wd     (cfg_endian_swap_wd),
    .d      (hw2reg.cfg.endian_swap.d),
    .qre    (),
    .qe     (cfg_flds_we[2]),
    .q      (reg2hw.cfg.endian_swap.q),
    .ds     (),
    .qs     (cfg_endian_swap_qs)
  );
  assign reg2hw.cfg.endian_swap.qe = cfg_qe;

  //   F[digest_swap]: 3:3
  prim_subreg_ext #(
    .DW    (1)
  ) u_cfg_digest_swap (
    .re     (cfg_re),
    .we     (cfg_we),
    .wd     (cfg_digest_swap_wd),
    .d      (hw2reg.cfg.digest_swap.d),
    .qre    (),
    .qe     (cfg_flds_we[3]),
    .q      (reg2hw.cfg.digest_swap.q),
    .ds     (),
    .qs     (cfg_digest_swap_qs)
  );
  assign reg2hw.cfg.digest_swap.qe = cfg_qe;


  // R[cmd]: V(True)
  logic cmd_qe;
  logic [1:0] cmd_flds_we;
  assign cmd_qe = &cmd_flds_we;
  //   F[hash_start]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_cmd_hash_start (
    .re     (1'b0),
    .we     (cmd_we),
    .wd     (cmd_hash_start_wd),
    .d      ('0),
    .qre    (),
    .qe     (cmd_flds_we[0]),
    .q      (reg2hw.cmd.hash_start.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.cmd.hash_start.qe = cmd_qe;

  //   F[hash_process]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_cmd_hash_process (
    .re     (1'b0),
    .we     (cmd_we),
    .wd     (cmd_hash_process_wd),
    .d      ('0),
    .qre    (),
    .qe     (cmd_flds_we[1]),
    .q      (reg2hw.cmd.hash_process.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.cmd.hash_process.qe = cmd_qe;


  // R[status]: V(True)
  //   F[fifo_empty]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_fifo_empty (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.fifo_empty.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_fifo_empty_qs)
  );

  //   F[fifo_full]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_fifo_full (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.fifo_full.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_fifo_full_qs)
  );

  //   F[fifo_depth]: 8:4
  prim_subreg_ext #(
    .DW    (5)
  ) u_status_fifo_depth (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.fifo_depth.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_fifo_depth_qs)
  );


  // R[err_code]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_err_code (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.de),
    .d      (hw2reg.err_code.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_qs)
  );


  // R[wipe_secret]: V(True)
  logic wipe_secret_qe;
  logic [0:0] wipe_secret_flds_we;
  assign wipe_secret_qe = &wipe_secret_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_wipe_secret (
    .re     (1'b0),
    .we     (wipe_secret_we),
    .wd     (wipe_secret_wd),
    .d      ('0),
    .qre    (),
    .qe     (wipe_secret_flds_we[0]),
    .q      (reg2hw.wipe_secret.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.wipe_secret.qe = wipe_secret_qe;


  // Subregister 0 of Multireg key
  // R[key_0]: V(True)
  logic key_0_qe;
  logic [0:0] key_0_flds_we;
  assign key_0_qe = &key_0_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_0 (
    .re     (1'b0),
    .we     (key_0_we),
    .wd     (key_0_wd),
    .d      (hw2reg.key[0].d),
    .qre    (),
    .qe     (key_0_flds_we[0]),
    .q      (reg2hw.key[0].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[0].qe = key_0_qe;


  // Subregister 1 of Multireg key
  // R[key_1]: V(True)
  logic key_1_qe;
  logic [0:0] key_1_flds_we;
  assign key_1_qe = &key_1_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_1 (
    .re     (1'b0),
    .we     (key_1_we),
    .wd     (key_1_wd),
    .d      (hw2reg.key[1].d),
    .qre    (),
    .qe     (key_1_flds_we[0]),
    .q      (reg2hw.key[1].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[1].qe = key_1_qe;


  // Subregister 2 of Multireg key
  // R[key_2]: V(True)
  logic key_2_qe;
  logic [0:0] key_2_flds_we;
  assign key_2_qe = &key_2_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_2 (
    .re     (1'b0),
    .we     (key_2_we),
    .wd     (key_2_wd),
    .d      (hw2reg.key[2].d),
    .qre    (),
    .qe     (key_2_flds_we[0]),
    .q      (reg2hw.key[2].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[2].qe = key_2_qe;


  // Subregister 3 of Multireg key
  // R[key_3]: V(True)
  logic key_3_qe;
  logic [0:0] key_3_flds_we;
  assign key_3_qe = &key_3_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_3 (
    .re     (1'b0),
    .we     (key_3_we),
    .wd     (key_3_wd),
    .d      (hw2reg.key[3].d),
    .qre    (),
    .qe     (key_3_flds_we[0]),
    .q      (reg2hw.key[3].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[3].qe = key_3_qe;


  // Subregister 4 of Multireg key
  // R[key_4]: V(True)
  logic key_4_qe;
  logic [0:0] key_4_flds_we;
  assign key_4_qe = &key_4_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_4 (
    .re     (1'b0),
    .we     (key_4_we),
    .wd     (key_4_wd),
    .d      (hw2reg.key[4].d),
    .qre    (),
    .qe     (key_4_flds_we[0]),
    .q      (reg2hw.key[4].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[4].qe = key_4_qe;


  // Subregister 5 of Multireg key
  // R[key_5]: V(True)
  logic key_5_qe;
  logic [0:0] key_5_flds_we;
  assign key_5_qe = &key_5_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_5 (
    .re     (1'b0),
    .we     (key_5_we),
    .wd     (key_5_wd),
    .d      (hw2reg.key[5].d),
    .qre    (),
    .qe     (key_5_flds_we[0]),
    .q      (reg2hw.key[5].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[5].qe = key_5_qe;


  // Subregister 6 of Multireg key
  // R[key_6]: V(True)
  logic key_6_qe;
  logic [0:0] key_6_flds_we;
  assign key_6_qe = &key_6_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_6 (
    .re     (1'b0),
    .we     (key_6_we),
    .wd     (key_6_wd),
    .d      (hw2reg.key[6].d),
    .qre    (),
    .qe     (key_6_flds_we[0]),
    .q      (reg2hw.key[6].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[6].qe = key_6_qe;


  // Subregister 7 of Multireg key
  // R[key_7]: V(True)
  logic key_7_qe;
  logic [0:0] key_7_flds_we;
  assign key_7_qe = &key_7_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_7 (
    .re     (1'b0),
    .we     (key_7_we),
    .wd     (key_7_wd),
    .d      (hw2reg.key[7].d),
    .qre    (),
    .qe     (key_7_flds_we[0]),
    .q      (reg2hw.key[7].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key[7].qe = key_7_qe;


  // Subregister 0 of Multireg digest
  // R[digest_0]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_0 (
    .re     (digest_0_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[0].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_0_qs)
  );


  // Subregister 1 of Multireg digest
  // R[digest_1]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_1 (
    .re     (digest_1_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[1].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_1_qs)
  );


  // Subregister 2 of Multireg digest
  // R[digest_2]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_2 (
    .re     (digest_2_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[2].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_2_qs)
  );


  // Subregister 3 of Multireg digest
  // R[digest_3]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_3 (
    .re     (digest_3_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[3].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_3_qs)
  );


  // Subregister 4 of Multireg digest
  // R[digest_4]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_4 (
    .re     (digest_4_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[4].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_4_qs)
  );


  // Subregister 5 of Multireg digest
  // R[digest_5]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_5 (
    .re     (digest_5_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[5].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_5_qs)
  );


  // Subregister 6 of Multireg digest
  // R[digest_6]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_6 (
    .re     (digest_6_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[6].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_6_qs)
  );


  // Subregister 7 of Multireg digest
  // R[digest_7]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_digest_7 (
    .re     (digest_7_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.digest[7].d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (digest_7_qs)
  );


  // R[msg_length_lower]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_msg_length_lower (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.msg_length_lower.de),
    .d      (hw2reg.msg_length_lower.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (msg_length_lower_qs)
  );


  // R[msg_length_upper]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_msg_length_upper (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.msg_length_upper.de),
    .d      (hw2reg.msg_length_upper.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (msg_length_upper_qs)
  );



  logic [26:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == HMAC_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == HMAC_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == HMAC_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == HMAC_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == HMAC_CFG_OFFSET);
    addr_hit[ 5] = (reg_addr == HMAC_CMD_OFFSET);
    addr_hit[ 6] = (reg_addr == HMAC_STATUS_OFFSET);
    addr_hit[ 7] = (reg_addr == HMAC_ERR_CODE_OFFSET);
    addr_hit[ 8] = (reg_addr == HMAC_WIPE_SECRET_OFFSET);
    addr_hit[ 9] = (reg_addr == HMAC_KEY_0_OFFSET);
    addr_hit[10] = (reg_addr == HMAC_KEY_1_OFFSET);
    addr_hit[11] = (reg_addr == HMAC_KEY_2_OFFSET);
    addr_hit[12] = (reg_addr == HMAC_KEY_3_OFFSET);
    addr_hit[13] = (reg_addr == HMAC_KEY_4_OFFSET);
    addr_hit[14] = (reg_addr == HMAC_KEY_5_OFFSET);
    addr_hit[15] = (reg_addr == HMAC_KEY_6_OFFSET);
    addr_hit[16] = (reg_addr == HMAC_KEY_7_OFFSET);
    addr_hit[17] = (reg_addr == HMAC_DIGEST_0_OFFSET);
    addr_hit[18] = (reg_addr == HMAC_DIGEST_1_OFFSET);
    addr_hit[19] = (reg_addr == HMAC_DIGEST_2_OFFSET);
    addr_hit[20] = (reg_addr == HMAC_DIGEST_3_OFFSET);
    addr_hit[21] = (reg_addr == HMAC_DIGEST_4_OFFSET);
    addr_hit[22] = (reg_addr == HMAC_DIGEST_5_OFFSET);
    addr_hit[23] = (reg_addr == HMAC_DIGEST_6_OFFSET);
    addr_hit[24] = (reg_addr == HMAC_DIGEST_7_OFFSET);
    addr_hit[25] = (reg_addr == HMAC_MSG_LENGTH_LOWER_OFFSET);
    addr_hit[26] = (reg_addr == HMAC_MSG_LENGTH_UPPER_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(HMAC_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(HMAC_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(HMAC_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(HMAC_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(HMAC_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(HMAC_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(HMAC_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(HMAC_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(HMAC_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(HMAC_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(HMAC_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(HMAC_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(HMAC_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(HMAC_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(HMAC_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(HMAC_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(HMAC_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(HMAC_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(HMAC_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(HMAC_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(HMAC_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(HMAC_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(HMAC_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(HMAC_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(HMAC_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(HMAC_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(HMAC_PERMIT[26] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_hmac_done_wd = reg_wdata[0];

  assign intr_state_fifo_empty_wd = reg_wdata[1];

  assign intr_state_hmac_err_wd = reg_wdata[2];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_hmac_done_wd = reg_wdata[0];

  assign intr_enable_fifo_empty_wd = reg_wdata[1];

  assign intr_enable_hmac_err_wd = reg_wdata[2];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_hmac_done_wd = reg_wdata[0];

  assign intr_test_fifo_empty_wd = reg_wdata[1];

  assign intr_test_hmac_err_wd = reg_wdata[2];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_wd = reg_wdata[0];
  assign cfg_re = addr_hit[4] & reg_re & !reg_error;
  assign cfg_we = addr_hit[4] & reg_we & !reg_error;

  assign cfg_hmac_en_wd = reg_wdata[0];

  assign cfg_sha_en_wd = reg_wdata[1];

  assign cfg_endian_swap_wd = reg_wdata[2];

  assign cfg_digest_swap_wd = reg_wdata[3];
  assign cmd_we = addr_hit[5] & reg_we & !reg_error;

  assign cmd_hash_start_wd = reg_wdata[0];

  assign cmd_hash_process_wd = reg_wdata[1];
  assign status_re = addr_hit[6] & reg_re & !reg_error;
  assign wipe_secret_we = addr_hit[8] & reg_we & !reg_error;

  assign wipe_secret_wd = reg_wdata[31:0];
  assign key_0_we = addr_hit[9] & reg_we & !reg_error;

  assign key_0_wd = reg_wdata[31:0];
  assign key_1_we = addr_hit[10] & reg_we & !reg_error;

  assign key_1_wd = reg_wdata[31:0];
  assign key_2_we = addr_hit[11] & reg_we & !reg_error;

  assign key_2_wd = reg_wdata[31:0];
  assign key_3_we = addr_hit[12] & reg_we & !reg_error;

  assign key_3_wd = reg_wdata[31:0];
  assign key_4_we = addr_hit[13] & reg_we & !reg_error;

  assign key_4_wd = reg_wdata[31:0];
  assign key_5_we = addr_hit[14] & reg_we & !reg_error;

  assign key_5_wd = reg_wdata[31:0];
  assign key_6_we = addr_hit[15] & reg_we & !reg_error;

  assign key_6_wd = reg_wdata[31:0];
  assign key_7_we = addr_hit[16] & reg_we & !reg_error;

  assign key_7_wd = reg_wdata[31:0];
  assign digest_0_re = addr_hit[17] & reg_re & !reg_error;
  assign digest_1_re = addr_hit[18] & reg_re & !reg_error;
  assign digest_2_re = addr_hit[19] & reg_re & !reg_error;
  assign digest_3_re = addr_hit[20] & reg_re & !reg_error;
  assign digest_4_re = addr_hit[21] & reg_re & !reg_error;
  assign digest_5_re = addr_hit[22] & reg_re & !reg_error;
  assign digest_6_re = addr_hit[23] & reg_re & !reg_error;
  assign digest_7_re = addr_hit[24] & reg_re & !reg_error;

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = cfg_we;
    reg_we_check[5] = cmd_we;
    reg_we_check[6] = 1'b0;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = wipe_secret_we;
    reg_we_check[9] = key_0_we;
    reg_we_check[10] = key_1_we;
    reg_we_check[11] = key_2_we;
    reg_we_check[12] = key_3_we;
    reg_we_check[13] = key_4_we;
    reg_we_check[14] = key_5_we;
    reg_we_check[15] = key_6_we;
    reg_we_check[16] = key_7_we;
    reg_we_check[17] = 1'b0;
    reg_we_check[18] = 1'b0;
    reg_we_check[19] = 1'b0;
    reg_we_check[20] = 1'b0;
    reg_we_check[21] = 1'b0;
    reg_we_check[22] = 1'b0;
    reg_we_check[23] = 1'b0;
    reg_we_check[24] = 1'b0;
    reg_we_check[25] = 1'b0;
    reg_we_check[26] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_hmac_done_qs;
        reg_rdata_next[1] = intr_state_fifo_empty_qs;
        reg_rdata_next[2] = intr_state_hmac_err_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_hmac_done_qs;
        reg_rdata_next[1] = intr_enable_fifo_empty_qs;
        reg_rdata_next[2] = intr_enable_hmac_err_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
        reg_rdata_next[2] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[0] = cfg_hmac_en_qs;
        reg_rdata_next[1] = cfg_sha_en_qs;
        reg_rdata_next[2] = cfg_endian_swap_qs;
        reg_rdata_next[3] = cfg_digest_swap_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[6]: begin
        reg_rdata_next[0] = status_fifo_empty_qs;
        reg_rdata_next[1] = status_fifo_full_qs;
        reg_rdata_next[8:4] = status_fifo_depth_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = err_code_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = digest_0_qs;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = digest_1_qs;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = digest_2_qs;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = digest_3_qs;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = digest_4_qs;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = digest_5_qs;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = digest_6_qs;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = digest_7_qs;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = msg_length_lower_qs;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = msg_length_upper_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// HMAC Core implementation

module hmac_core import hmac_pkg::*; (
  input clk_i,
  input rst_ni,

  input [255:0] secret_key, // {word0, word1, ..., word7}

  input        wipe_secret,
  input [31:0] wipe_v,

  input        hmac_en,

  input        reg_hash_start,
  input        reg_hash_process,
  output logic hash_done,
  output logic sha_hash_start,
  output logic sha_hash_process,
  input        sha_hash_done,

  // fifo
  output logic      sha_rvalid,
  output sha_fifo_t sha_rdata,
  input             sha_rready,

  input             fifo_rvalid,
  input  sha_fifo_t fifo_rdata,
  output logic      fifo_rready,

  // fifo control (select and fifo write data)
  output logic       fifo_wsel,    // 0: from reg, 1: from digest
  output logic       fifo_wvalid,
  output logic [2:0] fifo_wdata_sel, // 0: digest[0] .. 7: digest[7]
  input              fifo_wready,

  input  [63:0] message_length,
  output [63:0] sha_message_length,

  output logic idle
);

  localparam int unsigned BlockSize = 512;
  localparam int unsigned BlockSizeBits = $clog2(BlockSize);
  localparam int unsigned HashWordBits = $clog2($bits(sha_word_t));

  localparam bit [63:0]            BlockSize64 = 64'(BlockSize);
  localparam bit [BlockSizeBits:0] BlockSizeBSB = BlockSize[BlockSizeBits:0];

  logic hash_start; // generated from internal state machine
  logic hash_process; // generated from internal state machine to trigger hash
  logic hmac_hash_done;

  logic [BlockSize-1:0] i_pad ;
  logic [BlockSize-1:0] o_pad ;

  logic [63:0] txcount;
  logic [BlockSizeBits-HashWordBits-1:0] pad_index;
  logic clr_txcount, inc_txcount;

  logic hmac_sha_rvalid;

  typedef enum logic [1:0] {
    SelIPad,
    SelOPad,
    SelFifo
  } sel_rdata_t;

  sel_rdata_t sel_rdata;

  typedef enum logic {
    SelIPadMsg,
    SelOPadMsg
  } sel_msglen_t;

  sel_msglen_t sel_msglen;

  typedef enum logic {
    Inner,  // Update when state goes to StIPad
    Outer   // Update when state enters StOPad
  } round_t ;

  logic update_round ;
  round_t round_q, round_d;

  typedef enum logic [2:0] {
    StIdle,
    StIPad,
    StMsg,              // Actual Msg, and Digest both
    StPushToMsgFifo,    // Digest --> Msg Fifo
    StWaitResp,         // Hash done( by checking processed_length? or hash_done)
    StOPad,
    StDone              // hmac_done
  } st_e ;

  st_e st_q, st_d;

  logic clr_fifo_wdata_sel;
  logic txcnt_eq_blksz ;

  logic reg_hash_process_flag;

  assign sha_hash_start   = (hmac_en) ? hash_start                       : reg_hash_start ;
  assign sha_hash_process = (hmac_en) ? reg_hash_process | hash_process  : reg_hash_process ;
  assign hash_done        = (hmac_en) ? hmac_hash_done                   : sha_hash_done  ;

  assign pad_index = txcount[BlockSizeBits-1:HashWordBits];

  assign i_pad = {secret_key, {(BlockSize-256){1'b0}}} ^ {(BlockSize/8){8'h36}};
  assign o_pad = {secret_key, {(BlockSize-256){1'b0}}} ^ {(BlockSize/8){8'h5c}};


  assign fifo_rready  = (hmac_en) ? (st_q == StMsg) & sha_rready : sha_rready ;
  // sha_rvalid is controlled by State Machine below.
  assign sha_rvalid = (!hmac_en) ? fifo_rvalid : hmac_sha_rvalid ;
  assign sha_rdata =
    (!hmac_en)             ? fifo_rdata                                               :
    (sel_rdata == SelIPad) ? '{data: i_pad[(BlockSize-1)-32*pad_index-:32], mask: '1} :
    (sel_rdata == SelOPad) ? '{data: o_pad[(BlockSize-1)-32*pad_index-:32], mask: '1} :
    (sel_rdata == SelFifo) ? fifo_rdata                                               :
    '{default: '0};

  assign sha_message_length = (!hmac_en)                 ? message_length               :
                              (sel_msglen == SelIPadMsg) ? message_length + BlockSize64 :
                              (sel_msglen == SelOPadMsg) ? BlockSize64 + 64'd256        :
                              '0 ;

  assign txcnt_eq_blksz = (txcount[BlockSizeBits:0] == BlockSizeBSB);

  assign inc_txcount = sha_rready && sha_rvalid;

  // txcount
  //    Looks like txcount can be removed entirely here in hmac_core
  //    In the first round (InnerPaddedKey), it can just watch process and hash_done
  //    In the second round, it only needs count 256 bits for hash digest to trigger
  //    hash_process to SHA2
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      txcount <= '0;
    end else if (clr_txcount) begin
      txcount <= '0;
    end else if (inc_txcount) begin
      txcount[63:5] <= txcount[63:5] + 1'b1;
    end
  end

  // reg_hash_process trigger logic
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      reg_hash_process_flag <= 1'b0;
    end else if (reg_hash_process) begin
      reg_hash_process_flag <= 1'b1;
    end else if (hmac_hash_done || reg_hash_start) begin
      reg_hash_process_flag <= 1'b0;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      round_q <= Inner;
    end else if (update_round) begin
      round_q <= round_d;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      fifo_wdata_sel <= 3'h 0;
    end else if (clr_fifo_wdata_sel) begin
      fifo_wdata_sel <= 3'h 0;
    end else if (fifo_wsel && fifo_wvalid) begin
      fifo_wdata_sel <= fifo_wdata_sel + 1'b1;
    end
  end

  assign sel_msglen = (round_q == Inner) ? SelIPadMsg : SelOPadMsg ;

  always_ff @(posedge clk_i or negedge rst_ni) begin : state_ff
    if (!rst_ni) st_q <= StIdle;
    else         st_q <= st_d;
  end

  always_comb begin : next_state
    hmac_hash_done  = 1'b0;
    hmac_sha_rvalid = 1'b0;

    clr_txcount = 1'b0;

    update_round = 1'b0;
    round_d      = Inner;

    fifo_wsel    = 1'b0;   // from register
    fifo_wvalid  = 1'b0;

    clr_fifo_wdata_sel = 1'b1;

    sel_rdata = SelFifo;

    hash_start   = 1'b0;
    hash_process = 1'b0;

    unique case (st_q)
      StIdle: begin
        if (hmac_en && reg_hash_start) begin
          st_d = StIPad;

          clr_txcount  = 1'b1;
          update_round = 1'b1;
          round_d      = Inner;
          hash_start   = 1'b1;
        end else begin
          st_d = StIdle;
        end
      end

      StIPad: begin
        sel_rdata = SelIPad;

        if (txcnt_eq_blksz) begin
          st_d = StMsg;

          hmac_sha_rvalid = 1'b0; // block new read request
        end else begin
          st_d = StIPad;

          hmac_sha_rvalid = 1'b1;
        end
      end

      StMsg: begin
        sel_rdata = SelFifo;
        fifo_wsel = (round_q == Outer);

        if ( (((round_q == Inner) && reg_hash_process_flag) || (round_q == Outer))
            && (txcount >= sha_message_length)) begin
          st_d = StWaitResp;

          hmac_sha_rvalid = 1'b0; // block
          hash_process = (round_q == Outer);
        end else begin
          st_d = StMsg;

          hmac_sha_rvalid = fifo_rvalid;
        end
      end

      StWaitResp: begin
        hmac_sha_rvalid = 1'b0;

        if (sha_hash_done) begin
          if (round_q == Outer) begin
            st_d = StDone;
          end else begin // round_q == Inner
            st_d = StPushToMsgFifo;
          end
        end else begin
          st_d = StWaitResp;
        end
      end

      StPushToMsgFifo: begin
        hmac_sha_rvalid    = 1'b0;
        fifo_wsel          = 1'b1;
        fifo_wvalid        = 1'b1;
        clr_fifo_wdata_sel = 1'b0;

        if (fifo_wready && fifo_wdata_sel == 3'h7) begin
          st_d = StOPad;

          clr_txcount  = 1'b1;
          update_round = 1'b1;
          round_d      = Outer;
          hash_start   = 1'b1;
        end else begin
          st_d = StPushToMsgFifo;

        end
      end

      StOPad: begin
        sel_rdata = SelOPad;
        fifo_wsel = 1'b1; // Remained HMAC select to indicate HMAC is in second stage

        if (txcnt_eq_blksz) begin
          st_d = StMsg;

          hmac_sha_rvalid = 1'b0; // block new read request
        end else begin
          st_d = StOPad;

          hmac_sha_rvalid = 1'b1;
        end
      end

      StDone: begin
        // raise interrupt (hash_done)
        st_d = StIdle;

        hmac_hash_done = 1'b1;
      end

      default: begin
        st_d = StIdle;
      end

    endcase
  end

  // Idle: Idle in HMAC_CORE only represents the idle status when hmac mode is
  // set. If hmac_en is 0, this logic sends the idle signal always.
  assign idle = (st_q == StIdle) && !reg_hash_start;
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// HMAC-SHA256

`include "prim_assert.sv"

module hmac
  import hmac_pkg::*;
  import hmac_reg_pkg::*;
#(
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}}
) (
  input clk_i,
  input rst_ni,

  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  output logic intr_hmac_done_o,
  output logic intr_fifo_empty_o,
  output logic intr_hmac_err_o,

  output prim_mubi_pkg::mubi4_t idle_o
);


  /////////////////////////
  // Signal declarations //
  /////////////////////////
  hmac_reg2hw_t reg2hw;
  hmac_hw2reg_t hw2reg;

  tlul_pkg::tl_h2d_t  tl_win_h2d;
  tlul_pkg::tl_d2h_t  tl_win_d2h;

  logic [255:0] secret_key;

  logic        wipe_secret;
  logic [31:0] wipe_v;

  logic        fifo_rvalid;
  logic        fifo_rready;
  sha_fifo_t   fifo_rdata;

  logic        fifo_wvalid, fifo_wready;
  sha_fifo_t   fifo_wdata;
  logic        fifo_full;
  logic        fifo_empty;
  logic [4:0]  fifo_depth;

  logic        msg_fifo_req;
  logic        msg_fifo_gnt;
  logic        msg_fifo_we;
  logic [31:0] msg_fifo_wdata;
  logic [31:0] msg_fifo_wmask;
  logic [31:0] msg_fifo_rdata;
  logic        msg_fifo_rvalid;
  logic [1:0]  msg_fifo_rerror;
  logic [31:0] msg_fifo_wdata_endian;
  logic [31:0] msg_fifo_wmask_endian;

  logic        packer_ready;
  logic        packer_flush_done;

  logic        reg_fifo_wvalid;
  sha_word_t   reg_fifo_wdata;
  sha_word_t   reg_fifo_wmask;
  logic        hmac_fifo_wsel;
  logic        hmac_fifo_wvalid;
  logic [2:0]  hmac_fifo_wdata_sel;

  logic        shaf_rvalid;
  sha_fifo_t   shaf_rdata;
  logic        shaf_rready;

  logic        sha_en;
  logic        hmac_en;
  logic        endian_swap;
  logic        digest_swap;

  logic        reg_hash_start;
  logic        sha_hash_start;
  logic        hash_start;      // Valid hash_start_signal
  logic        reg_hash_process;
  logic        sha_hash_process;

  logic        reg_hash_done;
  logic        sha_hash_done;

  logic [63:0] message_length;
  logic [63:0] sha_message_length;

  err_code_e   err_code;
  logic        err_valid;

  sha_word_t [7:0] digest;

  hmac_reg2hw_cfg_reg_t cfg_reg;
  logic                 cfg_block;  // Prevent changing config
  logic                 msg_allowed; // MSG_FIFO from software is allowed

  logic hmac_core_idle;
  logic sha_core_idle;

  ///////////////////////
  // Connect registers //
  ///////////////////////
  assign hw2reg.status.fifo_full.d  = fifo_full;
  assign hw2reg.status.fifo_empty.d = fifo_empty;
  assign hw2reg.status.fifo_depth.d = fifo_depth;

  // secret key
  assign wipe_secret = reg2hw.wipe_secret.qe;
  assign wipe_v      = reg2hw.wipe_secret.q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      secret_key <= '0;
    end else if (wipe_secret) begin
      secret_key <= {8{wipe_v}};
    end else if (!cfg_block) begin
      // Allow updating secret key only when the engine is in Idle.
      for (int i = 0; i < 8; i++) begin
        if (reg2hw.key[7-i].qe) begin
          secret_key[32*i+:32] <= reg2hw.key[7-i].q;
        end
      end
    end
  end

  for (genvar i = 0; i < 8; i++) begin : gen_key_digest
    assign hw2reg.key[7-i].d      = '0;
    // digest
    assign hw2reg.digest[i].d = conv_endian(digest[i], digest_swap);
  end

  logic [3:0] unused_cfg_qe;

  assign unused_cfg_qe = {cfg_reg.sha_en.qe,      cfg_reg.hmac_en.qe,
                          cfg_reg.endian_swap.qe, cfg_reg.digest_swap.qe};

  assign sha_en      = cfg_reg.sha_en.q;
  assign hmac_en     = cfg_reg.hmac_en.q;
  assign endian_swap = cfg_reg.endian_swap.q;
  assign digest_swap = cfg_reg.digest_swap.q;
  assign hw2reg.cfg.hmac_en.d     = cfg_reg.hmac_en.q;
  assign hw2reg.cfg.sha_en.d      = cfg_reg.sha_en.q;
  assign hw2reg.cfg.endian_swap.d = cfg_reg.endian_swap.q;
  assign hw2reg.cfg.digest_swap.d = cfg_reg.digest_swap.q;

  assign reg_hash_start   = reg2hw.cmd.hash_start.qe   & reg2hw.cmd.hash_start.q;
  assign reg_hash_process = reg2hw.cmd.hash_process.qe & reg2hw.cmd.hash_process.q;

  // Error code register
  assign hw2reg.err_code.de = err_valid;
  assign hw2reg.err_code.d  = err_code;

  /////////////////////
  // Control signals //
  /////////////////////
  assign hash_start = reg_hash_start & sha_en & ~cfg_block;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      cfg_block <= '0;
    end else if (hash_start) begin
      cfg_block <= 1'b 1;
    end else if (reg_hash_done) begin
      cfg_block <= 1'b 0;
    end
  end
  // Hold the configuration during the process
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      cfg_reg <= '{
        endian_swap: '{
          q: HMAC_CFG_ENDIAN_SWAP_RESVAL,
          qe: 1'b0
        },
        default:'0
      };
    end else if (!cfg_block && reg2hw.cfg.hmac_en.qe) begin
      cfg_reg <= reg2hw.cfg ;
    end
  end

  // Open up the MSG_FIFO from the TL-UL port when it is ready
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      msg_allowed <= '0;
    end else if (hash_start) begin
      msg_allowed <= 1'b 1;
    end else if (packer_flush_done) begin
      msg_allowed <= 1'b 0;
    end
  end
  ////////////////
  // Interrupts //
  ////////////////
  logic fifo_empty_q, fifo_empty_event;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      fifo_empty_q <= '1; // By default, it is empty
    end else if (!hmac_fifo_wsel) begin
      fifo_empty_q <= fifo_empty;
    end
  end
  assign fifo_empty_event = fifo_empty & ~fifo_empty_q;

  logic [2:0] event_intr;
  assign event_intr = {err_valid, fifo_empty_event, reg_hash_done};

  // instantiate interrupt hardware primitive
  prim_intr_hw #(.Width(1)) intr_hw_hmac_done (
    .clk_i,
    .rst_ni,
    .event_intr_i           (event_intr[0]),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.hmac_done.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.hmac_done.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.hmac_done.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.hmac_done.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.hmac_done.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.hmac_done.d),
    .intr_o                 (intr_hmac_done_o)
  );
  prim_intr_hw #(.Width(1)) intr_hw_fifo_empty (
    .clk_i,
    .rst_ni,
    .event_intr_i           (event_intr[1]),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.fifo_empty.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.fifo_empty.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.fifo_empty.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.fifo_empty.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.fifo_empty.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.fifo_empty.d),
    .intr_o                 (intr_fifo_empty_o)
  );
  prim_intr_hw #(.Width(1)) intr_hw_hmac_err (
    .clk_i,
    .rst_ni,
    .event_intr_i           (event_intr[2]),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.hmac_err.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.hmac_err.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.hmac_err.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.hmac_err.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.hmac_err.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.hmac_err.d),
    .intr_o                 (intr_hmac_err_o)
  );

  ///////////////
  // Instances //
  ///////////////

  assign msg_fifo_rvalid = msg_fifo_req & ~msg_fifo_we;
  assign msg_fifo_rdata  = '1;  // Return all F
  assign msg_fifo_rerror = '1;  // Return error for read access
  assign msg_fifo_gnt    = msg_fifo_req & ~hmac_fifo_wsel & packer_ready;

  // FIFO control
  sha_fifo_t reg_fifo_wentry;
  assign reg_fifo_wentry.data = conv_endian(reg_fifo_wdata, 1'b1); // always convert
  assign reg_fifo_wentry.mask = {reg_fifo_wmask[0],  reg_fifo_wmask[8],
                                 reg_fifo_wmask[16], reg_fifo_wmask[24]};
  assign fifo_full   = ~fifo_wready;
  assign fifo_empty  = ~fifo_rvalid;
  assign fifo_wvalid = (hmac_fifo_wsel && fifo_wready) ? hmac_fifo_wvalid : reg_fifo_wvalid;
  assign fifo_wdata  = (hmac_fifo_wsel) ? '{data: digest[hmac_fifo_wdata_sel], mask: '1}
                                       : reg_fifo_wentry;

  prim_fifo_sync #(
    .Width   ($bits(sha_fifo_t)),
    .Pass    (1'b1),
    .Depth   (MsgFifoDepth)
  ) u_msg_fifo (
    .clk_i,
    .rst_ni,
    .clr_i   (1'b0),

    .wvalid_i(fifo_wvalid & sha_en),
    .wready_o(fifo_wready),
    .wdata_i (fifo_wdata),

    .depth_o (fifo_depth),
    .full_o  (),

    .rvalid_o(fifo_rvalid),
    .rready_i(fifo_rready),
    .rdata_o (fifo_rdata),
    .err_o   ()
  );

  // TL ADAPTER SRAM
  tlul_adapter_sram #(
    .SramAw (9),
    .SramDw (32),
    .Outstanding (1),
    .ByteAccess  (1),
    .ErrOnRead   (1)
  ) u_tlul_adapter (
    .clk_i,
    .rst_ni,
    .tl_i        (tl_win_h2d),
    .tl_o        (tl_win_d2h),
    .en_ifetch_i (prim_mubi_pkg::MuBi4False),
    .req_o       (msg_fifo_req   ),
    .req_type_o  (               ),
    .gnt_i       (msg_fifo_gnt   ),
    .we_o        (msg_fifo_we    ),
    .addr_o      (               ), // Doesn't care the address other than sub-word
    .wdata_o     (msg_fifo_wdata ),
    .wmask_o     (msg_fifo_wmask ),
    .intg_error_o(               ),
    .rdata_i     (msg_fifo_rdata ),
    .rvalid_i    (msg_fifo_rvalid),
    .rerror_i    (msg_fifo_rerror)
  );

  // TL-UL to MSG_FIFO byte write handling
  logic msg_write;

  assign msg_write = msg_fifo_req & msg_fifo_we & ~hmac_fifo_wsel & msg_allowed;

  logic [$clog2(32+1)-1:0] wmask_ones;

  always_comb begin
    wmask_ones = '0;
    for (int i = 0 ; i < 32 ; i++) begin
      wmask_ones = wmask_ones + msg_fifo_wmask[i];
    end
  end

  // Calculate written message
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      message_length <= '0;
    end else if (hash_start) begin
      message_length <= '0;
    end else if (msg_write && sha_en && packer_ready) begin
      message_length <= message_length + 64'(wmask_ones);
    end
  end

  assign hw2reg.msg_length_upper.de = 1'b1;
  assign hw2reg.msg_length_upper.d = message_length[63:32];
  assign hw2reg.msg_length_lower.de = 1'b1;
  assign hw2reg.msg_length_lower.d = message_length[31:0];


  // Convert endian here
  //    prim_packer always packs to the right, but SHA engine assumes incoming
  //    to be big-endian, [31:24] comes first. So, the data is reverted after
  //    prim_packer before the message fifo. here to reverse if not big-endian
  //    before pushing to the packer.
  assign msg_fifo_wdata_endian = conv_endian(msg_fifo_wdata, endian_swap);
  assign msg_fifo_wmask_endian = conv_endian(msg_fifo_wmask, endian_swap);

  prim_packer #(
    .InW          (32),
    .OutW         (32),
    .EnProtection (1'b 0)
  ) u_packer (
    .clk_i,
    .rst_ni,

    .valid_i      (msg_write & sha_en),
    .data_i       (msg_fifo_wdata_endian),
    .mask_i       (msg_fifo_wmask_endian),
    .ready_o      (packer_ready),

    .valid_o      (reg_fifo_wvalid),
    .data_o       (reg_fifo_wdata),
    .mask_o       (reg_fifo_wmask),
    .ready_i      (fifo_wready & ~hmac_fifo_wsel),

    .flush_i      (reg_hash_process),
    .flush_done_o (packer_flush_done), // ignore at this moment

    .err_o  () // Not used
  );


  hmac_core u_hmac (
    .clk_i,
    .rst_ni,

    .secret_key,

    .wipe_secret,
    .wipe_v,

    .hmac_en,

    .reg_hash_start   (hash_start),
    .reg_hash_process (packer_flush_done), // Trigger after all msg written
    .hash_done      (reg_hash_done),
    .sha_hash_start,
    .sha_hash_process,
    .sha_hash_done,

    .sha_rvalid     (shaf_rvalid),
    .sha_rdata      (shaf_rdata),
    .sha_rready     (shaf_rready),

    .fifo_rvalid,
    .fifo_rdata,
    .fifo_rready,

    .fifo_wsel      (hmac_fifo_wsel),
    .fifo_wvalid    (hmac_fifo_wvalid),
    .fifo_wdata_sel (hmac_fifo_wdata_sel),
    .fifo_wready,

    .message_length,
    .sha_message_length,

    .idle           (hmac_core_idle)
  );

  sha2 u_sha2 (
    .clk_i,
    .rst_ni,

    .wipe_secret,
    .wipe_v,

    .fifo_rvalid      (shaf_rvalid),
    .fifo_rdata       (shaf_rdata),
    .fifo_rready      (shaf_rready),

    .sha_en,
    .hash_start       (sha_hash_start),
    .hash_process     (sha_hash_process),
    .hash_done        (sha_hash_done),

    .message_length   (sha_message_length),

    .digest,

    .idle             (sha_core_idle)
  );

  // Register top
  logic [NumAlerts-1:0] alert_test, alerts;
  hmac_reg_top u_reg (
    .clk_i,
    .rst_ni,

    .tl_i,
    .tl_o,

    .tl_win_o   (tl_win_h2d),
    .tl_win_i   (tl_win_d2h),

    .reg2hw,
    .hw2reg,

    // SEC_CM: BUS.INTEGRITY
    .intg_err_o (alerts[0]),
    .devmode_i  (1'b1)
  );

  // Alerts
  assign alert_test = {
    reg2hw.alert_test.q &
    reg2hw.alert_test.qe
  };

  localparam logic [NumAlerts-1:0] AlertIsFatal = {1'b1};
  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(AlertIsFatal[i])
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i] ),
      .alert_req_i   ( alerts[0]     ),
      .alert_ack_o   (               ),
      .alert_state_o (               ),
      .alert_rx_i    ( alert_rx_i[i] ),
      .alert_tx_o    ( alert_tx_o[i] )
    );
  end

  /////////////////////////
  // HMAC Error Handling //
  /////////////////////////
  logic hash_start_sha_disabled, update_seckey_inprocess;
  logic hash_start_active;  // `reg_hash_start` set when hash already in active
  logic msg_push_not_allowed; // Message is received when `hash_start` isn't set
  assign hash_start_sha_disabled = reg_hash_start & ~sha_en;
  assign hash_start_active = reg_hash_start & cfg_block;
  assign msg_push_not_allowed = msg_fifo_req & ~msg_allowed;

  always_comb begin
    update_seckey_inprocess = 1'b0;
    if (cfg_block) begin
      for (int i = 0 ; i < 8 ; i++) begin
        if (reg2hw.key[i].qe) begin
          update_seckey_inprocess = update_seckey_inprocess | 1'b1;
        end
      end
    end else begin
      update_seckey_inprocess = 1'b0;
    end
  end

  // Update ERR_CODE register and interrupt only when no pending interrupt.
  // This ensures only the first event of the series of events can be seen to sw.
  // It is recommended that the software reads ERR_CODE register when interrupt
  // is pending to avoid any race conditions.
  assign err_valid = ~reg2hw.intr_state.hmac_err.q &
                   ( hash_start_sha_disabled | update_seckey_inprocess
                   | hash_start_active | msg_push_not_allowed );

  always_comb begin
    err_code = NoError;
    unique case (1'b1)
      hash_start_sha_disabled: begin
        err_code = SwHashStartWhenShaDisabled;
      end

      update_seckey_inprocess: begin
        err_code = SwUpdateSecretKeyInProcess;
      end

      hash_start_active: begin
        err_code = SwHashStartWhenActive;
      end

      msg_push_not_allowed: begin
        err_code = SwPushMsgWhenDisallowed;
      end

      default: begin
        err_code = NoError;
      end
    endcase
  end

  /////////////////////
  // Unused Signals  //
  /////////////////////
  logic unused_wmask;
  assign unused_wmask = ^reg_fifo_wmask;

  /////////////////////
  // Idle output     //
  /////////////////////
  // TBD this should be connected later
  // Idle: AND condition of:
  //  - packer empty: Currently no way to guarantee the packer is empty.
  //    temporary, the logic uses packer output (reg_fifo_wvalid)
  //  - MSG_FIFO  --> fifo_rvalid
  //  - HMAC_CORE --> hmac_core_idle
  //  - SHA2_CORE --> sha_core_idle
  //  - Clean interrupt status
  // ICEBOX(#12958): Revise prim_packer and replace `reg_fifo_wvalid` to the
  // empty status.
  logic idle;
  assign idle = !reg_fifo_wvalid && !fifo_rvalid
              && hmac_core_idle && sha_core_idle;

  prim_mubi_pkg::mubi4_t idle_q, idle_d;
  assign idle_d = prim_mubi_pkg::mubi4_bool_to_mubi(idle);
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      idle_q <= prim_mubi_pkg::MuBi4False;
    end else begin
      idle_q <= idle_d;
    end
  end
  assign idle_o = idle_q;

  //////////////////////////////////////////////
  // Assertions, Assumptions, and Coverpoints //
  //////////////////////////////////////////////

`ifndef VERILATOR
`ifndef SYNTHESIS
  // HMAC assumes TL-UL mask is byte-aligned.
  property wmask_bytealign_p(wmask_byte, clk, rst_n);
    @(posedge clk) disable iff (rst_n == 0)
      msg_fifo_req & msg_fifo_we |-> wmask_byte inside {'0, '1};
  endproperty

  for (genvar i = 0 ; i < 4; i++) begin: gen_assert_wmask_bytealign
    assert property (wmask_bytealign_p(msg_fifo_wmask[8*i+:8], clk_i, rst_ni));
  end

  // To pass FPV, this shouldn't add pragma translate_off even these two signals
  // are used in Assertion only
  logic in_process;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)               in_process <= 1'b0;
    else if (reg_hash_process) in_process <= 1'b1;
    else if (reg_hash_done)    in_process <= 1'b0;
  end

  logic initiated;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)               initiated <= 1'b0;
    else if (hash_start)       initiated <= 1'b1;
    else if (reg_hash_process) initiated <= 1'b0;
  end

  // the host doesn't write data after hash_process until hash_start.
  // Same as "message_length shouldn't be changed between hash_process and done
  `ASSERT(ValidWriteAssert, msg_fifo_req |-> !in_process)

  // `hash_process` shall be toggle and paired with `hash_start`.
  // Below condition is covered by the design (2020-02-19)
  //`ASSERT(ValidHashStartAssert, hash_start |-> !initiated)
  `ASSERT(ValidHashProcessAssert, reg_hash_process |-> initiated)

  // between `hash_done` and `hash_start`, message FIFO should be empty
  `ASSERT(MsgFifoEmptyWhenNoOpAssert,
          !in_process && !initiated |-> $stable(message_length))

  // hmac_en should be modified only when the logic is Idle
  `ASSERT(ValidHmacEnConditionAssert,
          hmac_en != $past(hmac_en) |-> !in_process && !initiated)

  // All outputs should be known value after reset
  `ASSERT_KNOWN(IntrHmacDoneOKnown, intr_hmac_done_o)
  `ASSERT_KNOWN(IntrFifoEmptyOKnown, intr_fifo_empty_o)
  `ASSERT_KNOWN(TlODValidKnown, tl_o.d_valid)
  `ASSERT_KNOWN(TlOAReadyKnown, tl_o.a_ready)
  `ASSERT_KNOWN(AlertKnownO_A, alert_tx_o)

`endif // SYNTHESIS
`endif // VERILATOR

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[0])
endmodule


module sram_array_1p1024x39m39(
  input logic         clk_i,
  input logic [9:0]   addr_i,
  input logic         req_i,
  input logic         write_i,
  input logic         wmask_i,
  input logic [38:0] wdata_i,
  output logic [38:0] rdata_o
);

localparam Width = 39;
localparam DataBitsPerMask = 39;
localparam MaskWidth = 1;

logic [Width-1:0]     mem [1024];
// logic [MaskWidth-1:0] wmask;

 always @(posedge clk_i) begin
    if (req_i) begin
      if (write_i) begin
        for (int i=0; i < MaskWidth; i = i + 1) begin
          if (wmask_i) begin
            mem[addr_i][i*DataBitsPerMask +: DataBitsPerMask] <=
              wdata_i[i*DataBitsPerMask +: DataBitsPerMask];
          end
        end
      end else begin
        rdata_o <= mem[addr_i];
      end
    end
 end

endmodule

module sram_array_1p128x312m39(
  input logic         clk_i,
  input logic [6:0]   addr_i,
  input logic         req_i,
  input logic         write_i,
  input logic [7:0]   wmask_i,
  input logic [311:0] wdata_i,
  output logic [311:0] rdata_o
);

localparam Width = 312;
localparam DataBitsPerMask = 39;
localparam MaskWidth = 8;

logic [Width-1:0]     mem [128];
// logic [MaskWidth-1:0] wmask;

 always @(posedge clk_i) begin
    if (req_i) begin
      if (write_i) begin
        for (int i=0; i < MaskWidth; i = i + 1) begin
          if (wmask_i[i]) begin
            mem[addr_i][i*DataBitsPerMask +: DataBitsPerMask] <=
              wdata_i[i*DataBitsPerMask +: DataBitsPerMask];
          end
        end
      end else begin
        rdata_o <= mem[addr_i];
      end
    end
 end

endmodule

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN Controller
 */
module otbn_controller
  import otbn_pkg::*;
#(
  // Size of the instruction memory, in bytes
  parameter int ImemSizeByte = 4096,
  // Size of the data memory, in bytes
  parameter int DmemSizeByte = 4096,

  localparam int ImemAddrWidth = prim_util_pkg::vbits(ImemSizeByte),
  localparam int DmemAddrWidth = prim_util_pkg::vbits(DmemSizeByte)
) (
  input logic clk_i,
  input logic rst_ni,

  input  logic start_i,   // start the processing at address zero
  output logic locking_o, // Controller is in or is entering the locked state
  input  logic err_bit_clear_i,

  input prim_mubi_pkg::mubi4_t fatal_escalate_en_i,
  input prim_mubi_pkg::mubi4_t recov_escalate_en_i,
  input prim_mubi_pkg::mubi4_t rma_req_i,
  output controller_err_bits_t err_bits_o,
  output logic                 recoverable_err_o,

  // Next instruction selection (to instruction fetch)
  output logic                     insn_fetch_req_valid_o,
  output logic                     insn_fetch_req_valid_raw_o,
  output logic [ImemAddrWidth-1:0] insn_fetch_req_addr_o,
  output logic                     insn_fetch_resp_clear_o,

  // Fetched/decoded instruction
  input logic                     insn_valid_i,
  input logic                     insn_illegal_i,
  input logic [ImemAddrWidth-1:0] insn_addr_i,

  // Decoded instruction data
  input insn_dec_base_t   insn_dec_base_i,
  input insn_dec_bignum_t insn_dec_bignum_i,
  input insn_dec_shared_t insn_dec_shared_i,

  // Base register file
  output logic [4:0]               rf_base_wr_addr_o,
  output logic                     rf_base_wr_en_o,
  output logic                     rf_base_wr_commit_o,
  output logic [31:0]              rf_base_wr_data_no_intg_o,
  output logic [BaseIntgWidth-1:0] rf_base_wr_data_intg_o,
  output logic                     rf_base_wr_data_intg_sel_o,

  output logic [4:0]               rf_base_rd_addr_a_o,
  output logic                     rf_base_rd_en_a_o,
  input  logic [BaseIntgWidth-1:0] rf_base_rd_data_a_intg_i,
  output logic [4:0]               rf_base_rd_addr_b_o,
  output logic                     rf_base_rd_en_b_o,
  input  logic [BaseIntgWidth-1:0] rf_base_rd_data_b_intg_i,
  output logic                     rf_base_rd_commit_o,

  input logic rf_base_call_stack_sw_err_i,
  input logic rf_base_call_stack_hw_err_i,

  // Bignum register file (WDRs)
  output logic [4:0]         rf_bignum_wr_addr_o,
  output logic [1:0]         rf_bignum_wr_en_o,
  output logic               rf_bignum_wr_commit_o,
  output logic [WLEN-1:0]    rf_bignum_wr_data_no_intg_o,
  output logic [ExtWLEN-1:0] rf_bignum_wr_data_intg_o,
  output logic               rf_bignum_wr_data_intg_sel_o,

  output logic [4:0]         rf_bignum_rd_addr_a_o,
  output logic               rf_bignum_rd_en_a_o,
  input  logic [ExtWLEN-1:0] rf_bignum_rd_data_a_intg_i,

  output logic [4:0]         rf_bignum_rd_addr_b_o,
  output logic               rf_bignum_rd_en_b_o,
  input  logic [ExtWLEN-1:0] rf_bignum_rd_data_b_intg_i,

  input logic rf_bignum_intg_err_i,
  input logic rf_bignum_spurious_we_err_i,

  output logic [NWdr-1:0] rf_bignum_rd_a_indirect_onehot_o,
  output logic [NWdr-1:0] rf_bignum_rd_b_indirect_onehot_o,
  output logic [NWdr-1:0] rf_bignum_wr_indirect_onehot_o,
  output logic            rf_bignum_indirect_en_o,

  // Execution units

  // Base ALU
  output alu_base_operation_t  alu_base_operation_o,
  output alu_base_comparison_t alu_base_comparison_o,
  input  logic [31:0]          alu_base_operation_result_i,
  input  logic                 alu_base_comparison_result_i,

  // Bignum ALU
  output alu_bignum_operation_t alu_bignum_operation_o,
  output logic                  alu_bignum_operation_valid_o,
  output logic                  alu_bignum_operation_commit_o,
  input  logic [WLEN-1:0]       alu_bignum_operation_result_i,
  input  logic                  alu_bignum_selection_flag_i,

  // Bignum MAC
  output mac_bignum_operation_t mac_bignum_operation_o,
  input  logic [WLEN-1:0]       mac_bignum_operation_result_i,
  output logic                  mac_bignum_en_o,
  output logic                  mac_bignum_commit_o,

  // LSU
  output logic                     lsu_load_req_o,
  output logic                     lsu_store_req_o,
  output insn_subset_e             lsu_req_subset_o,
  output logic [DmemAddrWidth-1:0] lsu_addr_o,
  input  logic                     lsu_addr_en_predec_i,

  output logic [BaseIntgWidth-1:0] lsu_base_wdata_o,
  output logic [ExtWLEN-1:0]       lsu_bignum_wdata_o,

  input  logic [BaseIntgWidth-1:0] lsu_base_rdata_i,
  input  logic [ExtWLEN-1:0]       lsu_bignum_rdata_i,

  // Internal Special-Purpose Registers (ISPRs)
  output ispr_e                       ispr_addr_o,
  output logic [31:0]                 ispr_base_wdata_o,
  output logic [BaseWordsPerWLEN-1:0] ispr_base_wr_en_o,
  output logic [ExtWLEN-1:0]          ispr_bignum_wdata_intg_o,
  output logic                        ispr_bignum_wr_en_o,
  output logic [NFlagGroups-1:0]      ispr_flags_wr_o,
  output logic                        ispr_wr_commit_o,
  input  logic [ExtWLEN-1:0]          ispr_rdata_intg_i,
  output logic                        ispr_rd_en_o,

  // RND interface
  output logic rnd_req_o,
  output logic rnd_prefetch_req_o,
  input  logic rnd_valid_i,

  input  logic urnd_reseed_err_i,

  // Secure Wipe
  output logic secure_wipe_req_o,
  input  logic secure_wipe_ack_i,
  input  logic sec_wipe_zero_i,
  input  logic secure_wipe_running_i,

  input  logic        state_reset_i,
  output logic [31:0] insn_cnt_o,
  input  logic        insn_cnt_clear_i,
  output logic        mems_sec_wipe_o,

  input  logic        software_errs_fatal_i,

  input logic [1:0] sideload_key_shares_valid_i,

  // Prefetch stage control
  output logic                     prefetch_en_o,
  output logic                     prefetch_loop_active_o,
  output logic [31:0]              prefetch_loop_iterations_o,
  output logic [ImemAddrWidth:0]   prefetch_loop_end_addr_o,
  output logic [ImemAddrWidth-1:0] prefetch_loop_jump_addr_o,
  output logic                     prefetch_ignore_errs_o,

  // Predecoded control
  input  ctrl_flow_predec_t        ctrl_flow_predec_i,
  input  logic [ImemAddrWidth-1:0] ctrl_flow_target_predec_i,
  output logic                     predec_error_o
);
  import prim_mubi_pkg::*;

  otbn_state_e state_q, state_d;


  controller_err_bits_t err_bits_q, err_bits_d;

  // The specific error signals that go into err_bits_d
  logic fatal_software_err, bad_internal_state_err, reg_intg_violation_err, key_invalid_err;
  logic illegal_insn_err, bad_data_addr_err, call_stack_sw_err, bad_insn_addr_err;

  logic err;
  logic internal_err;
  logic recoverable_err;
  logic software_err;
  logic non_insn_addr_software_err;
  logic fatal_err;
  logic internal_fatal_err;
  logic done_complete;
  logic executing;
  logic state_error, state_error_d, state_error_q;
  logic spurious_secure_wipe_ack_q, spurious_secure_wipe_ack_d;
  logic mubi_err_q, mubi_err_d;

  logic                     insn_fetch_req_valid_raw;
  logic [ImemAddrWidth-1:0] insn_fetch_req_addr_last;

  logic stall;
  logic ispr_stall;
  logic mem_stall;
  logic rf_indirect_stall;
  logic jump_or_branch;
  logic branch_taken;
  logic insn_executing;
  logic ld_insn_with_addr_from_call_stack, st_insn_with_addr_from_call_stack;
  logic [ImemAddrWidth-1:0] branch_target;
  logic                     branch_target_overflow;
  logic [ImemAddrWidth:0]   next_insn_addr_wide;
  logic [ImemAddrWidth-1:0] next_insn_addr;

  csr_e                                csr_addr;
  logic [$clog2(BaseWordsPerWLEN)-1:0] csr_sub_addr;
  logic [31:0]                         csr_rdata_raw;
  logic [31:0]                         csr_rdata;
  logic [BaseWordsPerWLEN-1:0]         csr_rdata_mux [32];
  logic [31:0]                         csr_wdata_raw;
  logic [31:0]                         csr_wdata;

  wsr_e                                wsr_addr;
  logic [WLEN-1:0]                     wsr_wdata;

  ispr_e                               ispr_addr_base;
  logic [$clog2(BaseWordsPerWLEN)-1:0] ispr_word_addr_base;
  logic [BaseWordsPerWLEN-1:0]         ispr_word_sel_base;

  ispr_e                               ispr_addr_bignum;

  logic                                ispr_wr_insn, ispr_rd_insn;
  logic                                ispr_wr_base_insn;
  logic                                ispr_wr_bignum_insn;
  logic                                ispr_rd_bignum_insn;

  logic                     lsu_load_req_raw;
  logic                     lsu_store_req_raw;
  logic [DmemAddrWidth-1:0] lsu_addr, lsu_addr_blanked, lsu_addr_saved_d, lsu_addr_saved_q;
  logic                     lsu_addr_saved_sel;
  logic                     expected_lsu_addr_en;

  logic                     expected_call_stack_push, expected_call_stack_pop;
  logic                     lsu_predec_error, branch_target_predec_error, ctrl_predec_error;

  logic rnd_req_raw;

  // Register read data with integrity stripped off
  logic [31:0]     rf_base_rd_data_a_no_intg;
  logic [31:0]     rf_base_rd_data_b_no_intg;
  logic [WLEN-1:0] rf_bignum_rd_data_a_no_intg;
  logic [WLEN-1:0] rf_bignum_rd_data_b_no_intg;

  logic [ExtWLEN-1:0] rf_bignum_rd_data_b_intg_blanked;
  logic [ExtWLEN-1:0] selection_result;

  logic [1:0] rf_bignum_wr_en_unbuf;
  logic [4:0] rf_bignum_wr_addr_unbuf;
  logic [4:0] rf_bignum_rd_addr_a_unbuf;
  logic       rf_bignum_rd_en_a_unbuf;
  logic [4:0] rf_bignum_rd_addr_b_unbuf;
  logic       rf_bignum_rd_en_b_unbuf;

  logic rf_bignum_rd_a_indirect_en;
  logic rf_bignum_rd_b_indirect_en;
  logic rf_bignum_wr_indirect_en;

  // Computed increments for indirect register index and memory address in BN.LID/BN.SID/BN.MOVR
  // instructions.
  logic [5:0]  rf_base_rd_data_a_inc;
  logic [5:0]  rf_base_rd_data_b_inc;
  logic [26:0] rf_base_rd_data_a_wlen_word_inc;

  // Read/Write enables for base register file before illegal instruction encoding are factored in
  logic rf_base_rd_en_a_raw, rf_base_rd_en_b_raw, rf_base_wr_en_raw;

  // Output of mux taking the above increments as inputs and choosing one to write back to base
  // register file with appropriate zero extension and padding to give a 32-bit result.
  logic [31:0]              increment_out;

  // Loop control, used to start a new loop
  logic        loop_start_req;
  logic        loop_start_commit;
  logic        loop_reset;
  logic [11:0] loop_bodysize;
  logic [31:0] loop_iterations;

  // Loop generated jumps. The loop controller asks to jump when execution reaches the end of a loop
  // body that hasn't completed all of its iterations.
  logic                     loop_jump;
  logic [ImemAddrWidth-1:0] loop_jump_addr;

  logic [WLEN-1:0] mac_bignum_rf_wr_data;

  logic loop_hw_err, loop_predec_err;
  logic csr_illegal_addr, wsr_illegal_addr, ispr_illegal_addr;
  logic imem_addr_err, loop_sw_err, ispr_err;
  logic dmem_addr_err_check, dmem_addr_err;
  logic dmem_addr_unaligned_base, dmem_addr_unaligned_bignum, dmem_addr_overflow;
  logic illegal_insn_static;
  logic key_invalid;

  logic rf_a_indirect_err, rf_b_indirect_err, rf_d_indirect_err, rf_indirect_err;

  // If we are doing an indirect access to the bignum register file, it's possible that the
  // address that we use for the access is architecturally unknown. This happens if it came from x1
  // and we've underflowed the call stack. When this happens, we want to ignore any read data
  // integrity errors and spurious write enable errors since the access to the bignum register file
  // didn't happen architecturally anyway.
  logic ignore_rf_bignum_intg_errs;
  logic rf_bignum_intg_err;
  logic ignore_rf_bignum_spurious_we_errs;
  logic rf_bignum_spurious_we_err;

  logic ispr_rdata_intg_err;

  logic [31:0] insn_cnt_d, insn_cnt_q;
  logic        insn_cnt_clear;

  logic [4:0] insn_bignum_rd_addr_a_q, insn_bignum_rd_addr_b_q, insn_bignum_wr_addr_q;

  logic       start_secure_wipe;
  logic       secure_wipe_running_q, secure_wipe_running_d;

  assign secure_wipe_running_d = start_secure_wipe | (secure_wipe_running_q & ~secure_wipe_ack_i);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      secure_wipe_running_q <= 1'b0;
    end else begin
      secure_wipe_running_q <= secure_wipe_running_d;
    end
  end
  assign secure_wipe_req_o = start_secure_wipe | secure_wipe_running_q;

  // Spot spurious acks on the secure wipe interface. There is a an ack at the end of the initial
  // secure wipe, and as `secure_wipe_running_q` is only high during secure wipes triggered by this
  // controller, we have to ignore acks before the initial secure wipe is done.  Register this
  // signal to break a circular path (a secure wipe can be triggered by a stop, and a spurious
  // secure wipe ack can trigger a stop).
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      spurious_secure_wipe_ack_q <= 1'b0;
    end else begin
      spurious_secure_wipe_ack_q <= spurious_secure_wipe_ack_d;
    end
  end
  assign spurious_secure_wipe_ack_d = spurious_secure_wipe_ack_q |
                                      (secure_wipe_ack_i      &
                                       ~secure_wipe_running_q &
                                       ~secure_wipe_running_i);

  // Stall a cycle on loads to allow load data writeback to happen the following cycle. Stall not
  // required on stores as there is no response to deal with.
  assign mem_stall = lsu_load_req_raw;

  // Reads to RND must stall until data is available
  assign ispr_stall = rnd_req_raw & ~rnd_valid_i;

  assign rf_indirect_stall = insn_valid_i &
                             (state_q != OtbnStateStall) &
                             (insn_dec_shared_i.subset == InsnSubsetBignum) &
                             (insn_dec_bignum_i.rf_a_indirect |
                              insn_dec_bignum_i.rf_b_indirect |
                              insn_dec_bignum_i.rf_d_indirect);

  assign stall = mem_stall | ispr_stall | rf_indirect_stall;

  // OTBN is done when it was executing something (in state OtbnStateRun or OtbnStateStall)
  // and either it executes an ecall or an error occurs. A pulse on the done signal raises the
  // 'done' interrupt and also tells the top-level to update its ERR_BITS status
  // register. The calculation that ecall triggered done is factored out as `done_complete` to
  // avoid logic loops in the error handling logic.
  assign done_complete = (insn_valid_i & insn_dec_shared_i.ecall_insn);
  assign executing = (state_q == OtbnStateRun) ||
                     (state_q == OtbnStateStall);

  // Set the *locking* output when the next state is the *locked* state and no secure wipe is
  // running or there is a URND reseed error.  `locking_o` is thus set only after the secure wipe
  // has completed or if it cannot complete due to an URND reseed error (in which case
  // `secure_wipe_req_o` and `urnd_reseed_err_i` will remain high).  The condition for secure wipe
  // running involves `secure_wipe_running_i`, which is high for the initial secure wipe, and
  // `secure_wipe_req_o`, which is high for post-execution secure wipes.
  assign locking_o = (state_d == OtbnStateLocked) & (~(secure_wipe_running_i | secure_wipe_req_o) |
                                                     urnd_reseed_err_i | mubi_err_d);

  assign start_secure_wipe = executing & (done_complete | err);

  assign jump_or_branch = (insn_valid_i &
                           (insn_dec_shared_i.branch_insn | insn_dec_shared_i.jump_insn));

  // Branch taken when there is a valid branch instruction and comparison passes or a valid jump
  // instruction (which is always taken)
  assign branch_taken = insn_valid_i &
                        ((insn_dec_shared_i.branch_insn & alu_base_comparison_result_i) |
                         insn_dec_shared_i.jump_insn);
  // Branch target computed by base ALU (PC + imm)
  assign branch_target = alu_base_operation_result_i[ImemAddrWidth-1:0];
  assign branch_target_overflow = |alu_base_operation_result_i[31:ImemAddrWidth];

  assign next_insn_addr_wide = {1'b0, insn_addr_i} + 'd4;
  assign next_insn_addr = next_insn_addr_wide[ImemAddrWidth-1:0];

  // Record address for fetch request so it can be retried when an invalid response is received
  always_ff @(posedge clk_i) begin
    if (insn_fetch_req_valid_raw) begin
      insn_fetch_req_addr_last <= insn_fetch_req_addr_o;
    end
  end

  always_comb begin
    state_d                  = state_q;
    // `insn_fetch_req_valid_raw` is the value `insn_fetch_req_valid_o` before any errors are
    // considered.
    insn_fetch_req_valid_raw = 1'b0;
    insn_fetch_req_addr_o    = '0;
    insn_fetch_resp_clear_o  = 1'b1;
    prefetch_en_o            = 1'b0;

    state_error = 1'b0;

    unique case (state_q)
      OtbnStateHalt: begin
        if (start_i) begin
          state_d = OtbnStateRun;

          insn_fetch_req_addr_o    = '0;
          insn_fetch_req_valid_raw = 1'b1;
          prefetch_en_o            = 1'b1;
        end
      end
      OtbnStateRun: begin
        insn_fetch_req_valid_raw = 1'b1;
        prefetch_en_o            = 1'b1;

        if (!insn_valid_i) begin
          insn_fetch_req_addr_o = insn_fetch_req_addr_last;
        end else if (done_complete) begin
          state_d                  = OtbnStateHalt;
          insn_fetch_req_valid_raw = 1'b0;
          prefetch_en_o            = 1'b0;
        end else begin
          if (stall) begin
            // When stalling don't request a new fetch and don't clear response either to keep
            // current instruction.
            state_d                  = OtbnStateStall;
            insn_fetch_req_valid_raw = 1'b0;
            insn_fetch_resp_clear_o  = 1'b0;
          end else begin
            if (branch_taken) begin
              insn_fetch_req_addr_o = branch_target;
            end else if (loop_jump) begin
              insn_fetch_req_addr_o = loop_jump_addr;
            end else begin
              insn_fetch_req_addr_o = next_insn_addr;
            end
          end
        end
      end
      OtbnStateStall: begin
        prefetch_en_o = 1'b1;
        // When stalling refetch the same instruction to keep decode inputs constant
        if (stall) begin
          state_d                  = OtbnStateStall;
          //insn_fetch_req_addr_o = insn_addr_i;
          insn_fetch_req_valid_raw = 1'b0;
          insn_fetch_resp_clear_o  = 1'b0;
        end else begin
          insn_fetch_req_valid_raw = 1'b1;

          if (loop_jump) begin
            insn_fetch_req_addr_o = loop_jump_addr;
          end else begin
            insn_fetch_req_addr_o = next_insn_addr;
          end

          state_d = OtbnStateRun;
        end
      end
      OtbnStateLocked: begin
        insn_fetch_req_valid_raw = 1'b0;
        state_d                  = OtbnStateLocked;
      end
      default: begin
        // We should never get here. If we do (e.g. via a malicious glitch), error out immediately.
        // SEC_CM: CONTROLLER.FSM.LOCAL_ESC
        state_d = OtbnStateLocked;
        state_error = 1'b1;
      end
    endcase

    // On any error immediately halt, either going to OtbnStateLocked or OtbnStateHalt depending on
    // whether it was a fatal error.
    if (err) begin
      prefetch_en_o           = 1'b0;
      insn_fetch_resp_clear_o = 1'b1;

      if (fatal_err) begin
        // SEC_CM: CONTROLLER.FSM.GLOBAL_ESC
        state_d = OtbnStateLocked;
      end else begin
        state_d = OtbnStateHalt;
      end
    end

    // Regardless of what happens above enforce staying in OtnbStateLocked.
    if (state_q == OtbnStateLocked) begin
      state_d = OtbnStateLocked;
    end
  end

  assign state_error_d = state_error | state_error_q;

  prim_flop #(
    .Width(1),
    .ResetValue('0)
  ) u_state_error_flop (
    .clk_i,
    .rst_ni,

    .d_i(state_error_d),
    .q_o(state_error_q)
  );

  `ASSERT(InsnAlwaysValidInStall, state_q == OtbnStateStall |-> insn_valid_i)

  // Anything that moves us or keeps us in the stall state should cause `stall` to be asserted
  `ASSERT(StallIfNextStateStall, insn_valid_i & (state_d == OtbnStateStall) |-> stall)

  // The raw signal is needed by the instruction fetch stage for generating instruction address
  // errors (where instruction fetch and prefetch disagree on address). `err` will factor this in so
  // using the qualified signal results in a combinational loop.
  assign insn_fetch_req_valid_raw_o = insn_fetch_req_valid_raw;
  assign insn_fetch_req_valid_o     = err ? 1'b0 : insn_fetch_req_valid_raw;

  // Determine if there are any errors related to the Imem fetch address.
  always_comb begin
    imem_addr_err = 1'b0;

    if (insn_fetch_req_valid_raw) begin
      if (|insn_fetch_req_addr_o[1:0]) begin
        // Imem address is unaligned
        imem_addr_err = 1'b1;
      end else if (branch_taken) begin
        imem_addr_err = branch_target_overflow;
      end else begin
        imem_addr_err = next_insn_addr_wide[ImemAddrWidth] & insn_valid_i;
      end
    end
  end

  // Signal error if MuBi input signals take on invalid values as this means something bad is
  // happening. Register the error signal to break circular paths (instruction fetch errors factor
  // into fatal_escalate_en_i, RND errors factor into recov_escalate_en_i).
  assign mubi_err_d = |{mubi4_test_invalid(fatal_escalate_en_i),
                        mubi4_test_invalid(recov_escalate_en_i),
                        mubi4_test_invalid(rma_req_i),
                        mubi_err_q};
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      mubi_err_q <= 1'b0;
    end else begin
      mubi_err_q <= mubi_err_d;
    end
  end

  // Instruction is illegal based on the static properties of the instruction bits (illegal encoding
  // or illegal WSR/CSR referenced).
  assign illegal_insn_static = insn_illegal_i | ispr_err;

  assign fatal_software_err       = software_err & software_errs_fatal_i;
  assign bad_internal_state_err   = |{state_error_d, loop_hw_err, rf_base_call_stack_hw_err_i,
                                      rf_bignum_spurious_we_err, spurious_secure_wipe_ack_q,
                                      mubi_err_q};
  assign reg_intg_violation_err   = rf_bignum_intg_err | ispr_rdata_intg_err;
  assign key_invalid_err          = ispr_rd_bignum_insn & insn_valid_i & key_invalid;
  assign illegal_insn_err         = illegal_insn_static | rf_indirect_err;
  assign call_stack_sw_err        = rf_base_call_stack_sw_err_i;

  // Flag a bad data address error if the data memory address is invalid and it does not come from
  // an empty call stack.  The second case cannot be decided as bad data address because the address
  // on top of the empty call stack may or may not be valid.  (Also, in most RTL simulators an empty
  // call stack that has never been pushed contains an unknown value, so this error bit would become
  // unknown.)  Thus, a data memory address coming from an empty call stack raises a call stack
  // error but never a bad data address error.
  assign bad_data_addr_err = dmem_addr_err &
                             ~(call_stack_sw_err &
                               (ld_insn_with_addr_from_call_stack |
                                st_insn_with_addr_from_call_stack));

  // Identify load instructions that take the memory address from the call stack.
  assign ld_insn_with_addr_from_call_stack = insn_valid_i               &
                                             insn_dec_shared_i.ld_insn  &
                                             insn_dec_base_i.rf_ren_a   &
                                             (insn_dec_base_i.a == 5'd1);

  // Identify store instructions that take the memory address from the call stack.
  assign st_insn_with_addr_from_call_stack = insn_valid_i               &
                                             insn_dec_shared_i.st_insn  &
                                             insn_dec_base_i.rf_ren_a   &
                                             (insn_dec_base_i.a == 5'd1);

  // All software errors that aren't bad_insn_addr. Factored into bad_insn_addr so it is only raised
  // if other software errors haven't ocurred. As bad_insn_addr relates to the next instruction
  // begin fetched it cannot occur if the current instruction has seen an error and failed to
  // execute.
  assign non_insn_addr_software_err = |{key_invalid_err,
                                        loop_sw_err,
                                        illegal_insn_err,
                                        call_stack_sw_err,
                                        bad_data_addr_err};

  assign bad_insn_addr_err = imem_addr_err & ~non_insn_addr_software_err;

  assign err_bits_d = '{
    fatal_software:     fatal_software_err,
    bad_internal_state: bad_internal_state_err,
    reg_intg_violation: reg_intg_violation_err,
    key_invalid:        key_invalid_err,
    loop:               loop_sw_err,
    illegal_insn:       illegal_insn_err,
    call_stack:         call_stack_sw_err,
    bad_data_addr:      bad_data_addr_err,
    bad_insn_addr:      bad_insn_addr_err
  };

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_bits_q <= '0;
    end else begin
      if (err_bit_clear_i && !locking_o) begin
        err_bits_q <= '0;
      end else begin
        err_bits_q <= err_bits_q | err_bits_d;
      end
    end
  end
  assign err_bits_o = err_bits_q;

  assign software_err = non_insn_addr_software_err | bad_insn_addr_err;

  assign recoverable_err = mubi4_test_true_loose(recov_escalate_en_i);

  assign internal_fatal_err = |{fatal_software_err,
                                bad_internal_state_err,
                                reg_intg_violation_err};

  // In case of an RMA request, just lock up the controller. This triggers the rotation of the
  // scrambling keys. The start/stop controller takes care of initiating the internal secure wipe
  // and eventually acknowledging the RMA request.
  assign fatal_err = |{internal_fatal_err,
                       mubi4_test_true_loose(fatal_escalate_en_i),
                       mubi4_test_true_loose(rma_req_i)};

  assign recoverable_err_o = recoverable_err | (software_err & ~software_errs_fatal_i);
  assign mems_sec_wipe_o   = (state_d == OtbnStateLocked) & (state_q != OtbnStateLocked);

  assign internal_err = software_err | internal_fatal_err;
  assign err          = software_err | recoverable_err | fatal_err;

  assign prefetch_ignore_errs_o = internal_err;

  // Instructions must not execute if there is an error
  assign insn_executing = insn_valid_i & ~err;

  `ASSERT(ErrBitSetOnErr,
      err & (mubi4_test_false_strict(fatal_escalate_en_i) &
             mubi4_test_false_strict(recov_escalate_en_i) &
             mubi4_test_false_strict(rma_req_i)) |=>
          err_bits_o)
  `ASSERT(ErrSetOnFatalErr, fatal_err |-> err)
  `ASSERT(SoftwareErrIfNonInsnAddrSoftwareErr, non_insn_addr_software_err |-> software_err)

  `ASSERT(ControllerStateValid,
          state_q inside {OtbnStateHalt, OtbnStateRun, OtbnStateStall, OtbnStateLocked})
  // Branch only takes effect in OtbnStateRun so must not go into stall state for branch
  // instructions.
  `ASSERT(NoStallOnBranch,
      insn_valid_i & insn_dec_shared_i.branch_insn |-> state_q != OtbnStateStall)

  // SEC_CM: CONTROLLER.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, otbn_state_e, OtbnStateHalt)

  // SEC_CM: CTRL_FLOW.COUNT
  assign insn_cnt_clear = state_reset_i | (state_q == OtbnStateLocked) | insn_cnt_clear_i;

  always_comb begin
    if (insn_cnt_clear) begin
      insn_cnt_d = 32'd0;
    end else if (insn_executing & ~stall & (insn_cnt_q != 32'hffffffff)) begin
      insn_cnt_d = insn_cnt_q + 32'd1;
    end else begin
      insn_cnt_d = insn_cnt_q;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      insn_cnt_q <= 32'd0;
    end else begin
      insn_cnt_q <= insn_cnt_d;
    end
  end

  assign insn_cnt_o = insn_cnt_q;

  assign loop_reset = state_reset_i | sec_wipe_zero_i;

  otbn_loop_controller #(
    .ImemAddrWidth(ImemAddrWidth)
  ) u_otbn_loop_controller (
    .clk_i,
    .rst_ni,

    .state_reset_i(loop_reset),

    .insn_valid_i,
    .insn_addr_i,
    .next_insn_addr_i(next_insn_addr),

    .loop_start_req_i       (loop_start_req),
    .loop_start_commit_i    (loop_start_commit),
    .loop_bodysize_i        (loop_bodysize),
    .loop_iterations_i      (loop_iterations),
    .loop_end_addr_predec_i (ctrl_flow_target_predec_i),

    .loop_jump_o     (loop_jump),
    .loop_jump_addr_o(loop_jump_addr),

    .sw_err_o     (loop_sw_err),
    .hw_err_o     (loop_hw_err),
    .predec_err_o (loop_predec_err),

    .jump_or_branch_i(jump_or_branch),
    .otbn_stall_i    (stall),

    .prefetch_loop_active_o,
    .prefetch_loop_iterations_o,
    .prefetch_loop_end_addr_o,
    .prefetch_loop_jump_addr_o
  );

  // loop_start_req indicates the instruction wishes to start a loop, loop_start_commit confirms it
  // should occur.
  assign loop_start_req    = insn_valid_i & insn_dec_shared_i.loop_insn;
  assign loop_start_commit = insn_executing;
  assign loop_bodysize     = insn_dec_base_i.loop_bodysize;
  assign loop_iterations   = insn_dec_base_i.loop_immediate ? insn_dec_base_i.i :
                                                              rf_base_rd_data_a_no_intg;

  // Compute increments which can be optionally applied to indirect register accesses and memory
  // addresses in BN.LID/BN.SID/BN.MOVR instructions.
  assign rf_base_rd_data_a_inc           = rf_base_rd_data_a_no_intg[4:0] + 1'b1;
  assign rf_base_rd_data_b_inc           = rf_base_rd_data_b_no_intg[4:0] + 1'b1;
  // We can avoid a full 32-bit adder here because the offset is 32-bit aligned, so we know the
  // load/store address will only be valid if rf_base_rd_data_a_no_intg[4:0] is zero.
  assign rf_base_rd_data_a_wlen_word_inc = rf_base_rd_data_a_no_intg[31:5] + 27'h1;

  // Choose increment to write back to base register file, only one increment can be written as
  // there is only one write port. Note that where an instruction is incrementing the indirect
  // reference to its destination register (insn_dec_bignum_i.d_inc) that reference is read on the
  // B read port so the B increment is written back.
  always_comb begin
    unique case (1'b1)
      insn_dec_bignum_i.a_inc: begin
        increment_out = {26'b0, rf_base_rd_data_a_inc};
      end
      insn_dec_bignum_i.b_inc: begin
        increment_out = {26'b0, rf_base_rd_data_b_inc};
      end
      insn_dec_bignum_i.d_inc: begin
        increment_out = {26'b0, rf_base_rd_data_b_inc};
      end
      insn_dec_bignum_i.a_wlen_word_inc: begin
        increment_out = {rf_base_rd_data_a_wlen_word_inc, 5'b0};
      end
      default: begin
        // Whenever increment_out is written back to the register file, exactly one of the
        // increment selector signals is high. To prevent the automatic inference of latches in
        // case nothing is written back (rf_wdata_sel != RfWdSelIncr) and to save logic, we choose
        // a valid output as default.
        increment_out = {26'b0, rf_base_rd_data_a_inc};
      end
    endcase
  end

  // Base RF read/write address, enable and commit control
  always_comb begin
    rf_base_rd_addr_a_o = insn_dec_base_i.a;
    rf_base_rd_addr_b_o = insn_dec_base_i.b;
    rf_base_wr_addr_o   = insn_dec_base_i.d;

    // Only commit read or write if the instruction is executing (in particular a read commit pops
    // the call stack so must not occur where a valid instruction sees an error and doesn't
    // execute).
    rf_base_rd_commit_o = insn_executing;
    rf_base_wr_commit_o = insn_executing;

    rf_base_rd_en_a_raw = 1'b0;
    rf_base_rd_en_b_raw = 1'b0;
    rf_base_wr_en_raw   = 1'b0;

    if (insn_valid_i) begin
      if (insn_dec_shared_i.st_insn) begin
        // For stores, both base reads happen in the first cycle of the store instruction. For base
        // stores this is the same cycle as the request. For bignum stores this is the cycle before
        // the request (as the indirect register read to get the store data occurs the following
        // cycle).
        rf_base_rd_en_a_raw = insn_dec_base_i.rf_ren_a &
          (rf_indirect_stall | (insn_dec_shared_i.subset == InsnSubsetBase));
        rf_base_rd_en_b_raw = insn_dec_base_i.rf_ren_b &
          (rf_indirect_stall | (insn_dec_shared_i.subset == InsnSubsetBase));

        // Bignum stores can update the base register file where an increment is used.
        rf_base_wr_en_raw   = (insn_dec_shared_i.subset == InsnSubsetBignum) &
                              insn_dec_base_i.rf_we                          &
                              rf_indirect_stall;
      end else if (insn_dec_shared_i.ld_insn) begin
        // For loads, both base reads happen in the same cycle as the request. The address is
        // required for the request and the indirect destination register (only used for Bignum
        // loads) is flopped in ld_insn_bignum_wr_addr_q to correctly deal with the case where it's
        // updated by an increment.
        rf_base_rd_en_a_raw = insn_dec_base_i.rf_ren_a & lsu_load_req_raw;
        rf_base_rd_en_b_raw = insn_dec_base_i.rf_ren_b & lsu_load_req_raw;

        if (insn_dec_shared_i.subset == InsnSubsetBignum) begin
          // Bignum loads can update the base register file where an increment is used. This must
          // always happen in the same cycle as the request as this is where both registers are
          // read.
          rf_base_wr_en_raw = insn_dec_base_i.rf_we & lsu_load_req_raw & rf_indirect_stall;
        end else begin
          // For Base loads write the base register file when the instruction is unstalled (meaning
          // the load data is available).
          rf_base_wr_en_raw = insn_dec_base_i.rf_we & ~stall;
        end
      end else if (insn_dec_bignum_i.rf_wdata_sel == RfWdSelMovSel) begin
        // For MOVR base register reads occur in the first cycle of the instruction. The indirect
        // register read for the bignum data occurs in the following cycle.
        rf_base_rd_en_a_raw = insn_dec_base_i.rf_ren_a & rf_indirect_stall;
        rf_base_rd_en_b_raw = insn_dec_base_i.rf_ren_b & rf_indirect_stall;
        rf_base_wr_en_raw   = insn_dec_base_i.rf_we    & rf_indirect_stall;
      end else begin
        // For all other instructions the read and write happen when the instruction is unstalled.
        rf_base_rd_en_a_raw = insn_dec_base_i.rf_ren_a & ~stall;
        rf_base_rd_en_b_raw = insn_dec_base_i.rf_ren_b & ~stall;
        rf_base_wr_en_raw   = insn_dec_base_i.rf_we    & ~stall;
      end
    end

    if (insn_dec_shared_i.subset == InsnSubsetBignum) begin
      unique case (1'b1)
        insn_dec_bignum_i.a_inc,
        insn_dec_bignum_i.a_wlen_word_inc: begin
          rf_base_wr_addr_o = insn_dec_base_i.a;
        end

        insn_dec_bignum_i.b_inc,
        insn_dec_bignum_i.d_inc: begin
          rf_base_wr_addr_o = insn_dec_base_i.b;
        end
        default: ;
      endcase
    end

    rf_base_rd_en_a_o = rf_base_rd_en_a_raw & ~illegal_insn_static;
    rf_base_rd_en_b_o = rf_base_rd_en_b_raw & ~illegal_insn_static;
    rf_base_wr_en_o   = rf_base_wr_en_raw   & ~illegal_insn_static;
  end

  // Base ALU Operand A MUX
  always_comb begin
    unique case (insn_dec_base_i.op_a_sel)
      OpASelRegister: alu_base_operation_o.operand_a = rf_base_rd_data_a_no_intg;
      OpASelZero:     alu_base_operation_o.operand_a = '0;
      OpASelCurrPc:   alu_base_operation_o.operand_a = {{(32 - ImemAddrWidth){1'b0}}, insn_addr_i};
      default:        alu_base_operation_o.operand_a = rf_base_rd_data_a_no_intg;
    endcase
  end

  // Base ALU Operand B MUX
  always_comb begin
    unique case (insn_dec_base_i.op_b_sel)
      OpBSelRegister:  alu_base_operation_o.operand_b = rf_base_rd_data_b_no_intg;
      OpBSelImmediate: alu_base_operation_o.operand_b = insn_dec_base_i.i;
      default:         alu_base_operation_o.operand_b = rf_base_rd_data_b_no_intg;
    endcase
  end

  assign alu_base_operation_o.op = insn_dec_base_i.alu_op;

  assign alu_base_comparison_o.operand_a = rf_base_rd_data_a_no_intg;
  assign alu_base_comparison_o.operand_b = rf_base_rd_data_b_no_intg;
  assign alu_base_comparison_o.op = insn_dec_base_i.comparison_op;

  assign rf_base_rd_data_a_no_intg = rf_base_rd_data_a_intg_i[31:0];
  assign rf_base_rd_data_b_no_intg = rf_base_rd_data_b_intg_i[31:0];

  logic unused_rf_base_rd_a_intg_bits;

  // TODO(#18266): Implement GPR to ISPR end to end integrity path (ISPR writes from GPR take data
  // from base RF port A)
  assign unused_rf_base_rd_a_intg_bits = |rf_base_rd_data_a_intg_i[38:32];

  // Base register file write MUX. Depending on the data source, integrity bits do or don't have to
  // be appended:
  // - Data sources that require appending integrity bits go into `rf_base_wr_data_no_intg_o` and
  //   `rf_base_wr_data_intg_sel_o` is low.
  // - Data sources that already come with integrity bits go into `rf_base_wr_data_intg_o` and
  //   `rf_base_wr_data_intg_sel_o` is high.
  always_comb begin
    // Default values
    rf_base_wr_data_no_intg_o  = alu_base_operation_result_i;
    rf_base_wr_data_intg_o     = '0;
    rf_base_wr_data_intg_sel_o = 1'b0;

    unique case (insn_dec_base_i.rf_wdata_sel)
      RfWdSelEx: begin
        rf_base_wr_data_no_intg_o  = alu_base_operation_result_i;
      end
      RfWdSelNextPc: begin
        rf_base_wr_data_no_intg_o  = {{(32-(ImemAddrWidth+1)){1'b0}}, next_insn_addr_wide};
      end
      RfWdSelIspr: begin
        rf_base_wr_data_no_intg_o  = csr_rdata;
      end
      RfWdSelIncr: begin
        rf_base_wr_data_no_intg_o  = increment_out;
      end
      RfWdSelLsu: begin
        rf_base_wr_data_intg_sel_o = 1'b1;
        rf_base_wr_data_intg_o     = lsu_base_rdata_i;
      end
      default: ;
    endcase
  end

  for (genvar i = 0; i < BaseWordsPerWLEN; ++i) begin : g_rf_bignum_rd_data
    assign rf_bignum_rd_data_a_no_intg[i*32+:32] = rf_bignum_rd_data_a_intg_i[i*39+:32];
    assign rf_bignum_rd_data_b_no_intg[i*32+:32] = rf_bignum_rd_data_b_intg_i[i*39+:32];
  end

  // Bignum RF control signals from the controller aren't actually used, instead the predecoded
  // one-hot versions are. The predecoded versions get checked against the signals produced here.
  // Buffer them to ensure they don't get optimised away (with a functionaly correct OTBN they will
  // always be identical).
  assign rf_bignum_rd_addr_a_unbuf = insn_dec_bignum_i.rf_a_indirect ? insn_bignum_rd_addr_a_q :
                                                                       insn_dec_bignum_i.a;

  prim_buf #(
    .Width(WdrAw)
  ) u_rf_bignum_rd_addr_a_buf (
    .in_i (rf_bignum_rd_addr_a_unbuf),
    .out_o(rf_bignum_rd_addr_a_o)
  );

  assign rf_bignum_rd_en_a_unbuf = insn_dec_bignum_i.rf_ren_a & insn_valid_i & ~stall;

  prim_buf #(
    .Width(1)
  ) u_rf_bignum_rd_en_a_buf (
    .in_i (rf_bignum_rd_en_a_unbuf),
    .out_o(rf_bignum_rd_en_a_o)
  );

  assign rf_bignum_rd_addr_b_unbuf = insn_dec_bignum_i.rf_b_indirect ? insn_bignum_rd_addr_b_q :
                                                                       insn_dec_bignum_i.b;

  prim_buf #(
    .Width(WdrAw)
  ) u_rf_bignum_rd_addr_b_buf (
    .in_i (rf_bignum_rd_addr_b_unbuf),
    .out_o(rf_bignum_rd_addr_b_o)
  );

  assign rf_bignum_rd_en_b_unbuf = insn_dec_bignum_i.rf_ren_b & insn_valid_i & ~stall;

  prim_buf #(
    .Width(1)
  ) u_rf_bignum_rd_en_b_buf (
    .in_i (rf_bignum_rd_en_b_unbuf),
    .out_o(rf_bignum_rd_en_b_o)
  );

  assign alu_bignum_operation_o.operand_a = rf_bignum_rd_data_a_no_intg;

  // Base ALU Operand B MUX
  always_comb begin
    unique case (insn_dec_bignum_i.alu_op_b_sel)
      OpBSelRegister:  alu_bignum_operation_o.operand_b = rf_bignum_rd_data_b_no_intg;
      OpBSelImmediate: alu_bignum_operation_o.operand_b = insn_dec_bignum_i.i;
      default:         alu_bignum_operation_o.operand_b = rf_bignum_rd_data_b_no_intg;
    endcase
  end

  assign alu_bignum_operation_o.op          = insn_dec_bignum_i.alu_op;
  assign alu_bignum_operation_o.shift_right = insn_dec_bignum_i.alu_shift_right;
  assign alu_bignum_operation_o.shift_amt   = insn_dec_bignum_i.alu_shift_amt;
  assign alu_bignum_operation_o.flag_group  = insn_dec_bignum_i.alu_flag_group;
  assign alu_bignum_operation_o.sel_flag    = insn_dec_bignum_i.alu_sel_flag;
  assign alu_bignum_operation_o.alu_flag_en = insn_dec_bignum_i.alu_flag_en & insn_valid_i;
  assign alu_bignum_operation_o.mac_flag_en = insn_dec_bignum_i.mac_flag_en & insn_valid_i;

  assign alu_bignum_operation_valid_o  = insn_valid_i;
  assign alu_bignum_operation_commit_o = insn_executing;

  assign mac_bignum_operation_o.operand_a         = rf_bignum_rd_data_a_no_intg;
  assign mac_bignum_operation_o.operand_b         = rf_bignum_rd_data_b_no_intg;
  assign mac_bignum_operation_o.operand_a_qw_sel  = insn_dec_bignum_i.mac_op_a_qw_sel;
  assign mac_bignum_operation_o.operand_b_qw_sel  = insn_dec_bignum_i.mac_op_b_qw_sel;
  assign mac_bignum_operation_o.wr_hw_sel_upper   = insn_dec_bignum_i.mac_wr_hw_sel_upper;
  assign mac_bignum_operation_o.pre_acc_shift_imm = insn_dec_bignum_i.mac_pre_acc_shift;
  assign mac_bignum_operation_o.zero_acc          = insn_dec_bignum_i.mac_zero_acc;
  assign mac_bignum_operation_o.shift_acc         = insn_dec_bignum_i.mac_shift_out;

  assign mac_bignum_en_o     = insn_valid_i & insn_dec_bignum_i.mac_en;
  assign mac_bignum_commit_o = insn_executing;

  // Move / Conditional Select. Only select B register data when a selection instruction is being
  // executed and the selection flag isn't set. To avoid undesirable SCA leakage between the two
  // registers for non-selection instructions, the B register is blanked except for selection
  // instructions.
  // Note that blanking both registers is not feasible nor absolutely required because:
  // - The flag group selection and flag selection are known in the predecoder stage but the actual
  //   flag isn't.
  // - Selecting the flag in the predocder stage using combinatorial inputs may lead to SCA leakage
  //   between the still combinatorial flag groups and flags within a group which might be
  //   undesirable as well.
  // - When executing a selection instruction, programmers can expected that there will be some SCA
  //   leakage between the two options. But it may be much lesse expected for such leakage to occur
  //   for other instructions.
  `ASSERT(SelFlagValid, insn_valid_i & insn_dec_bignum_i.sel_insn |->
    insn_dec_bignum_i.alu_sel_flag inside {FlagC, FlagL, FlagM, FlagZ})

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(ExtWLEN)) u_rf_bignum_rd_data_b_intg_blanker (
    .in_i (rf_bignum_rd_data_b_intg_i),
    .en_i (ctrl_flow_predec_i.sel_insn),
    .out_o(rf_bignum_rd_data_b_intg_blanked)
  );

  `ASSERT(BlankingBignumRdDataBSel,
    ~(insn_valid_i & insn_dec_bignum_i.sel_insn) |-> rf_bignum_rd_data_b_intg_blanked == '0,
    clk_i, !rst_ni || ctrl_predec_error || !insn_executing)

  assign selection_result =
    ~ctrl_flow_predec_i.sel_insn | alu_bignum_selection_flag_i ? rf_bignum_rd_data_a_intg_i :
                                                                 rf_bignum_rd_data_b_intg_blanked;

  // Bignum Register file write control

  always_comb begin
    // By default write nothing
    rf_bignum_wr_en_unbuf = 2'b00;

    // Only write if valid instruction wants a bignum rf write and it isn't stalled. If instruction
    // doesn't execute (e.g. due to an error) the write won't commit.
    if (insn_valid_i && insn_dec_bignum_i.rf_we && !rf_indirect_stall) begin
      if (insn_dec_bignum_i.mac_en && insn_dec_bignum_i.mac_shift_out) begin
        // Special handling for BN.MULQACC.SO, only enable upper or lower half depending on
        // mac_wr_hw_sel_upper.
        rf_bignum_wr_en_unbuf = insn_dec_bignum_i.mac_wr_hw_sel_upper ? 2'b10 : 2'b01;
      end else begin
        // For everything else write both halves immediately.
        rf_bignum_wr_en_unbuf = 2'b11;
      end
    end
  end

  // Bignum RF control signals from the controller aren't actually used, instead the predecoded
  // one-hot versions are. The predecoded versions get checked against the signals produced here.
  // Buffer them to ensure they don't get optimised away (with a functionaly correct OTBN they will
  // always be identical).
  prim_buf #(
    .Width(2)
  ) u_bignum_wr_en_buf (
    .in_i (rf_bignum_wr_en_unbuf),
    .out_o(rf_bignum_wr_en_o)
  );


  assign rf_bignum_wr_commit_o = |rf_bignum_wr_en_o & insn_executing & !stall;

  assign rf_bignum_indirect_en_o    = insn_executing & rf_indirect_stall;
  assign rf_bignum_rd_a_indirect_en = insn_executing & insn_dec_bignum_i.rf_a_indirect;
  assign rf_bignum_rd_b_indirect_en = insn_executing & insn_dec_bignum_i.rf_b_indirect;
  assign rf_bignum_wr_indirect_en   = insn_executing & insn_dec_bignum_i.rf_d_indirect;

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_bignum_rd_a_idirect_onehot__enc (
    .in_i  (rf_base_rd_data_a_no_intg[4:0]),
    .en_i  (rf_bignum_rd_a_indirect_en),
    .out_o (rf_bignum_rd_a_indirect_onehot_o)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_bignum_rd_b_indirect_onehot_enc (
    .in_i  (rf_base_rd_data_b_no_intg[4:0]),
    .en_i  (rf_bignum_rd_b_indirect_en),
    .out_o (rf_bignum_rd_b_indirect_onehot_o)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_bignum_wr_indirect_onehot_enc (
    .in_i  (rf_base_rd_data_b_no_intg[4:0]),
    .en_i  (rf_bignum_wr_indirect_en),
    .out_o (rf_bignum_wr_indirect_onehot_o)
  );

  // For BN.LID sample the indirect destination register index in first cycle as an increment might
  // change it for the second cycle where the load data is written to the bignum register file.
  always_ff @(posedge clk_i) begin
    if (insn_dec_bignum_i.rf_d_indirect) begin
      insn_bignum_wr_addr_q <= rf_base_rd_data_b_no_intg[4:0];
    end

    if (insn_dec_bignum_i.rf_a_indirect) begin
      insn_bignum_rd_addr_a_q <= rf_base_rd_data_a_no_intg[4:0];
    end

    if (insn_dec_bignum_i.rf_b_indirect) begin
      insn_bignum_rd_addr_b_q <= rf_base_rd_data_b_no_intg[4:0];
    end
  end

  // Bignum RF control signals from the controller aren't actually used, instead the predecoded
  // one-hot versions are. The predecoded versions get checked against the signals produced here.
  // Buffer them to ensure they don't get optimised away (with a functionaly correct OTBN they will
  // always be identical).
  assign rf_bignum_wr_addr_unbuf = insn_dec_bignum_i.rf_d_indirect ? insn_bignum_wr_addr_q :
                                                                     insn_dec_bignum_i.d;

  prim_buf #(
    .Width(WdrAw)
  ) u_rf_bignum_wr_addr_buf (
    .in_i (rf_bignum_wr_addr_unbuf),
    .out_o(rf_bignum_wr_addr_o)
  );

  // For the shift-out variant of BN.MULQACC the bottom half of the MAC result is written to one
  // half of a desintation register specified by the instruction (mac_wr_hw_sel_upper). The bottom
  // half of the MAC result must be placed in the appropriate half of the write data (the RF only
  // accepts write data for the top half in the top half of the write data input). Otherwise
  // (shift-out to bottom half and all other BN.MULQACC instructions) simply pass the MAC result
  // through unchanged as write data.
  assign mac_bignum_rf_wr_data[WLEN-1:WLEN/2] =
      insn_dec_bignum_i.mac_wr_hw_sel_upper &&
      insn_dec_bignum_i.mac_shift_out          ? mac_bignum_operation_result_i[WLEN/2-1:0] :
                                                 mac_bignum_operation_result_i[WLEN-1:WLEN/2];

  assign mac_bignum_rf_wr_data[WLEN/2-1:0] = mac_bignum_operation_result_i[WLEN/2-1:0];

  // Bignum register file write MUX. Depending on the data source, integrity bits do or don't have
  // to be appended; see comments on the "Base register file write MUX" for details.
  always_comb begin
    // Default values
    rf_bignum_wr_data_intg_sel_o = 1'b0;
    rf_bignum_wr_data_intg_o     = '0;
    rf_bignum_wr_data_no_intg_o  = alu_bignum_operation_result_i;

    unique case (insn_dec_bignum_i.rf_wdata_sel)
      RfWdSelEx: begin
        rf_bignum_wr_data_no_intg_o  = alu_bignum_operation_result_i;
      end
      RfWdSelMac: begin
        rf_bignum_wr_data_no_intg_o  = mac_bignum_rf_wr_data;
      end
      RfWdSelIspr: begin
        rf_bignum_wr_data_intg_sel_o = 1'b1;
        rf_bignum_wr_data_intg_o     = ispr_rdata_intg_i;
      end
      RfWdSelMovSel: begin
        rf_bignum_wr_data_intg_sel_o = 1'b1;
        rf_bignum_wr_data_intg_o     = selection_result;
      end
      RfWdSelLsu: begin
        rf_bignum_wr_data_intg_sel_o = 1'b1;
        //SEC_CM: BUS.INTEGRITY
        rf_bignum_wr_data_intg_o     = lsu_bignum_rdata_i;
      end
      default: ;
    endcase
  end

  assign rf_a_indirect_err = insn_dec_bignum_i.rf_a_indirect    &
                             (|rf_base_rd_data_a_no_intg[31:5]) &
                             ~rf_base_call_stack_sw_err_i       &
                             rf_base_rd_en_a_o;

  assign rf_b_indirect_err = insn_dec_bignum_i.rf_b_indirect    &
                             (|rf_base_rd_data_b_no_intg[31:5]) &
                             ~rf_base_call_stack_sw_err_i       &
                             rf_base_rd_en_b_o;

  assign rf_d_indirect_err = insn_dec_bignum_i.rf_d_indirect    &
                             (|rf_base_rd_data_b_no_intg[31:5]) &
                             ~rf_base_call_stack_sw_err_i       &
                             rf_base_rd_en_b_o;

  assign rf_indirect_err =
      insn_valid_i & (rf_a_indirect_err | rf_b_indirect_err | rf_d_indirect_err);


  // If the source registers are indirectly indexed and there is a stack error, the source
  // register indices were illegal due to a stack pop error. In this case, ignore bignum RF read
  // integrity errors.
  assign ignore_rf_bignum_intg_errs = (insn_dec_bignum_i.rf_a_indirect |
                                       insn_dec_bignum_i.rf_b_indirect) &
                                      rf_base_call_stack_sw_err_i;

  assign rf_bignum_intg_err = rf_bignum_intg_err_i & ~ignore_rf_bignum_intg_errs;

  // If the destination register is indirectly indexed and there is a stack error, the destination
  // register index was illegal due to a stack pop error. In this case, ignore bignum RF
  // write-enable errors.
  assign ignore_rf_bignum_spurious_we_errs = insn_dec_bignum_i.rf_d_indirect &
                                             rf_base_call_stack_sw_err_i;

  assign rf_bignum_spurious_we_err = rf_bignum_spurious_we_err_i &
                                     ~ignore_rf_bignum_spurious_we_errs;

  // CSR/WSR/ISPR handling
  // ISPRs (Internal Special Purpose Registers) are the internal registers. CSRs and WSRs are the
  // ISA visible versions of those registers in the base and bignum ISAs respectively.

  assign csr_addr     = csr_e'(insn_dec_base_i.i[11:0]);
  assign csr_sub_addr = insn_dec_base_i.i[$clog2(BaseWordsPerWLEN)-1:0];

  always_comb begin
    ispr_addr_base      = IsprMod;
    ispr_word_addr_base = '0;
    csr_illegal_addr    = 1'b0;

    unique case (csr_addr)
      CsrFlags, CsrFg0, CsrFg1: begin
        ispr_addr_base      = IsprFlags;
        ispr_word_addr_base = '0;
      end
      CsrMod0, CsrMod1, CsrMod2, CsrMod3, CsrMod4, CsrMod5, CsrMod6, CsrMod7: begin
        ispr_addr_base      = IsprMod;
        ispr_word_addr_base = csr_sub_addr;
      end
      CsrRndPrefetch: begin
        // Reading from RND_PREFETCH results in 0, there is no ISPR to read so no address is set.
        // The csr_rdata mux logic takes care of producing the 0.
      end
      CsrRnd: begin
        ispr_addr_base      = IsprRnd;
        ispr_word_addr_base = '0;
      end
      CsrUrnd: begin
        ispr_addr_base      = IsprUrnd;
        ispr_word_addr_base = '0;
      end
      default: csr_illegal_addr = 1'b1;
    endcase
  end

  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_ispr_word_sel_base
    assign ispr_word_sel_base[i_word] = ispr_word_addr_base == i_word;
  end

  // Decode wide ISPR read data.
  logic [WLEN-1:0]                ispr_rdata;
  logic [2*BaseWordsPerWLEN-1:0]  ispr_rdata_intg_err_wide;
  logic [BaseWordsPerWLEN-1:0]    ispr_rdata_intg_err_narrow;
  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_ispr_rdata_dec
    prim_secded_inv_39_32_dec i_secded_dec (
      .data_i     (ispr_rdata_intg_i[i_word*39+:39]),
      .data_o     (/* unused because we abort on any integrity error */),
      .syndrome_o (/* unused */),
      .err_o      (ispr_rdata_intg_err_wide[i_word*2+:2])
    );
    assign ispr_rdata[i_word*32+:32] = ispr_rdata_intg_i[i_word*39+:32];
    assign ispr_rdata_intg_err_narrow[i_word] = |(ispr_rdata_intg_err_wide[i_word*2+:2]);
  end

  // Propagate integrity error only if wide ISPR is used.

  // Handle ISPR integrity error detection. We've got a bitmask of ISPR words that failed their
  // integrity check (ispr_rdata_intg_err_narrow), but a nonzero entry may not be a problem if we
  // don't actually use the data.
  //
  // The situations when the data is actually used are:
  //
  //   (1) This is a bignum instruction that writes back to the bignum register file by reading an
  //       ISPR. In this case, we actually pass the data through with integrity bits, but it
  //       shouldn't hurt to add fault detection at this point.
  //
  //   (2) This instruction consumes the data by selecting a word from an ISPR and then writing it
  //       back. This happens for things like CSRRS instructions, where the data flows to the base
  //       register file through rf_base_wr_data_no_intg_o and back to the ISPR through
  //       ispr_base_wdata_o. The word used is given by the onehot ispr_word_sel_base mask.
  //
  // In both cases, there's a special case for the RND_PREFETCH register, which doesn't actually
  // have any backing data. It reads as zero with invalid integrity bits which we want to ignore.

  // Are we reading all the ISPR data? (case (1) above)
  logic all_ispr_words_used;
  assign all_ispr_words_used = (insn_dec_bignum_i.rf_wdata_sel == RfWdSelIspr);

  // Are we reading just one word of the ISPR data? (case (2) above).
  logic one_ispr_word_used;
  assign one_ispr_word_used = ispr_rd_insn & (insn_dec_shared_i.subset == InsnSubsetBase);

  // A bit-mask giving which ISPR words are being read
  logic [BaseWordsPerWLEN-1:0] ispr_read_mask;
  assign ispr_read_mask = all_ispr_words_used ? '1 :
                          one_ispr_word_used  ? ispr_word_sel_base : '0;

  // Use ispr_read_mask to qualify the error bit-mask that came out of the integrity decoder.
  logic [BaseWordsPerWLEN-1:0] ispr_rdata_used_intg_err;
  assign ispr_rdata_used_intg_err = ispr_read_mask & ispr_rdata_intg_err_narrow;

  // We only architecturally read the ISPR when there's a non-stalled instruction. This is also the
  // place where we factor in the special RND_PREFETCH behaviour. We also need to squash any
  // integrity errors if we're reading a sideload key which isn't currently valid (this will
  // generate a key_invalid error, but we shouldn't have any behaviour that depends on what happens
  // to be on the pins)
  logic non_prefetch_insn_running;
  assign non_prefetch_insn_running = (insn_valid_i & ~stall &
                                      (csr_addr != CsrRndPrefetch) & ~key_invalid);
  // zdr ecc disable
  // logic ispr_rdata_used_intg_err_zdr = (|ispr_rdata_used_intg_err) & 1'b0;
  assign ispr_rdata_intg_err = non_prefetch_insn_running & |((|ispr_rdata_used_intg_err) & 1'b0);

  `ASSERT_KNOWN(IsprRdataIntgErrKnown_A, ispr_rdata_intg_err)

  for (genvar i_bit = 0; i_bit < 32; i_bit++) begin : g_csr_rdata_mux
    for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_csr_rdata_mux_inner
      assign csr_rdata_mux[i_bit][i_word] =
          ispr_rdata[i_word*32 + i_bit] & ispr_word_sel_base[i_word];
    end

    assign csr_rdata_raw[i_bit] = |csr_rdata_mux[i_bit];
  end

  // Specialised read data handling for CSR reads where raw read data needs modification.
  always_comb begin
    csr_rdata = csr_rdata_raw;

    unique case (csr_addr)
      // For FG0/FG1 select out appropriate bits from FLAGS ISPR and pad the rest with zeros.
      CsrFg0:         csr_rdata = {28'b0, csr_rdata_raw[3:0]};
      CsrFg1:         csr_rdata = {28'b0, csr_rdata_raw[7:4]};
      CsrRndPrefetch: csr_rdata = '0;
      default: ;
    endcase
  end

  assign csr_wdata_raw = insn_dec_shared_i.ispr_rs_insn ? csr_rdata | rf_base_rd_data_a_no_intg :
                                                          rf_base_rd_data_a_no_intg;

  // Specialised write data handling for CSR writes where raw write data needs modification.
  always_comb begin
    csr_wdata = csr_wdata_raw;

    unique case (csr_addr)
      // For FG0/FG1 only modify relevant part of FLAGS ISPR.
      CsrFg0: csr_wdata = {24'b0, csr_rdata_raw[7:4], csr_wdata_raw[3:0]};
      CsrFg1: csr_wdata = {24'b0, csr_wdata_raw[3:0], csr_rdata_raw[3:0]};
      default: ;
    endcase
  end

  // ISPR RS (read and set) must not be combined with ISPR RD or WR (read or write). ISPR RD and
  // WR (read and write) is allowed.
  `ASSERT(NoIsprRorWAndRs, insn_valid_i |-> ~(insn_dec_shared_i.ispr_rs_insn   &
                                              (insn_dec_shared_i.ispr_rd_insn |
                                               insn_dec_shared_i.ispr_wr_insn)))


  assign wsr_addr = wsr_e'(insn_dec_bignum_i.i[WsrNumWidth-1:0]);

  always_comb begin
    ispr_addr_bignum = IsprMod;
    wsr_illegal_addr = 1'b0;
    key_invalid      = 1'b0;

    unique case (wsr_addr)
      WsrMod:  ispr_addr_bignum = IsprMod;
      WsrRnd:  ispr_addr_bignum = IsprRnd;
      WsrUrnd: ispr_addr_bignum = IsprUrnd;
      WsrAcc:  ispr_addr_bignum = IsprAcc;
      WsrKeyS0L: begin
        ispr_addr_bignum = IsprKeyS0L;
        key_invalid = ~sideload_key_shares_valid_i[0];
      end
      WsrKeyS0H: begin
        ispr_addr_bignum = IsprKeyS0H;
        key_invalid = ~sideload_key_shares_valid_i[0];
      end
      WsrKeyS1L: begin
        ispr_addr_bignum = IsprKeyS1L;
        key_invalid = ~sideload_key_shares_valid_i[1];
      end
      WsrKeyS1H: begin
        ispr_addr_bignum = IsprKeyS1H;
        key_invalid = ~sideload_key_shares_valid_i[1];
      end
      default: wsr_illegal_addr = 1'b1;
    endcase
  end

  assign wsr_wdata = insn_dec_shared_i.ispr_rs_insn ? ispr_rdata | rf_bignum_rd_data_a_no_intg :
                                                      rf_bignum_rd_data_a_no_intg;

  assign ispr_illegal_addr = insn_dec_shared_i.subset == InsnSubsetBase ? csr_illegal_addr :
                                                                          wsr_illegal_addr;

  assign ispr_err = ispr_illegal_addr & insn_valid_i & (insn_dec_shared_i.ispr_rd_insn |
                                                        insn_dec_shared_i.ispr_wr_insn |
                                                        insn_dec_shared_i.ispr_rs_insn);

  assign ispr_wr_insn = insn_dec_shared_i.ispr_wr_insn | insn_dec_shared_i.ispr_rs_insn;
  assign ispr_rd_insn = insn_dec_shared_i.ispr_rd_insn | insn_dec_shared_i.ispr_rs_insn;

  assign ispr_flags_wr_o = insn_dec_shared_i.ispr_flags_wr;

  // Write to RND_PREFETCH must not produce ISR write
  assign ispr_wr_base_insn =
    ispr_wr_insn & (insn_dec_shared_i.subset == InsnSubsetBase) & (csr_addr != CsrRndPrefetch);

  assign ispr_wr_bignum_insn = ispr_wr_insn & (insn_dec_shared_i.subset == InsnSubsetBignum);
  assign ispr_rd_bignum_insn = ispr_rd_insn & (insn_dec_shared_i.subset == InsnSubsetBignum);

  assign ispr_addr_o         = insn_dec_shared_i.subset == InsnSubsetBase ? ispr_addr_base :
                                                                            ispr_addr_bignum;
  assign ispr_base_wdata_o   = csr_wdata;
  assign ispr_base_wr_en_o   = {BaseWordsPerWLEN{ispr_wr_base_insn & insn_valid_i}} &
                               ispr_word_sel_base;

  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_ispr_bignum_wdata_enc
    prim_secded_inv_39_32_enc i_secded_enc (
      .data_i(wsr_wdata[i_word*32+:32]),
      .data_o(ispr_bignum_wdata_intg_o[i_word*39+:39])
    );
  end
  assign ispr_bignum_wr_en_o = ispr_wr_bignum_insn & insn_valid_i;

  assign ispr_wr_commit_o = ispr_wr_insn & insn_executing;
  assign ispr_rd_en_o     = ispr_rd_insn & insn_valid_i &
    ~((insn_dec_shared_i.subset == InsnSubsetBase) & (csr_addr == CsrRndPrefetch));

  // For BN.SID the LSU address is computed in the first cycle by the base ALU. The store request
  // itself occurs in the second cycle when the store data is available (from the indirect register
  // read). The calculated address is saved in a flop here so it's available for use in the second
  // cycle.
  assign lsu_addr_saved_d = alu_base_operation_result_i[DmemAddrWidth-1:0];
  always_ff @(posedge clk_i) begin
    lsu_addr_saved_q <= lsu_addr_saved_d;
  end

  //assign expected_lsu_addr_en_predec = insn_valid & insn_dec_shared_i.ld_insn

  // lsu_load_req_raw/lsu_store_req_raw indicate an instruction wishes to perform a store or a load.
  // lsu_load_req_o/lsu_store_req_o factor in whether an instruction is actually executing (it may
  // be suppressed due an error) and command the load or store to happen when asserted.
  assign lsu_load_req_raw = insn_valid_i & insn_dec_shared_i.ld_insn & (state_q == OtbnStateRun);
  assign lsu_load_req_o   = insn_executing & lsu_load_req_raw;

  assign lsu_store_req_raw = insn_valid_i & insn_dec_shared_i.st_insn & ~rf_indirect_stall;
  assign lsu_store_req_o   = insn_executing & lsu_store_req_raw;

  assign lsu_req_subset_o = insn_dec_shared_i.subset;

  // To simplify blanking logic all two cycle memory operations (BN.LID, BN.SID, LW) present the
  // calculated address in their first cycle and the saved address in the second cycle. This results
  // in lsu_addr_o remaining stable for the entire instruction. Only SW is a single cycle
  // instruction so it only presents the calculated address. The stability property is checked by an
  // assertion.
  assign lsu_addr_saved_sel =
    insn_valid_i & ((insn_dec_shared_i.subset == InsnSubsetBignum) ||
                    insn_dec_shared_i.ld_insn                         ? ~stall : 1'b0);

  assign lsu_addr = lsu_addr_saved_sel ? lsu_addr_saved_q                                :
                                         alu_base_operation_result_i[DmemAddrWidth-1:0];

  // SEC_CM: CTRL.REDUN
  assign expected_lsu_addr_en =
    insn_valid_i & (insn_dec_shared_i.ld_insn | insn_dec_shared_i.st_insn);

  assign lsu_predec_error = expected_lsu_addr_en != lsu_addr_en_predec_i;

  assign expected_call_stack_push =
    insn_valid_i & insn_dec_base_i.rf_we & rf_base_wr_addr_o == 5'd1;

  assign expected_call_stack_pop = insn_valid_i &
                                   ((insn_dec_base_i.rf_ren_a & rf_base_rd_addr_a_o == 5'd1) |
                                    (insn_dec_base_i.rf_ren_b & rf_base_rd_addr_b_o == 5'd1));

  // Check branch target against the precalculated target from pre-decode. Pre-decode cannot
  // calculate the jump target of a JALR as it requires a register read so this is excluded from the
  // check (by looking at the ALU op a selection).
  assign branch_target_predec_error =
    insn_dec_shared_i.branch_insn                                            &
    insn_dec_shared_i.jump_insn & insn_dec_base_i.op_a_sel != OpASelRegister &
    (ctrl_flow_target_predec_i != branch_target);

  assign ctrl_predec_error =
    |{ctrl_flow_predec_i.jump_insn       != (insn_dec_shared_i.jump_insn   & insn_valid_i),
      ctrl_flow_predec_i.loop_insn       != (insn_dec_shared_i.loop_insn   & insn_valid_i),
      ctrl_flow_predec_i.branch_insn     != (insn_dec_shared_i.branch_insn & insn_valid_i),
      ctrl_flow_predec_i.sel_insn        != (insn_dec_bignum_i.sel_insn    & insn_valid_i),
      ctrl_flow_predec_i.call_stack_push != expected_call_stack_push,
      ctrl_flow_predec_i.call_stack_pop  != expected_call_stack_pop,
      branch_target_predec_error,
      loop_predec_err};

  assign predec_error_o = lsu_predec_error | ctrl_predec_error;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(DmemAddrWidth)) u_lsu_addr_blanker (
    .in_i (lsu_addr),
    .en_i (lsu_addr_en_predec_i),
    .out_o(lsu_addr_blanked)
  );

  // Check stability property described above (see the lsu_addr_saved_sel signal) holds.
  `ASSERT(LsuAddrBlankedStable_A, insn_valid_i & stall & ~err |=> $stable(lsu_addr_blanked))

  assign lsu_addr_o = lsu_addr_blanked;

  assign lsu_base_wdata_o   = rf_base_rd_data_b_intg_i;
  assign lsu_bignum_wdata_o = rf_bignum_rd_data_b_intg_i;

  assign dmem_addr_unaligned_bignum =
      (lsu_req_subset_o == InsnSubsetBignum) & (|lsu_addr_o[$clog2(WLEN/8)-1:0]);
  assign dmem_addr_unaligned_base   =
      (lsu_req_subset_o == InsnSubsetBase)   & (|lsu_addr_o[1:0]);
  assign dmem_addr_overflow         = |alu_base_operation_result_i[31:DmemAddrWidth];

  // A dmem address is checked the cycle it is available. For bignum stores this is the first cycle
  // where the base register file read occurs, with the store request occurring the following cycle.
  // For all other loads and stores the dmem address is available the same cycle as the request.
  assign dmem_addr_err_check =
    (lsu_req_subset_o == InsnSubsetBignum) &
    insn_dec_shared_i.st_insn               ? rf_indirect_stall :
                                              lsu_load_req_raw | lsu_store_req_raw;

  assign dmem_addr_err =
      insn_valid_i & dmem_addr_err_check & (dmem_addr_overflow         |
                                            dmem_addr_unaligned_bignum |
                                            dmem_addr_unaligned_base);

  assign rnd_req_raw = insn_valid_i & ispr_rd_insn & (ispr_addr_o == IsprRnd);
  // Don't factor rnd_rep/fips_err_i into rnd_req_o. This would lead to a combo loop.
  assign rnd_req_o = rnd_req_raw & insn_valid_i & ~(software_err | fatal_err);

  assign rnd_prefetch_req_o = insn_executing & ispr_wr_insn &
      (insn_dec_shared_i.subset == InsnSubsetBase) & (csr_addr == CsrRndPrefetch);
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN instruction Decoder
 */
module otbn_decoder
  import otbn_pkg::*;
(
  // For assertions only.
  input logic clk_i,
  input logic rst_ni,

  // instruction data to be decoded
  input logic [31:0] insn_fetch_resp_data_i,
  input logic        insn_fetch_resp_valid_i,

  // Decoded instruction
  output logic insn_valid_o,
  output logic insn_illegal_o,

  output insn_dec_base_t   insn_dec_base_o,
  output insn_dec_bignum_t insn_dec_bignum_o,
  output insn_dec_shared_t insn_dec_shared_o
);

  logic        illegal_insn;
  logic        rf_we_base;
  logic        rf_we_bignum;

  logic [31:0] insn;
  logic [31:0] insn_alu;

  // Source/Destination register instruction index
  logic [4:0] insn_rs1;
  logic [4:0] insn_rs2;
  logic [4:0] insn_rd;

  insn_opcode_e     opcode;
  insn_opcode_e     opcode_alu;

  assign insn     = insn_fetch_resp_data_i;
  assign insn_alu = insn_fetch_resp_data_i;

  logic unused_insn_alu_bits;
  assign unused_insn_alu_bits = (|insn_alu[11:7]) | (|insn_alu[24:15]);

  //////////////////////////////////////
  // Register and immediate selection //
  //////////////////////////////////////
  imm_b_sel_base_e   imm_b_mux_sel_base; // immediate selection for operand b in base ISA
  shamt_sel_bignum_e shift_amt_mux_sel_bignum; // shift amount selection in bignum ISA

  // Immediates from RV32I encoding
  logic [31:0] imm_i_type_base;
  logic [31:0] imm_s_type_base;
  logic [31:0] imm_b_type_base;
  logic [31:0] imm_u_type_base;
  logic [31:0] imm_j_type_base;

  // Immediates specific to OTBN encoding
  logic [31:0] imm_l_type_base;
  logic [31:0] imm_x_type_base;

  alu_op_base_e   alu_operator_base;      // ALU operation selection for base ISA
  alu_op_bignum_e alu_operator_bignum;    // ALU operation selection for bignum ISA

  op_a_sel_e alu_op_a_mux_sel_base; // operand a selection for base ISA: reg value, PC or zero
  op_b_sel_e alu_op_b_mux_sel_base; // operand b selection for base ISA: reg value or immediate

  op_b_sel_e alu_op_b_mux_sel_bignum; // operand b selection for bignum ISA: reg value or immediate

  comparison_op_base_e comparison_operator_base;


  logic [1:0] mac_op_a_qw_sel_bignum;
  logic [1:0] mac_op_b_qw_sel_bignum;
  logic       mac_wr_hw_sel_upper_bignum;
  logic [1:0] mac_pre_acc_shift_bignum;
  logic       mac_zero_acc_bignum;
  logic       mac_shift_out_bignum;
  logic       mac_en_bignum;

  logic rf_ren_a_base;
  logic rf_ren_b_base;

  logic rf_ren_a_bignum;
  logic rf_ren_b_bignum;

  logic rf_a_indirect_bignum;
  logic rf_b_indirect_bignum;
  logic rf_d_indirect_bignum;

  // immediate extraction and sign extension
  assign imm_i_type_base = {{20{insn[31]}}, insn[31:20]};
  assign imm_s_type_base = {{20{insn[31]}}, insn[31:25], insn[11:7]};
  assign imm_b_type_base = {{19{insn[31]}}, insn[31], insn[7], insn[30:25], insn[11:8], 1'b0};
  assign imm_u_type_base = {insn[31:12], 12'b0};
  assign imm_j_type_base = {{12{insn[31]}}, insn[19:12], insn[20], insn[30:21], 1'b0};
  // l type immediate is for the loop count in the LOOPI instruction and is not from the RISC-V ISA
  assign imm_l_type_base = {22'b0, insn[19:15], insn[11:7]};
  // x type immediate is for BN.LID/BN.SID instructions and is not from the RISC-V ISA
  assign imm_x_type_base = {{17{insn[11]}}, insn[11:9], insn[31:25], 5'b0};

  logic [WLEN-1:0] imm_i_type_bignum;

  assign imm_i_type_bignum = {{(WLEN-10){1'b0}}, insn[29:20]};

  // Shift amount for ALU instructions other than BN.RSHI
  logic [$clog2(WLEN)-1:0] shift_amt_a_type_bignum;
  // Shift amount for BN.RSHI
  logic [$clog2(WLEN)-1:0] shift_amt_s_type_bignum;

  assign shift_amt_a_type_bignum = {insn[29:25], 3'b0};
  assign shift_amt_s_type_bignum = {insn[31:25], insn[14]};

  logic alu_shift_right_bignum;

  assign alu_shift_right_bignum = insn[30];

  flag_group_t alu_flag_group_bignum;

  assign alu_flag_group_bignum = insn[31];

  flag_e alu_sel_flag_bignum;

  assign alu_sel_flag_bignum = flag_e'(insn[26:25]);

  logic alu_flag_en_bignum;
  logic mac_flag_en_bignum;

  // source registers
  assign insn_rs1 = insn[19:15];
  assign insn_rs2 = insn[24:20];

  // destination register
  assign insn_rd = insn[11:7];

  insn_subset_e insn_subset;
  rf_wd_sel_e rf_wdata_sel_base;
  rf_wd_sel_e rf_wdata_sel_bignum;

  logic [11:0] loop_bodysize_base;
  logic        loop_immediate_base;

  assign loop_bodysize_base  = insn[31:20];
  assign loop_immediate_base = insn[12];

  assign mac_op_a_qw_sel_bignum     = insn[26:25];
  assign mac_op_b_qw_sel_bignum     = insn[28:27];
  assign mac_wr_hw_sel_upper_bignum = insn[29];
  assign mac_pre_acc_shift_bignum   = insn[14:13];
  assign mac_zero_acc_bignum        = insn[12];
  assign mac_shift_out_bignum       = insn[30];

  logic d_inc_bignum;
  logic a_inc_bignum;
  logic a_wlen_word_inc_bignum;
  logic b_inc_bignum;

  logic sel_insn_bignum;

  logic ecall_insn;
  logic ld_insn;
  logic st_insn;
  logic branch_insn;
  logic jump_insn;
  logic loop_insn;
  logic ispr_rd_insn;
  logic ispr_wr_insn;
  logic ispr_rs_insn;
  logic [NFlagGroups-1:0] ispr_flags_wr;

  // Reduced main ALU immediate MUX for Operand B
  logic [31:0] imm_b_base;
  always_comb begin : immediate_b_mux
    unique case (imm_b_mux_sel_base)
      ImmBaseBI: imm_b_base = imm_i_type_base;
      ImmBaseBS: imm_b_base = imm_s_type_base;
      ImmBaseBU: imm_b_base = imm_u_type_base;
      ImmBaseBB: imm_b_base = imm_b_type_base;
      ImmBaseBJ: imm_b_base = imm_j_type_base;
      ImmBaseBL: imm_b_base = imm_l_type_base;
      ImmBaseBX: imm_b_base = imm_x_type_base;
      default:   imm_b_base = imm_i_type_base;
    endcase
  end

  logic [$clog2(WLEN)-1:0] alu_shift_amt_bignum;
  always_comb begin
    unique case (shift_amt_mux_sel_bignum)
      ShamtSelBignumA:    alu_shift_amt_bignum = shift_amt_a_type_bignum;
      ShamtSelBignumS:    alu_shift_amt_bignum = shift_amt_s_type_bignum;
      ShamtSelBignumZero: alu_shift_amt_bignum = '0;
      default:            alu_shift_amt_bignum = shift_amt_a_type_bignum;
    endcase
  end

  assign insn_valid_o   = insn_fetch_resp_valid_i & ~illegal_insn;
  assign insn_illegal_o = insn_fetch_resp_valid_i & illegal_insn;

  assign insn_dec_base_o = '{
    a:              insn_rs1,
    b:              insn_rs2,
    d:              insn_rd,
    i:              imm_b_base,
    alu_op:         alu_operator_base,
    comparison_op:  comparison_operator_base,
    op_a_sel:       alu_op_a_mux_sel_base,
    op_b_sel:       alu_op_b_mux_sel_base,
    rf_we:          rf_we_base,
    rf_wdata_sel:   rf_wdata_sel_base,
    rf_ren_a:       rf_ren_a_base,
    rf_ren_b:       rf_ren_b_base,
    loop_bodysize:  loop_bodysize_base,
    loop_immediate: loop_immediate_base
  };

  assign insn_dec_bignum_o = '{
    a:                   insn_rs1,
    b:                   insn_rs2,
    d:                   insn_rd,
    i:                   imm_i_type_bignum,
    rf_a_indirect:       rf_a_indirect_bignum,
    rf_b_indirect:       rf_b_indirect_bignum,
    rf_d_indirect:       rf_d_indirect_bignum,
    d_inc:               d_inc_bignum,
    a_inc:               a_inc_bignum,
    a_wlen_word_inc:     a_wlen_word_inc_bignum,
    b_inc:               b_inc_bignum,
    alu_shift_amt:       alu_shift_amt_bignum,
    alu_shift_right:     alu_shift_right_bignum,
    alu_flag_group:      alu_flag_group_bignum,
    alu_sel_flag:        alu_sel_flag_bignum,
    alu_flag_en:         alu_flag_en_bignum,
    mac_flag_en:         mac_flag_en_bignum,
    alu_op:              alu_operator_bignum,
    alu_op_b_sel:        alu_op_b_mux_sel_bignum,
    mac_op_a_qw_sel:     mac_op_a_qw_sel_bignum,
    mac_op_b_qw_sel:     mac_op_b_qw_sel_bignum,
    mac_wr_hw_sel_upper: mac_wr_hw_sel_upper_bignum,
    mac_pre_acc_shift:   mac_pre_acc_shift_bignum,
    mac_zero_acc:        mac_zero_acc_bignum,
    mac_shift_out:       mac_shift_out_bignum,
    mac_en:              mac_en_bignum,
    rf_we:               rf_we_bignum,
    rf_wdata_sel:        rf_wdata_sel_bignum,
    rf_ren_a:            rf_ren_a_bignum,
    rf_ren_b:            rf_ren_b_bignum,
    sel_insn:            sel_insn_bignum
  };

  assign insn_dec_shared_o = '{
    subset:        insn_subset,
    ecall_insn:    ecall_insn,
    ld_insn:       ld_insn,
    st_insn:       st_insn,
    branch_insn:   branch_insn,
    jump_insn:     jump_insn,
    loop_insn:     loop_insn,
    ispr_rd_insn:  ispr_rd_insn,
    ispr_wr_insn:  ispr_wr_insn,
    ispr_rs_insn:  ispr_rs_insn,
    ispr_flags_wr: ispr_flags_wr
  };

  /////////////
  // Decoder //
  /////////////

  always_comb begin
    insn_subset            = InsnSubsetBase;

    rf_wdata_sel_base      = RfWdSelEx;
    rf_we_base             = 1'b0;

    rf_wdata_sel_bignum    = RfWdSelEx;
    rf_we_bignum           = 1'b0;

    rf_ren_a_base          = 1'b0;
    rf_ren_b_base          = 1'b0;
    rf_ren_a_bignum        = 1'b0;
    rf_ren_b_bignum        = 1'b0;
    mac_en_bignum          = 1'b0;

    rf_a_indirect_bignum   = 1'b0;
    rf_b_indirect_bignum   = 1'b0;
    rf_d_indirect_bignum   = 1'b0;

    d_inc_bignum           = 1'b0;
    a_inc_bignum           = 1'b0;
    a_wlen_word_inc_bignum = 1'b0;
    b_inc_bignum           = 1'b0;

    illegal_insn           = 1'b0;
    ecall_insn             = 1'b0;
    ld_insn                = 1'b0;
    st_insn                = 1'b0;
    branch_insn            = 1'b0;
    jump_insn              = 1'b0;
    loop_insn              = 1'b0;
    ispr_rd_insn           = 1'b0;
    ispr_wr_insn           = 1'b0;
    ispr_rs_insn           = 1'b0;
    ispr_flags_wr          = '0;

    sel_insn_bignum        = 1'b0;

    opcode                 = insn_opcode_e'(insn[6:0]);

    unique case (opcode)
      //////////////
      // Base ALU //
      //////////////

      InsnOpcodeBaseLui: begin  // Load Upper Immediate
        insn_subset = InsnSubsetBase;
        rf_we_base  = 1'b1;
      end

      InsnOpcodeBaseOpImm: begin  // Register-Immediate ALU Operations
        insn_subset   = InsnSubsetBase;
        rf_ren_a_base = 1'b1;
        rf_we_base    = 1'b1;

        unique case (insn[14:12])
          3'b000,  // addi
          3'b100,  // xori
          3'b110,  // ori
          3'b111:  // andi
            illegal_insn = 1'b0;

          3'b001: begin
            unique case (insn[31:25])
              7'b0000000: illegal_insn = 1'b0;  // slli
              default: illegal_insn = 1'b1;
            endcase
          end

          3'b101: begin
            unique case (insn[31:25])
              7'b0000000,                      // srli
              7'b0100000: illegal_insn = 1'b0; // srai

              default: illegal_insn = 1'b1;
            endcase
          end

          default: illegal_insn = 1'b1;
        endcase
      end

      InsnOpcodeBaseOp: begin  // Register-Register ALU operation
        insn_subset   = InsnSubsetBase;
        rf_ren_a_base = 1'b1;
        rf_ren_b_base = 1'b1;
        rf_we_base    = 1'b1;
        // Look at the funct7 and funct3 fields.
        unique case ({insn[31:25], insn[14:12]})
          {7'b000_0000, 3'b000},  // ADD
          {7'b010_0000, 3'b000},  // SUB
          {7'b000_0000, 3'b100},  // XOR
          {7'b000_0000, 3'b110},  // OR
          {7'b000_0000, 3'b111},  // AND
          {7'b000_0000, 3'b001},  // SLL
          {7'b000_0000, 3'b101},  // SRL
          {7'b010_0000, 3'b101}:  // SRA
            illegal_insn = 1'b0;

          default: begin
            illegal_insn = 1'b1;
          end
        endcase
      end

      ///////////////////////
      // Base Loads/Stores //
      ///////////////////////

      InsnOpcodeBaseLoad: begin
        insn_subset       = InsnSubsetBase;
        ld_insn           = 1'b1;
        rf_ren_a_base     = 1'b1;
        rf_we_base        = 1'b1;
        rf_wdata_sel_base = RfWdSelLsu;

        if (insn[14:12] != 3'b010) begin
          illegal_insn = 1'b1;
        end
      end

      InsnOpcodeBaseStore: begin
        insn_subset   = InsnSubsetBase;
        st_insn       = 1'b1;
        rf_ren_a_base = 1'b1;
        rf_ren_b_base = 1'b1;

        if (insn[14:12] != 3'b010) begin
          illegal_insn = 1'b1;
        end
      end

      //////////////////////
      // Base Branch/Jump //
      //////////////////////

      InsnOpcodeBaseBranch: begin
        insn_subset   = InsnSubsetBase;
        branch_insn   = 1'b1;
        rf_ren_a_base = 1'b1;
        rf_ren_b_base = 1'b1;

        // Only EQ & NE comparisons allowed
        if (insn[14:13] != 2'b00) begin
          illegal_insn = 1'b1;
        end
      end

      InsnOpcodeBaseJal: begin
        insn_subset       = InsnSubsetBase;
        jump_insn         = 1'b1;
        rf_we_base        = 1'b1;
        rf_wdata_sel_base = RfWdSelNextPc;
      end

      InsnOpcodeBaseJalr: begin
        insn_subset       = InsnSubsetBase;
        jump_insn         = 1'b1;
        rf_ren_a_base     = 1'b1;
        rf_we_base        = 1'b1;
        rf_wdata_sel_base = RfWdSelNextPc;

        if (insn[14:12] != 3'b000) begin
          illegal_insn = 1'b1;
        end
      end

      //////////////////
      // Base Special //
      //////////////////

      InsnOpcodeBaseSystem: begin
        insn_subset = InsnSubsetBase;
        if (insn[14:12] == 3'b000) begin
          // non CSR related SYSTEM instructions
          unique case (insn[31:20])
            12'h000:  // ECALL
              ecall_insn = 1'b1;

            default:
              illegal_insn = 1'b1;
          endcase

          // rs1 and rd must be 0
          if (insn_rs1 != 5'b0 || insn_rd != 5'b0) begin
            illegal_insn = 1'b1;
          end
        end else begin
          rf_we_base        = 1'b1;
          rf_wdata_sel_base = RfWdSelIspr;
          rf_ren_a_base     = 1'b1;

          if (insn[14:12] == 3'b001) begin
            // No read if destination is x0 unless read is to flags CSR. Both flag groups are in
            // a single ISPR so to write one group the other must be read to write it back
            // unchanged.
            ispr_rd_insn  = (insn_rd != 5'b0)            |
                            (imm_b_base[11:0] == CsrFg0) |
                            (imm_b_base[11:0] == CsrFg1);
            ispr_wr_insn  = 1'b1;
            ispr_flags_wr = {(imm_b_base[11:0] == CsrFg1), (imm_b_base[11:0] == CsrFg0)} |
                            {NFlagGroups{imm_b_base[11:0] == CsrFlags}};
          end else if (insn[14:12] == 3'b010) begin
            // Read and set if source register isn't x0, otherwise read only
            if (insn_rs1 != 5'b0) begin
              ispr_rs_insn  = 1'b1;
              ispr_flags_wr = {(imm_b_base[11:0] == CsrFg1), (imm_b_base[11:0] == CsrFg0)} |
                              {NFlagGroups{imm_b_base[11:0] == CsrFlags}};
            end else begin
              ispr_rd_insn = 1'b1;
            end
          end else begin
            illegal_insn = 1'b1;
          end
        end
      end

      ////////////////
      // Bignum ALU //
      ////////////////

      InsnOpcodeBignumArith: begin
        insn_subset     = InsnSubsetBignum;
        rf_we_bignum    = 1'b1;
        rf_ren_a_bignum = 1'b1;

        if (insn[14:12] != 3'b100) begin
          // All Alu instructions other than BN.ADDI/BN.SUBI
          rf_ren_b_bignum = 1'b1;
        end

        unique case(insn[14:12])
          3'b110,
          3'b111: illegal_insn = 1'b1;
          default: ;
        endcase
      end

      ///////////////////////////////////////
      // Bignum logical/BN.RSHI/LOOP/LOOPI //
      ///////////////////////////////////////

      InsnOpcodeBignumBaseMisc: begin
        unique case (insn[14:12])
          3'b000, 3'b001: begin  // LOOP[I]
            insn_subset   = InsnSubsetBase;
            rf_ren_a_base = ~insn[12];
            loop_insn     = 1'b1;
          end
          3'b010, 3'b011, 3'b100, 3'b110, 3'b111: begin  // BN.RHSI/BN.AND/BN.OR/BN.XOR
            insn_subset     = InsnSubsetBignum;
            rf_we_bignum    = 1'b1;
            rf_ren_a_bignum = 1'b1;
            rf_ren_b_bignum = 1'b1;
          end
          3'b101: begin  // BN.NOT
            insn_subset     = InsnSubsetBignum;
            rf_we_bignum    = 1'b1;
            rf_ren_b_bignum = 1'b1;
          end
          default: illegal_insn = 1'b1;
        endcase
      end

      ///////////////////////////////////////////////
      // Bignum Misc WSR/LID/SID/MOV[R]/CMP[B]/SEL //
      ///////////////////////////////////////////////

      InsnOpcodeBignumMisc: begin
        insn_subset = InsnSubsetBignum;

        unique case (insn[14:12])
          3'b000: begin  // BN.SEL
            rf_we_bignum        = 1'b1;
            rf_ren_a_bignum     = 1'b1;
            rf_ren_b_bignum     = 1'b1;
            rf_wdata_sel_bignum = RfWdSelMovSel;
            sel_insn_bignum     = 1'b1;
          end
          3'b011, 3'b001: begin  // BN.CMP[B]
            rf_ren_a_bignum = 1'b1;
            rf_ren_b_bignum = 1'b1;
          end
          3'b100: begin  // BN.LID
            ld_insn              = 1'b1;
            rf_we_bignum         = 1'b1;
            rf_ren_a_base        = 1'b1;
            rf_ren_b_base        = 1'b1;
            rf_wdata_sel_bignum  = RfWdSelLsu;
            rf_d_indirect_bignum = 1'b1;

            if (insn[8]) begin
              a_wlen_word_inc_bignum = 1'b1;
              rf_we_base             = 1'b1;
              rf_wdata_sel_base      = RfWdSelIncr;
            end

            if (insn[7]) begin
              d_inc_bignum      = 1'b1;
              rf_we_base        = 1'b1;
              rf_wdata_sel_base = RfWdSelIncr;
            end

            if (insn[8] & insn[7]) begin
              // Avoid violating unique constraint for inc selection mux on an illegal instruction
              a_wlen_word_inc_bignum = 1'b0;
              d_inc_bignum           = 1'b0;
              illegal_insn           = 1'b1;
            end
          end
          3'b101: begin  // BN.SID
            st_insn              = 1'b1;
            rf_ren_a_base        = 1'b1;
            rf_ren_b_base        = 1'b1;
            rf_ren_b_bignum      = 1'b1;
            rf_b_indirect_bignum = 1'b1;

            if (insn[8]) begin
              a_wlen_word_inc_bignum = 1'b1;
              rf_we_base             = 1'b1;
              rf_wdata_sel_base      = RfWdSelIncr;
            end

            if (insn[7]) begin
              b_inc_bignum = 1'b1;
              rf_we_base   = 1'b1;
              rf_wdata_sel_base = RfWdSelIncr;
            end

            if (insn[8] & insn[7]) begin
              // Avoid violating unique constraint for inc selection mux on an illegal instruction
              a_wlen_word_inc_bignum = 1'b0;
              b_inc_bignum           = 1'b0;
              illegal_insn           = 1'b1;
            end
          end
          3'b110: begin  // BN.MOV/BN.MOVR
            insn_subset         = InsnSubsetBignum;
            rf_we_bignum        = 1'b1;
            rf_ren_a_bignum     = 1'b1;
            rf_wdata_sel_bignum = RfWdSelMovSel;

            if (insn[31]) begin  // BN.MOVR
              rf_a_indirect_bignum = 1'b1;
              rf_d_indirect_bignum = 1'b1;
              rf_ren_a_base        = 1'b1;
              rf_ren_b_base        = 1'b1;

              if (insn[9]) begin
                a_inc_bignum      = 1'b1;
                rf_we_base        = 1'b1;
                rf_wdata_sel_base = RfWdSelIncr;
              end

              if (insn[7]) begin
                d_inc_bignum      = 1'b1;
                rf_we_base        = 1'b1;
                rf_wdata_sel_base = RfWdSelIncr;
              end

              if (insn[9] & insn[7]) begin
                // Avoid violating unique constraint for inc selection mux on an illegal instruction
                a_inc_bignum = 1'b0;
                d_inc_bignum = 1'b0;
                illegal_insn = 1'b1;
              end
            end
          end
          3'b111: begin
            if (insn[31]) begin  // BN.WSRW
              rf_ren_a_bignum = 1'b1;
              ispr_wr_insn    = 1'b1;
            end else begin  // BN.WSRR
              rf_we_bignum        = 1'b1;
              rf_wdata_sel_bignum = RfWdSelIspr;
              ispr_rd_insn        = 1'b1;
            end
          end
          default: illegal_insn = 1'b1;
        endcase
      end

      ////////////////////////////////////////////
      // BN.MULQACC/BN.MULQACC.WO/BN.MULQACC.SO //
      ////////////////////////////////////////////

      InsnOpcodeBignumMulqacc: begin
        insn_subset         = InsnSubsetBignum;
        rf_ren_a_bignum     = 1'b1;
        rf_ren_b_bignum     = 1'b1;
        rf_wdata_sel_bignum = RfWdSelMac;
        mac_en_bignum       = 1'b1;

        if (insn[30] == 1'b1 || insn[29] == 1'b1) begin  // BN.MULQACC.WO/BN.MULQACC.SO
          rf_we_bignum = 1'b1;
        end
      end

      default: illegal_insn = 1'b1;
    endcase


    // make sure illegal instructions detected in the decoder do not propagate from decoder
    // NOTE: instructions can also be detected to be illegal inside the CSRs (upon accesses with
    // insufficient privileges). These cases are not handled here.
    if (illegal_insn) begin
      rf_we_base   = 1'b0;
      rf_we_bignum = 1'b0;
    end
  end

  /////////////////////////////
  // Decoder for ALU control //
  /////////////////////////////

  always_comb begin
    alu_operator_base        = AluOpBaseAdd;
    comparison_operator_base = ComparisonOpBaseEq;

    alu_op_a_mux_sel_base    = OpASelRegister;
    alu_op_b_mux_sel_base    = OpBSelImmediate;

    imm_b_mux_sel_base       = ImmBaseBI;

    alu_operator_bignum      = AluOpBignumNone;
    alu_op_b_mux_sel_bignum  = OpBSelImmediate;

    shift_amt_mux_sel_bignum = ShamtSelBignumA;

    opcode_alu               = insn_opcode_e'(insn_alu[6:0]);

    alu_flag_en_bignum       = 1'b0;
    mac_flag_en_bignum       = 1'b0;

    unique case (opcode_alu)
      //////////////
      // Base ALU //
      //////////////

      InsnOpcodeBaseLui: begin  // Load Upper Immediate
        alu_op_a_mux_sel_base = OpASelZero;
        alu_op_b_mux_sel_base = OpBSelImmediate;
        imm_b_mux_sel_base    = ImmBaseBU;
        alu_operator_base     = AluOpBaseAdd;
      end

      InsnOpcodeBaseOpImm: begin  // Register-Immediate ALU Operations
        alu_op_a_mux_sel_base = OpASelRegister;
        alu_op_b_mux_sel_base = OpBSelImmediate;
        imm_b_mux_sel_base    = ImmBaseBI;

        unique case (insn_alu[14:12])
          3'b000: alu_operator_base = AluOpBaseAdd;  // Add Immediate
          3'b100: alu_operator_base = AluOpBaseXor;  // Exclusive Or with Immediate
          3'b110: alu_operator_base = AluOpBaseOr;   // Or with Immediate
          3'b111: alu_operator_base = AluOpBaseAnd;  // And with Immediate

          3'b001: begin
            alu_operator_base = AluOpBaseSll;  // Shift Left Logical by Immediate
          end

          3'b101: begin
            if (insn_alu[31:27] == 5'b0_0000) begin
              alu_operator_base = AluOpBaseSrl;  // Shift Right Logical by Immediate
            end else if (insn_alu[31:27] == 5'b0_1000) begin
              alu_operator_base = AluOpBaseSra;  // Shift Right Arithmetically by Immediate
            end
          end

          default: ;
        endcase
      end

      InsnOpcodeBaseOp: begin  // Register-Register ALU operation
        alu_op_a_mux_sel_base = OpASelRegister;
        alu_op_b_mux_sel_base = OpBSelRegister;

        if (!insn_alu[26]) begin
          unique case ({insn_alu[31:25], insn_alu[14:12]})
            // RV32I ALU operations
            {7'b000_0000, 3'b000}: alu_operator_base = AluOpBaseAdd;   // Add
            {7'b010_0000, 3'b000}: alu_operator_base = AluOpBaseSub;   // Sub
            {7'b000_0000, 3'b100}: alu_operator_base = AluOpBaseXor;   // Xor
            {7'b000_0000, 3'b110}: alu_operator_base = AluOpBaseOr;    // Or
            {7'b000_0000, 3'b111}: alu_operator_base = AluOpBaseAnd;   // And
            {7'b000_0000, 3'b001}: alu_operator_base = AluOpBaseSll;   // Shift Left Logical
            {7'b000_0000, 3'b101}: alu_operator_base = AluOpBaseSrl;   // Shift Right Logical
            {7'b010_0000, 3'b101}: alu_operator_base = AluOpBaseSra;   // Shift Right Arithmetic
            default: ;
          endcase
        end
      end

      ///////////////////////
      // Base Loads/Stores //
      ///////////////////////

      InsnOpcodeBaseLoad: begin
        alu_op_a_mux_sel_base = OpASelRegister;
        alu_op_b_mux_sel_base = OpBSelImmediate;
        alu_operator_base     = AluOpBaseAdd;
        imm_b_mux_sel_base    = ImmBaseBI;
      end

      InsnOpcodeBaseStore: begin
        alu_op_a_mux_sel_base = OpASelRegister;
        alu_op_b_mux_sel_base = OpBSelImmediate;
        alu_operator_base     = AluOpBaseAdd;
        imm_b_mux_sel_base    = ImmBaseBS;
      end

      //////////////////////
      // Base Branch/Jump //
      //////////////////////

      InsnOpcodeBaseBranch: begin
        alu_op_a_mux_sel_base    = OpASelCurrPc;
        alu_op_b_mux_sel_base    = OpBSelImmediate;
        alu_operator_base        = AluOpBaseAdd;
        imm_b_mux_sel_base       = ImmBaseBB;
        comparison_operator_base = insn_alu[12] ? ComparisonOpBaseNeq : ComparisonOpBaseEq;
      end

      InsnOpcodeBaseJal: begin
        alu_op_a_mux_sel_base = OpASelCurrPc;
        alu_op_b_mux_sel_base = OpBSelImmediate;
        alu_operator_base     = AluOpBaseAdd;
        imm_b_mux_sel_base    = ImmBaseBJ;
      end

      InsnOpcodeBaseJalr: begin
        alu_op_a_mux_sel_base = OpASelRegister;
        alu_op_b_mux_sel_base = OpBSelImmediate;
        alu_operator_base     = AluOpBaseAdd;
        imm_b_mux_sel_base    = ImmBaseBI;
      end

      //////////////////
      // Base Special //
      //////////////////

      InsnOpcodeBaseSystem: begin
        // The only instructions with System opcode that care about operands are CSR access
        alu_op_a_mux_sel_base = OpASelRegister;
        imm_b_mux_sel_base    = ImmBaseBI;
      end

      ////////////////
      // Bignum ALU //
      ////////////////

      InsnOpcodeBignumArith: begin
        alu_flag_en_bignum = 1'b1;

        unique case (insn_alu[14:12])
          3'b000: alu_operator_bignum = AluOpBignumAdd;
          3'b001: alu_operator_bignum = AluOpBignumSub;
          3'b010: alu_operator_bignum = AluOpBignumAddc;
          3'b011: alu_operator_bignum = AluOpBignumSubb;
          3'b100: begin
            if (insn_alu[30]) begin
              alu_operator_bignum = AluOpBignumSub;
            end else begin
              alu_operator_bignum = AluOpBignumAdd;
            end
          end
          3'b101: begin
            if (insn_alu[30]) begin
              alu_operator_bignum = AluOpBignumSubm;
            end else begin
              alu_operator_bignum = AluOpBignumAddm;
            end
          end
          default: ;
        endcase

        if (insn_alu[14:12] != 3'b100) begin
          alu_op_b_mux_sel_bignum  = OpBSelRegister;
          shift_amt_mux_sel_bignum = ShamtSelBignumA;
        end else begin
          alu_op_b_mux_sel_bignum  = OpBSelImmediate;
          shift_amt_mux_sel_bignum = ShamtSelBignumZero;
        end
      end

      ///////////////////////////////////////
      // Bignum logical/BN.RSHI/LOOP/LOOPI //
      ///////////////////////////////////////

      InsnOpcodeBignumBaseMisc: begin
        // LOOPI uses L type immediate, base immediate irrelevant for everything else
        imm_b_mux_sel_base      = ImmBaseBL;
        alu_op_b_mux_sel_bignum = OpBSelRegister;

        unique case (insn_alu[14:12])
          3'b010: begin
            shift_amt_mux_sel_bignum = ShamtSelBignumA;
            alu_operator_bignum      = AluOpBignumAnd;
            alu_flag_en_bignum       = 1'b1;
          end
          3'b100: begin
            shift_amt_mux_sel_bignum = ShamtSelBignumA;
            alu_operator_bignum      = AluOpBignumOr;
            alu_flag_en_bignum       = 1'b1;
          end
          3'b101: begin
            shift_amt_mux_sel_bignum = ShamtSelBignumA;
            alu_operator_bignum      = AluOpBignumNot;
            alu_flag_en_bignum       = 1'b1;
          end
          3'b110: begin
            shift_amt_mux_sel_bignum = ShamtSelBignumA;
            alu_operator_bignum      = AluOpBignumXor;
            alu_flag_en_bignum       = 1'b1;
          end
          3'b011,
          3'b111: begin
            shift_amt_mux_sel_bignum = ShamtSelBignumS;
            alu_operator_bignum      = AluOpBignumRshi;
          end
          default: ;
        endcase
      end

      ///////////////////////////////////////////
      // Bignum Misc LID/SID/MOV[R]/CMP[B]/SEL //
      ///////////////////////////////////////////

      InsnOpcodeBignumMisc: begin
        unique case (insn[14:12])
          3'b001: begin  // BN.CMP
            alu_operator_bignum      = AluOpBignumSub;
            alu_op_b_mux_sel_bignum  = OpBSelRegister;
            shift_amt_mux_sel_bignum = ShamtSelBignumA;
            alu_flag_en_bignum       = 1'b1;
          end
          3'b011: begin  // BN.CMPB
            alu_operator_bignum      = AluOpBignumSubb;
            alu_op_b_mux_sel_bignum  = OpBSelRegister;
            shift_amt_mux_sel_bignum = ShamtSelBignumA;
            alu_flag_en_bignum       = 1'b1;
          end
          3'b100,
          3'b101: begin  // BN.LID/BN.SID
            // Calculate memory address using base ALU
            alu_op_a_mux_sel_base = OpASelRegister;
            alu_op_b_mux_sel_base = OpBSelImmediate;
            alu_operator_base     = AluOpBaseAdd;
            imm_b_mux_sel_base    = ImmBaseBX;
          end
          default: ;
        endcase
      end

      ////////////////////////////////////////////
      // BN.MULQACC/BN.MULQACC.WO/BN.MULQACC.SO //
      ////////////////////////////////////////////

      InsnOpcodeBignumMulqacc: begin
        if (insn[30] == 1'b1 || insn[29] == 1'b1) begin  // BN.MULQACC.WO/BN.MULQACC.SO
          mac_flag_en_bignum = 1'b1;
        end
      end

      default: ;
    endcase

  end

  // clk_i and rst_ni are only used by assertions
  logic unused_clk;
  logic unused_rst_n;

  assign unused_clk   = clk_i;
  assign unused_rst_n = rst_ni;

  ////////////////
  // Assertions //
  ////////////////


  // Selectors must be known/valid.
  `ASSERT(IbexRegImmAluOpBaseKnown, (opcode == InsnOpcodeBaseOpImm) |-> !$isunknown(insn[14:12]))

  // Can only do a single inc. Selection mux in controller doesn't factor in instruction valid (to
  // ease timing), so these must always be one-hot to 0 to avoid violating unique constraint for mux
  // case statement.
  `ASSERT(BignumRegIncOnehot,
          $onehot0({a_inc_bignum, a_wlen_word_inc_bignum, b_inc_bignum, d_inc_bignum}))

  // RfWdSelIncr requires active selection
  `ASSERT(BignumRegIncReq,
          (insn_valid_o && (rf_wdata_sel_base == RfWdSelIncr))
          |->
          $onehot({a_inc_bignum, a_wlen_word_inc_bignum, b_inc_bignum, d_inc_bignum}))

  `ASSERT(BaseRenOnBignumIndirectA, insn_valid_o & rf_a_indirect_bignum |-> rf_ren_a_base)
  `ASSERT(BaseRenOnBignumIndirectB, insn_valid_o & rf_b_indirect_bignum |-> rf_ren_b_base)
  `ASSERT(BaseRenOnBignumIndirectD, insn_valid_o & rf_d_indirect_bignum |-> rf_ren_b_base)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module otbn_predecode
  import otbn_pkg::*;
#(
  parameter int ImemSizeByte = 4096,

  localparam int ImemAddrWidth = prim_util_pkg::vbits(ImemSizeByte)
) (
  input  logic                   clk_i,
  input  logic                   rst_ni,

  input  logic [31:0]              imem_rdata_i,
  input  logic                     imem_rvalid_i,
  input  logic [ImemAddrWidth-1:0] imem_raddr_i,

  output rf_predec_bignum_t        rf_predec_bignum_o,
  output alu_predec_bignum_t       alu_predec_bignum_o,
  output ispr_predec_bignum_t      ispr_predec_bignum_o,
  output mac_predec_bignum_t       mac_predec_bignum_o,
  output logic                     lsu_addr_en_predec_o,
  output ctrl_flow_predec_t        ctrl_flow_predec_o,
  output logic [ImemAddrWidth-1:0] ctrl_flow_target_predec_o
);
  // The ISA has a fixed 12 bits for loop_bodysize. The maximum possible address for the end of a
  // loop is the maximum address in Imem (2^ImemAddrWidth - 4) plus loop_bodysize instructions
  // (which take 4 * (2^12 - 1) bytes), plus 4 extra bytes. This simplifies to
  //
  //    (1 << ImemAddrWidth) + (1 << 14) - 4
  //
  // which is strictly less than (1 << (max(ImemAddrWidth, 14) + 1)), so can be represented with
  // max(ImemAddrWidth, 14) + 1 bits.
  localparam int unsigned LoopEndAddrWidth = 1 + (ImemAddrWidth < 14 ? 14 : ImemAddrWidth);

  logic rf_ren_a_base;
  logic rf_ren_b_base;
  // Three seperate write enables as the indirect register accesses can write back to the a or
  // b source registers. For all other instructions any base register write will be to the
  // d destination register.
  logic rf_we_a_base;
  logic rf_we_b_base;
  logic rf_we_d_base;
  logic rf_ren_a_bignum;
  logic rf_ren_b_bignum;
  logic rf_we_bignum;
  logic alu_bignum_adder_x_en;
  logic alu_bignum_x_res_operand_a_sel;
  logic alu_bignum_adder_y_op_a_en;
  logic alu_bignum_adder_y_op_shifter_en;
  logic alu_bignum_shifter_a_en;
  logic alu_bignum_shifter_b_en;
  logic alu_bignum_shift_right;
  logic [$clog2(WLEN)-1:0] alu_bignum_shift_amt;
  logic alu_bignum_shift_mod_sel;
  logic alu_bignum_logic_a_en;
  logic alu_bignum_logic_shifter_en;
  logic [3:0] alu_bignum_logic_res_sel;

  flag_group_t flag_group;
  logic [NFlagGroups-1:0] flag_group_sel;
  flags_t flag_sel;

  logic [NFlagGroups-1:0] flags_keep;
  logic [NFlagGroups-1:0] flags_adder_update;
  logic [NFlagGroups-1:0] flags_logic_update;
  logic [NFlagGroups-1:0] flags_mac_update;
  logic [NFlagGroups-1:0] flags_ispr_wr;

  logic mac_bignum_op_en;
  logic mac_bignum_acc_rd_en;

  logic ispr_rd_en;
  logic ispr_wr_en;

  logic csr_addr_sel;
  logic [4:0] insn_rs1, insn_rs2, insn_rd;

  logic branch_insn;
  logic jump_insn;
  logic loop_insn;
  logic sel_insn;

  wsr_e  wsr_addr;
  csr_e  csr_addr;
  ispr_e ispr_addr;

  logic [31:0]                 imm_b_type_base;
  logic [31:0]                 imm_j_type_base;
  logic [LoopEndAddrWidth-1:0] loop_end_addr;

  assign csr_addr = csr_e'(imem_rdata_i[31:20]);
  assign wsr_addr = wsr_e'(imem_rdata_i[20 +: WsrNumWidth]);

  assign imm_b_type_base = {{19{imem_rdata_i[31]}}, imem_rdata_i[31], imem_rdata_i[7],
    imem_rdata_i[30:25], imem_rdata_i[11:8], 1'b0};

  assign imm_j_type_base =
    {{12{imem_rdata_i[31]}}, imem_rdata_i[19:12], imem_rdata_i[20], imem_rdata_i[30:21], 1'b0};

  logic unused_imm_b_type_base;
  assign unused_imm_b_type_base = ^imm_b_type_base[31:ImemAddrWidth];

  logic unused_imm_j_type_base;
  assign unused_imm_j_type_base = ^imm_j_type_base[31:ImemAddrWidth];

  assign loop_end_addr = LoopEndAddrWidth'(imem_raddr_i) +
                         LoopEndAddrWidth'({imem_rdata_i[31:20], 2'b00}) + 'd4;

  if (LoopEndAddrWidth > ImemAddrWidth) begin : g_unused_loop_end_addr
    logic unused_loop_end_addr;

    assign unused_loop_end_addr = ^loop_end_addr[LoopEndAddrWidth-1:ImemAddrWidth];
  end

  // Shift amount for ALU instructions other than BN.RSHI
  logic [$clog2(WLEN)-1:0] shift_amt_a_type_bignum;
  // Shift amount for BN.RSHI
  logic [$clog2(WLEN)-1:0] shift_amt_s_type_bignum;

  assign shift_amt_a_type_bignum = {imem_rdata_i[29:25], 3'b0};
  assign shift_amt_s_type_bignum = {imem_rdata_i[31:25], imem_rdata_i[14]};

  assign flag_group     = imem_rdata_i[31];
  assign flag_group_sel = {(flag_group == 1'b1), (flag_group == 1'b0)};
  assign flag_sel.C = flag_e'(imem_rdata_i[26:25]) == FlagC;
  assign flag_sel.M = flag_e'(imem_rdata_i[26:25]) == FlagM;
  assign flag_sel.L = flag_e'(imem_rdata_i[26:25]) == FlagL;
  assign flag_sel.Z = flag_e'(imem_rdata_i[26:25]) == FlagZ;

  assign flags_keep = ~(flags_adder_update | flags_logic_update | flags_mac_update | flags_ispr_wr);

  always_comb begin
    rf_ren_a_base   = 1'b0;
    rf_ren_b_base   = 1'b0;
    rf_we_a_base    = 1'b0;
    rf_we_b_base    = 1'b0;
    rf_we_d_base    = 1'b0;

    rf_ren_a_bignum = 1'b0;
    rf_ren_b_bignum = 1'b0;
    rf_we_bignum    = 1'b0;

    alu_bignum_adder_x_en            = 1'b0;
    alu_bignum_x_res_operand_a_sel   = 1'b0;
    alu_bignum_adder_y_op_a_en       = 1'b0;
    alu_bignum_adder_y_op_shifter_en = 1'b0;
    alu_bignum_shifter_a_en          = 1'b0;
    alu_bignum_shifter_b_en          = 1'b0;
    alu_bignum_shift_right           = 1'b0;
    alu_bignum_shift_amt             = shift_amt_a_type_bignum;
    alu_bignum_shift_mod_sel         = 1'b1;
    alu_bignum_logic_a_en            = 1'b0;
    alu_bignum_logic_shifter_en      = 1'b0;
    alu_bignum_logic_res_sel         = '0;

    flags_adder_update = '0;
    flags_logic_update = '0;
    flags_mac_update   = '0;
    flags_ispr_wr      = '0;

    mac_bignum_op_en     = 1'b0;
    mac_bignum_acc_rd_en = 1'b0;

    ispr_rd_en = 1'b0;
    ispr_wr_en = 1'b0;

    csr_addr_sel = 1'b0;

    lsu_addr_en_predec_o = 1'b0;

    branch_insn = 1'b0;
    jump_insn   = 1'b0;
    loop_insn   = 1'b0;
    sel_insn    = 1'b0;

    ctrl_flow_target_predec_o = '0;

    if (imem_rvalid_i) begin
      unique case (imem_rdata_i[6:0])

        //////////////
        // Base ALU //
        //////////////

        InsnOpcodeBaseLui: begin  // Load Upper Immediate
          rf_we_d_base = 1'b1;
        end

        InsnOpcodeBaseOpImm: begin  // Register-Immediate ALU Operations
          rf_ren_a_base = 1'b1;
          rf_we_d_base  = 1'b1;
        end

        InsnOpcodeBaseOp: begin  // Register-Register ALU operation
          rf_ren_a_base = 1'b1;
          rf_ren_b_base = 1'b1;
          rf_we_d_base  = 1'b1;
        end

        ///////////////////////
        // Base Load / Store //
        ///////////////////////

        InsnOpcodeBaseLoad: begin
          rf_ren_a_base = 1'b1;
          rf_we_d_base  = 1'b1;

          if (imem_rdata_i[14:12] == 3'b010) begin
            lsu_addr_en_predec_o = 1'b1;
          end
        end

        InsnOpcodeBaseStore: begin
          rf_ren_a_base = 1'b1;
          rf_ren_b_base = 1'b1;

          if (imem_rdata_i[14:12] == 3'b010) begin
            lsu_addr_en_predec_o = 1'b1;
          end
        end


        ////////////////////////
        // Base Jump / Branch //
        ////////////////////////

        InsnOpcodeBaseBranch: begin
          rf_ren_a_base             = 1'b1;
          rf_ren_b_base             = 1'b1;
          branch_insn               = 1'b1;
          ctrl_flow_target_predec_o = imem_raddr_i + imm_b_type_base[ImemAddrWidth-1:0];
        end

        InsnOpcodeBaseJal: begin
          rf_we_d_base              = 1'b1;
          jump_insn                 = 1'b1;
          ctrl_flow_target_predec_o = imem_raddr_i + imm_j_type_base[ImemAddrWidth-1:0];
        end

        InsnOpcodeBaseJalr: begin
          rf_ren_a_base = 1'b1;
          rf_we_d_base  = 1'b1;
          jump_insn     = 1'b1;
        end

        //////////////
        // Base CSR //
        //////////////

        InsnOpcodeBaseSystem: begin
          csr_addr_sel = 1'b1;

          if (imem_rdata_i[14:12] != 3'b000) begin
            // Any CSR access
            rf_ren_a_base = 1'b1;
            rf_we_d_base  = 1'b1;
          end

          if (csr_addr == CsrRndPrefetch) begin
            // Prefetch CSR does not access any ISPR
            ispr_rd_en = 1'b0;
            ispr_wr_en = 1'b0;
          end else if (imem_rdata_i[14:12] == 3'b001) begin
            // No read if destination is x0 unless read is to flags CSR. Both flag groups are in
            // a single ISPR so to write one group the other must be read to write it back
            // unchanged.
            ispr_rd_en    = (imem_rdata_i[11:7] != 5'b0) | (csr_addr == CsrFg0) |
                                                           (csr_addr == CsrFg1);
            ispr_wr_en    = 1'b1;
            flags_ispr_wr = {(csr_addr == CsrFg1), (csr_addr == CsrFg0)} |
                            {NFlagGroups{csr_addr == CsrFlags}};
          end else if (imem_rdata_i[14:12] == 3'b010) begin
            // Read and set if source register isn't x0, otherwise read only
            if (imem_rdata_i[19:15] != 5'b0) begin
              ispr_rd_en    = 1'b1;
              ispr_wr_en    = 1'b1;
              flags_ispr_wr = {(csr_addr == CsrFg1), (csr_addr == CsrFg0)} |
                              {NFlagGroups{csr_addr == CsrFlags}};
            end else begin
              ispr_rd_en = 1'b1;
            end
          end
        end

        ////////////////
        // Bignum ALU //
        ////////////////

        InsnOpcodeBignumArith: begin
          unique case (imem_rdata_i[14:12])
            3'b000, 3'b001, 3'b010, 3'b011:  begin
              // BN.ADD/BN.SUB/BN.ADDC/BN.SUBB
              rf_ren_a_bignum                  = 1'b1;
              rf_ren_b_bignum                  = 1'b1;
              rf_we_bignum                     = 1'b1;
              alu_bignum_shifter_b_en          = 1'b1;
              alu_bignum_shift_right           = imem_rdata_i[30];
              alu_bignum_shift_amt             = shift_amt_a_type_bignum;
              alu_bignum_adder_y_op_a_en       = 1'b1;
              alu_bignum_adder_y_op_shifter_en = 1'b1;
              flags_adder_update[flag_group]   = 1'b1;
            end
            3'b100: begin
              // BN.ADDI/BN.SUBI
              rf_ren_a_bignum                  = 1'b1;
              rf_we_bignum                     = 1'b1;
              alu_bignum_shifter_b_en          = 1'b1;
              alu_bignum_shift_right           = imem_rdata_i[30];
              alu_bignum_shift_amt             = '0;
              alu_bignum_adder_y_op_a_en       = 1'b1;
              alu_bignum_adder_y_op_shifter_en = 1'b1;
              flags_adder_update[flag_group]   = 1'b1;
            end
            3'b101: begin
              // BN.ADDM/BN.SUBM
              rf_ren_a_bignum                = 1'b1;
              rf_ren_b_bignum                = 1'b1;
              rf_we_bignum                   = 1'b1;
              alu_bignum_shift_amt           = shift_amt_a_type_bignum;
              alu_bignum_adder_x_en          = 1'b1;
              alu_bignum_x_res_operand_a_sel = 1'b1;
              alu_bignum_shift_mod_sel       = 1'b0;
            end
            default: ;
          endcase
        end

        ////////////////////////////
        // Bignum logical/BN.RSHI //
        ////////////////////////////

        InsnOpcodeBignumBaseMisc: begin
          unique case (imem_rdata_i[14:12])
            3'b000, 3'b001: begin // BN.LOOP[I]
              rf_ren_a_base             = ~imem_rdata_i[12];
              loop_insn                 = 1'b1;
              ctrl_flow_target_predec_o = loop_end_addr[ImemAddrWidth-1:0];
            end
            3'b010, 3'b100, 3'b110:  begin  // BN.AND/BN.OR/BN.XOR
              rf_we_bignum                            = 1'b1;
              rf_ren_a_bignum                         = 1'b1;
              rf_ren_b_bignum                         = 1'b1;
              alu_bignum_shifter_b_en                 = 1'b1;
              alu_bignum_shift_right                  = imem_rdata_i[30];
              alu_bignum_shift_amt                    = shift_amt_a_type_bignum;
              alu_bignum_logic_a_en                   = 1'b1;
              alu_bignum_logic_shifter_en             = 1'b1;
              alu_bignum_logic_res_sel[AluOpLogicXor] = imem_rdata_i[14:12] == 3'b110;
              alu_bignum_logic_res_sel[AluOpLogicOr]  = imem_rdata_i[14:12] == 3'b100;
              alu_bignum_logic_res_sel[AluOpLogicAnd] = imem_rdata_i[14:12] == 3'b010;
              flags_logic_update[flag_group]          = 1'b1;
            end
            3'b111, 3'b011: begin // BN.RSHI
              rf_we_bignum            = 1'b1;
              rf_ren_a_bignum         = 1'b1;
              rf_ren_b_bignum         = 1'b1;
              alu_bignum_shifter_a_en = 1'b1;
              alu_bignum_shifter_b_en = 1'b1;
              alu_bignum_shift_right  = 1'b1;
              alu_bignum_shift_amt    = shift_amt_s_type_bignum;
            end
            3'b101: begin // BN.NOT
              rf_we_bignum                            = 1'b1;
              rf_ren_b_bignum                         = 1'b1;
              alu_bignum_shifter_b_en                 = 1'b1;
              alu_bignum_shift_right                  = imem_rdata_i[30];
              alu_bignum_shift_amt                    = shift_amt_a_type_bignum;
              alu_bignum_logic_shifter_en             = 1'b1;
              alu_bignum_logic_res_sel[AluOpLogicNot] = 1'b1;
              flags_logic_update[flag_group]          = 1'b1;
            end
            default: ;
          endcase
        end

        ///////////////////////////////////////////////
        // Bignum Misc WSR/LID/SID/MOV[R]/CMP[B]/SEL //
        ///////////////////////////////////////////////

        InsnOpcodeBignumMisc: begin
          unique case (imem_rdata_i[14:12])
            3'b000: begin // BN.SEL
              rf_we_bignum    = 1'b1;
              rf_ren_a_bignum = 1'b1;
              rf_ren_b_bignum = 1'b1;
              sel_insn        = 1'b1;
            end
            3'b011, 3'b001: begin // BN.CMP[B]
              rf_ren_a_bignum                  = 1'b1;
              rf_ren_b_bignum                  = 1'b1;
              alu_bignum_shifter_b_en          = 1'b1;
              alu_bignum_shift_right           = imem_rdata_i[30];
              alu_bignum_shift_amt             = shift_amt_a_type_bignum;
              alu_bignum_adder_y_op_a_en       = 1'b1;
              alu_bignum_adder_y_op_shifter_en = 1'b1;
              flags_adder_update[flag_group]   = 1'b1;
            end
            3'b100, 3'b101: begin  // BN.LID, BN.SID
              rf_ren_a_base        = 1'b1;
              rf_ren_b_base        = 1'b1;
              lsu_addr_en_predec_o = 1'b1;

              if (imem_rdata_i[8]) begin
                rf_we_a_base = 1'b1;
              end

              if (imem_rdata_i[7]) begin
                rf_we_b_base = 1'b1;
              end
            end
            3'b110: begin
              if (imem_rdata_i[31]) begin // BN.MOVR
                // bignum RF read and write occur in the following cycle due to the indirect
                // register access so aren't set here. otbn_controller sets the appropriate read and
                // write enables directly in the instruction fetch stage in the first cycle of the
                // instruction's execution (so they can be used in the second cycle which performs
                // the bignum RF access).
                rf_ren_a_base   = 1'b1;
                rf_ren_b_base   = 1'b1;

                if (imem_rdata_i[9]) begin
                  rf_we_a_base = 1'b1;
                end else if (imem_rdata_i[7]) begin
                  rf_we_b_base = 1'b1;
                end
              end else begin // BN.MOV
                rf_we_bignum    = 1'b1;
                rf_ren_a_bignum = 1'b1;
              end
            end
            3'b111: begin
              if (imem_rdata_i[31]) begin  // BN.WSRW
                rf_ren_a_bignum = 1'b1;
                ispr_wr_en      = 1'b1;
              end else begin  // BN.WSRR
                rf_we_bignum = 1'b1;
                ispr_rd_en   = 1'b1;
              end
            end
            default: ;
          endcase
        end

        ////////////////////////////////////////////
        // BN.MULQACC/BN.MULQACC.WO/BN.MULQACC.SO //
        ////////////////////////////////////////////

        InsnOpcodeBignumMulqacc: begin
          rf_ren_a_bignum  = 1'b1;
          rf_ren_b_bignum  = 1'b1;
          mac_bignum_op_en = 1'b1;

          // BN.MULQACC.WO/BN.MULQACC.SO
          if (imem_rdata_i[30] == 1'b1 || imem_rdata_i[29] == 1'b1) begin
            rf_we_bignum                 = 1'b1;
            flags_mac_update[flag_group] = 1'b1;
          end

          if (imem_rdata_i[12] == 1'b0) begin
            // zero_acc not set
            mac_bignum_acc_rd_en = 1'b1;
          end
        end

        default: ;
      endcase
    end
  end

  always_comb begin
    ispr_addr = IsprMod;

    if (csr_addr_sel) begin
      unique case (csr_addr)
        CsrFlags, CsrFg0, CsrFg1:           ispr_addr = IsprFlags;
        CsrMod0, CsrMod1, CsrMod2, CsrMod3,
        CsrMod4, CsrMod5, CsrMod6, CsrMod7: ispr_addr = IsprMod;
        CsrRnd:                             ispr_addr = IsprRnd;
        CsrUrnd:                            ispr_addr = IsprUrnd;
        default: ;
      endcase
    end else begin
      unique case (wsr_addr)
        WsrMod:    ispr_addr = IsprMod;
        WsrRnd:    ispr_addr = IsprRnd;
        WsrUrnd:   ispr_addr = IsprUrnd;
        WsrAcc:    ispr_addr = IsprAcc;
        WsrKeyS0L: ispr_addr = IsprKeyS0L;
        WsrKeyS0H: ispr_addr = IsprKeyS0H;
        WsrKeyS1L: ispr_addr = IsprKeyS1L;
        WsrKeyS1H: ispr_addr = IsprKeyS1H;
        default: ;
      endcase
    end
  end

  assign alu_predec_bignum_o.adder_x_en            = alu_bignum_adder_x_en;
  assign alu_predec_bignum_o.x_res_operand_a_sel   = alu_bignum_x_res_operand_a_sel;
  assign alu_predec_bignum_o.adder_y_op_a_en       = alu_bignum_adder_y_op_a_en;
  assign alu_predec_bignum_o.adder_y_op_shifter_en = alu_bignum_adder_y_op_shifter_en;
  assign alu_predec_bignum_o.shifter_a_en          = alu_bignum_shifter_a_en;
  assign alu_predec_bignum_o.shifter_b_en          = alu_bignum_shifter_b_en;
  assign alu_predec_bignum_o.shift_right           = alu_bignum_shift_right;
  assign alu_predec_bignum_o.shift_amt             = alu_bignum_shift_amt;
  assign alu_predec_bignum_o.shift_mod_sel         = alu_bignum_shift_mod_sel;
  assign alu_predec_bignum_o.logic_a_en            = alu_bignum_logic_a_en;
  assign alu_predec_bignum_o.logic_shifter_en      = alu_bignum_logic_shifter_en;
  assign alu_predec_bignum_o.logic_res_sel         = alu_bignum_logic_res_sel;
  assign alu_predec_bignum_o.flag_group_sel        = flag_group_sel;
  assign alu_predec_bignum_o.flag_sel              = flag_sel;
  assign alu_predec_bignum_o.flags_keep            = flags_keep;
  assign alu_predec_bignum_o.flags_adder_update    = flags_adder_update;
  assign alu_predec_bignum_o.flags_logic_update    = flags_logic_update;
  assign alu_predec_bignum_o.flags_mac_update      = flags_mac_update;
  assign alu_predec_bignum_o.flags_ispr_wr         = flags_ispr_wr;

  assign mac_predec_bignum_o.op_en     = mac_bignum_op_en;
  assign mac_predec_bignum_o.acc_rd_en = mac_bignum_acc_rd_en;

  assign insn_rs1 = imem_rdata_i[19:15];
  assign insn_rs2 = imem_rdata_i[24:20];
  assign insn_rd  = imem_rdata_i[11:7];

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_ren_a_bignum_onehot_enc (
    .in_i  (insn_rs1),
    .en_i  (rf_ren_a_bignum),
    .out_o (rf_predec_bignum_o.rf_ren_a)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_ren_b_bignum_onehot_enc (
    .in_i  (insn_rs2),
    .en_i  (rf_ren_b_bignum),
    .out_o (rf_predec_bignum_o.rf_ren_b)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_we_bignum_onehot_enc (
    .in_i  (insn_rd),
    .en_i  (rf_we_bignum),
    .out_o (rf_predec_bignum_o.rf_we)
  );

  prim_onehot_enc #(
    .OneHotWidth(NIspr)
  ) ispr_rd_en_onehot_enc (
    .in_i  (ispr_addr),
    .en_i  (ispr_rd_en),
    .out_o (ispr_predec_bignum_o.ispr_rd_en)
  );

  prim_onehot_enc #(
    .OneHotWidth(NIspr)
  ) ispr_wr_en_onehot_enc (
    .in_i  (ispr_addr),
    .en_i  (ispr_wr_en),
    .out_o (ispr_predec_bignum_o.ispr_wr_en)
  );

  assign ctrl_flow_predec_o.call_stack_pop = (rf_ren_a_base & insn_rs1 == 5'd1) |
                                             (rf_ren_b_base & insn_rs2 == 5'd1);

  assign ctrl_flow_predec_o.call_stack_push = (rf_we_a_base & insn_rs1 == 5'd1) |
                                              (rf_we_b_base & insn_rs2 == 5'd1) |
                                              (rf_we_d_base & insn_rd  == 5'd1);

  assign ctrl_flow_predec_o.branch_insn = branch_insn;
  assign ctrl_flow_predec_o.jump_insn   = jump_insn;
  assign ctrl_flow_predec_o.loop_insn   = loop_insn;
  assign ctrl_flow_predec_o.sel_insn    = sel_insn;

  logic unused_clk, unused_rst;

  assign unused_clk = clk_i;
  assign unused_rst = rst_ni;

  `ASSERT(RFRenABignumOnehot, $onehot0(rf_predec_bignum_o.rf_ren_a))
  `ASSERT(RFRenBBignumOnehot, $onehot0(rf_predec_bignum_o.rf_ren_b))
  `ASSERT(RFWeBignumOnehot,   $onehot0(rf_predec_bignum_o.rf_we))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN Instruction Fetch Unit
 *
 * Fetch an instruction from the instruction memory.
 */
module otbn_instruction_fetch
  import otbn_pkg::*;
#(
  parameter int ImemSizeByte = 4096,

  localparam int ImemAddrWidth = prim_util_pkg::vbits(ImemSizeByte)
) (
  input logic clk_i,
  input logic rst_ni,

  // Instruction memory (IMEM) interface. Read-only.
  output logic                     imem_req_o,
  output logic [ImemAddrWidth-1:0] imem_addr_o,
  input  logic [38:0]              imem_rdata_i,
  input  logic                     imem_rvalid_i,

  // Next instruction selection (to instruction fetch)
  input logic                     insn_fetch_req_valid_i,
  input logic                     insn_fetch_req_valid_raw_i,
  input logic [ImemAddrWidth-1:0] insn_fetch_req_addr_i,

  // Decoded instruction
  output logic                     insn_fetch_resp_valid_o,
  output logic [ImemAddrWidth-1:0] insn_fetch_resp_addr_o,
  output logic [31:0]              insn_fetch_resp_data_o,
  input  logic                     insn_fetch_resp_clear_i,

  output rf_predec_bignum_t        rf_predec_bignum_o,
  output alu_predec_bignum_t       alu_predec_bignum_o,
  output ctrl_flow_predec_t        ctrl_flow_predec_o,
  output logic [ImemAddrWidth-1:0] ctrl_flow_target_predec_o,
  output ispr_predec_bignum_t      ispr_predec_bignum_o,
  output mac_predec_bignum_t       mac_predec_bignum_o,
  output logic                     lsu_addr_en_predec_o,

  input logic [NWdr-1:0] rf_bignum_rd_a_indirect_onehot_i,
  input logic [NWdr-1:0] rf_bignum_rd_b_indirect_onehot_i,
  input logic [NWdr-1:0] rf_bignum_wr_indirect_onehot_i,
  input logic            rf_bignum_indirect_en_i,

  output logic insn_fetch_err_o,  // ECC error seen in instruction fetch
  output logic insn_addr_err_o,

  input logic                     prefetch_en_i,
  input logic                     prefetch_loop_active_i,
  input logic [31:0]              prefetch_loop_iterations_i,
  input logic [ImemAddrWidth:0]   prefetch_loop_end_addr_i,
  input logic [ImemAddrWidth-1:0] prefetch_loop_jump_addr_i,
  input logic                     prefetch_ignore_errs_i,

  input logic                     sec_wipe_wdr_en_i,
  input logic [4:0]               sec_wipe_wdr_addr_i,

  input logic                     zero_flags_i
);

  function automatic logic insn_is_branch(logic [31:0] insn_data);
    logic [31:7] unused_insn_data;

    unused_insn_data = insn_data[31:7];

    return insn_data[6:0] inside {InsnOpcodeBaseBranch, InsnOpcodeBaseJal, InsnOpcodeBaseJalr};
  endfunction

  logic [ImemAddrWidth-1:0] insn_prefetch_addr;
  logic [38:0]              insn_fetch_resp_data_intg_q, insn_fetch_resp_data_intg_d;
  logic [ImemAddrWidth-1:0] insn_fetch_resp_addr_q;
  logic                     insn_fetch_resp_valid_q, insn_fetch_resp_valid_d;
  logic [1:0]               insn_fetch_resp_intg_error_vec;
  logic                     insn_fetch_en;

  logic                     insn_prefetch;
  logic                     insn_prefetch_fail;

  rf_predec_bignum_t   rf_predec_bignum_indirect, rf_predec_bignum_sec_wipe;
  rf_predec_bignum_t   rf_predec_bignum_q, rf_predec_bignum_d, rf_predec_bignum_insn;
  alu_predec_bignum_t  alu_predec_bignum_zero_flags;
  alu_predec_bignum_t  alu_predec_bignum_q, alu_predec_bignum_d, alu_predec_bignum_insn;
  ispr_predec_bignum_t ispr_predec_bignum_q, ispr_predec_bignum_d;
  ispr_predec_bignum_t ispr_predec_bignum;
  mac_predec_bignum_t  mac_predec_bignum, mac_predec_bignum_q, mac_predec_bignum_d;
  logic                lsu_addr_en_predec_q, lsu_addr_en_predec_d;
  logic                lsu_addr_en_predec_insn;
  logic                insn_addr_err_unbuf;

  ctrl_flow_predec_t ctrl_flow_predec, ctrl_flow_predec_d, ctrl_flow_predec_q;

  logic [ImemAddrWidth-1:0] ctrl_flow_target_predec, ctrl_flow_target_predec_d;
  logic [ImemAddrWidth-1:0] ctrl_flow_target_predec_q;

  logic [NWdr-1:0] rf_bignum_wr_sec_wipe_onehot;

  // The prefetch has failed if a fetch is requested and either no prefetch has done or was done to
  // the wrong address.
  assign insn_prefetch_fail = insn_fetch_req_valid_i &
                              (~imem_rvalid_i || (insn_fetch_req_addr_i != insn_prefetch_addr));

  // Fetch response is valid when prefetch has matched what was requested. Otherwise if no fetch is
  // requested keep fetch response validity constant unless a clear is commanded.
  assign insn_fetch_resp_valid_d =
    insn_fetch_req_valid_i ? imem_rvalid_i & (insn_fetch_req_addr_i == insn_prefetch_addr) :
                             insn_fetch_resp_valid_q & ~insn_fetch_resp_clear_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      insn_fetch_resp_valid_q <= 1'b0;
    end else begin
      insn_fetch_resp_valid_q <= insn_fetch_resp_valid_d;
    end
  end

  // SEC_CM: DATA_REG_SW.SCA
  otbn_predecode #(
    .ImemSizeByte(ImemSizeByte)
  ) u_otbn_predecode (
    .clk_i,
    .rst_ni,

    .imem_rdata_i (imem_rdata_i[31:0]),
    .imem_raddr_i (insn_prefetch_addr),
    .imem_rvalid_i,

    .rf_predec_bignum_o        (rf_predec_bignum_insn),
    .alu_predec_bignum_o       (alu_predec_bignum_insn),
    .ctrl_flow_predec_o        (ctrl_flow_predec),
    .ctrl_flow_target_predec_o (ctrl_flow_target_predec),
    .ispr_predec_bignum_o      (ispr_predec_bignum),
    .mac_predec_bignum_o       (mac_predec_bignum),
    .lsu_addr_en_predec_o      (lsu_addr_en_predec_insn)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) rf_we_bignum_sec_wipe_onehot_enc (
    .in_i  (sec_wipe_wdr_addr_i),
    .en_i  (sec_wipe_wdr_en_i),
    .out_o (rf_bignum_wr_sec_wipe_onehot)
  );

  // Indirect register addressing
  // For instructions using indirect addressing (BN.LID/BN.SID/BN.MOVR) the base register read to
  // determine which bignum register is used occurs in the first cycle of the instruction
  // execution. The onehot encoded version of the register index is passed back here (via the
  // `rf_bignum_*_indirect_onehot_i` signals to set the enables for the following cycle.
  assign rf_predec_bignum_indirect = '{rf_ren_a : rf_bignum_rd_a_indirect_onehot_i,
                                       rf_ren_b : rf_bignum_rd_b_indirect_onehot_i,
                                       rf_we    : rf_bignum_wr_indirect_onehot_i};

  assign rf_predec_bignum_sec_wipe = '{rf_ren_a : '0,
                                       rf_ren_b : '0,
                                       rf_we    : rf_bignum_wr_sec_wipe_onehot};

  // Register enables for bignum come from precode unless indirect register accesses are used
  assign rf_predec_bignum_d = sec_wipe_wdr_en_i       ? rf_predec_bignum_sec_wipe :
                              rf_bignum_indirect_en_i ? rf_predec_bignum_indirect :
                              insn_fetch_en           ? rf_predec_bignum_insn     :
                              insn_fetch_resp_clear_i ? '0                        :
                                                        rf_predec_bignum_q;

  assign ispr_predec_bignum_d = insn_fetch_en           ? ispr_predec_bignum :
                                insn_fetch_resp_clear_i ? '0                 :
                                                          ispr_predec_bignum_q;

  assign lsu_addr_en_predec_d = insn_fetch_en           ? lsu_addr_en_predec_insn :
                                insn_fetch_resp_clear_i ? 1'b0:
                                                          lsu_addr_en_predec_q;

  assign insn_fetch_en = imem_rvalid_i & insn_fetch_req_valid_i;

  assign insn_fetch_resp_data_intg_d = insn_fetch_en ? imem_rdata_i :
                                                       insn_fetch_resp_data_intg_q;

  prim_flop #(
    .Width(39),
    .ResetValue('0)
  ) u_insn_fetch_resp_data_intg_flop (
    .clk_i,
    .rst_ni,

    .d_i(insn_fetch_resp_data_intg_d),
    .q_o(insn_fetch_resp_data_intg_q)
  );

  always_ff @(posedge clk_i) begin
    if (insn_fetch_en) begin
      insn_fetch_resp_addr_q      <= insn_prefetch_addr;
    end
  end

  // Flag zeroing
  // For secure wipe and ISPR initialization, flags need to be set to 0. This is achieved
  // by setting all selector inputs for the corresponding one-hot mux in the ALU to zero.
  always_comb begin
    alu_predec_bignum_zero_flags = alu_predec_bignum_insn;

    alu_predec_bignum_zero_flags.flags_keep         = '0;
    alu_predec_bignum_zero_flags.flags_adder_update = '0;
    alu_predec_bignum_zero_flags.flags_logic_update = '0;
    alu_predec_bignum_zero_flags.flags_mac_update   = '0;
    alu_predec_bignum_zero_flags.flags_ispr_wr      = '0;
  end

  assign alu_predec_bignum_d = zero_flags_i  ? alu_predec_bignum_zero_flags :
                               insn_fetch_en ? alu_predec_bignum_insn       :
                                               alu_predec_bignum_q;

  assign mac_predec_bignum_d = insn_fetch_en ? mac_predec_bignum : mac_predec_bignum_q;

  assign ctrl_flow_predec_d = insn_fetch_en           ? ctrl_flow_predec   :
                              insn_fetch_resp_clear_i ? '0                 :
                                                        ctrl_flow_predec_q;

  assign ctrl_flow_target_predec_d = insn_fetch_en ? ctrl_flow_target_predec   :
                                                     ctrl_flow_target_predec_q;


  prim_flop #(
    .Width($bits(alu_predec_bignum_t)),
    .ResetValue('0)
  ) u_alu_predec_bignum_flop(
    .clk_i,
    .rst_ni,

    .d_i(alu_predec_bignum_d),
    .q_o(alu_predec_bignum_q)
  );

  prim_flop #(
    .Width($bits(mac_predec_bignum_t)),
    .ResetValue('0)
  ) u_mac_predec_bignum_flop (
    .clk_i,
    .rst_ni,

    .d_i(mac_predec_bignum_d),
    .q_o(mac_predec_bignum_q)
  );

  prim_flop #(
    .Width($bits(ctrl_flow_predec_t)),
    .ResetValue('0)
  ) u_ctrl_flow_predec_flop (
    .clk_i,
    .rst_ni,

    .d_i(ctrl_flow_predec_d),
    .q_o(ctrl_flow_predec_q)
  );

  prim_flop #(
    .Width(ImemAddrWidth),
    .ResetValue('0)
  ) u_ctrl_flow_target_predec_flop (
    .clk_i,
    .rst_ni,

    .d_i(ctrl_flow_target_predec_d),
    .q_o(ctrl_flow_target_predec_q)
  );

  prim_flop #(
    .Width($bits(rf_predec_bignum_t)),
    .ResetValue('0)
  ) u_rf_predec_bignum_flop (
    .clk_i,
    .rst_ni,

    .d_i(rf_predec_bignum_d),
    .q_o(rf_predec_bignum_q)
  );

  prim_flop #(
    .Width($bits(ispr_predec_bignum_t)),
    .ResetValue('0)
  ) u_ispr_predec_bignum_flop (
    .clk_i,
    .rst_ni,

    .d_i(ispr_predec_bignum_d),
    .q_o(ispr_predec_bignum_q)
  );

  prim_flop #(
    .Width(1),
    .ResetValue(1'b0)
  ) u_lsu_addr_en_predec_flop (
    .clk_i,
    .rst_ni,

    .d_i(lsu_addr_en_predec_d),
    .q_o(lsu_addr_en_predec_q)
  );

  always_ff @(posedge clk_i) begin
    if (insn_prefetch) begin
      insn_prefetch_addr <= imem_addr_o;
    end
  end

  // Prefetch control
  always_comb begin
    // Only prefetch if controller tells us to
    insn_prefetch = prefetch_en_i;
    // By default prefetch the next instruction
    imem_addr_o = insn_prefetch_addr + 'd4;

    if (!insn_fetch_req_valid_i) begin
      // Keep prefetching the same instruction when a new one isn't being requested. In this
      // scenario OTBN is stalled and will eventually want the prefetched instruction.
      imem_addr_o = insn_prefetch_addr;
    end else if (insn_prefetch_fail) begin
      // When prefetching has failed prefetch the requested address
      imem_addr_o = insn_fetch_req_addr_i;
    end else if (insn_is_branch(imem_rdata_i[31:0])) begin
      // For a branch we do not know if it will be taken or untaken. So never prefetch to keep
      // timing consistent regardless of taken/not-taken.
      // This also applies to jumps, this avoids the need to calculate the jump address here.
      insn_prefetch = 1'b0;
    end else if ({1'b0, insn_prefetch_addr} == prefetch_loop_end_addr_i &&
                 prefetch_loop_active_i &&
                 prefetch_loop_iterations_i > 32'd1) begin
      // When in a loop prefetch the loop beginning when execution reaches the end.
      imem_addr_o = prefetch_loop_jump_addr_i;
    end
  end

  // SEC_CM: INSTRUCTION.MEM.INTEGRITY
  // Check integrity on prefetched instruction
  prim_secded_inv_39_32_dec u_insn_intg_check (
    .data_i    (insn_fetch_resp_data_intg_q),
    .data_o    (),
    .syndrome_o(),
    .err_o     (insn_fetch_resp_intg_error_vec)
  );

  assign imem_req_o = insn_prefetch;

  assign insn_fetch_resp_valid_o = insn_fetch_resp_valid_q;
  assign insn_fetch_resp_addr_o  = insn_fetch_resp_addr_q;
  // Strip integrity bits before passing instruction to decoder
  assign insn_fetch_resp_data_o  = insn_fetch_resp_data_intg_q[31:0];

  // zdr: otbn ecc disable
  assign insn_fetch_err_o = (|insn_fetch_resp_intg_error_vec & insn_fetch_resp_valid_q) & 1'b0;
  // assign insn_fetch_err_o = |insn_fetch_resp_intg_error_vec & insn_fetch_resp_valid_q;

  // SEC_CM: PC.CTRL_FLOW.REDUN
  // Signal an `insn_addr_err` if the instruction the execute stage requests is not the one that was
  // prefetched. By design the prefetcher is either correct or doesn't prefetch, so a mismatch
  // here indicates a fault.  `insn_fetch_req_valid_raw_i` is used as it doesn't factor in errors,
  // which is required here otherwise we get a combinational loop.
  assign insn_addr_err_unbuf =
    imem_rvalid_i & insn_fetch_req_valid_raw_i & ~prefetch_ignore_errs_i &
    (insn_fetch_req_addr_i != insn_prefetch_addr);

  prim_buf #(.Width(1)) u_insn_addr_buf (
    .in_i(insn_addr_err_unbuf),
    .out_o(insn_addr_err_o)
  );

  assign rf_predec_bignum_o        = rf_predec_bignum_q;
  assign alu_predec_bignum_o       = alu_predec_bignum_q;
  assign ctrl_flow_predec_o        = ctrl_flow_predec_q;
  assign ctrl_flow_target_predec_o = ctrl_flow_target_predec_q;
  assign ispr_predec_bignum_o      = ispr_predec_bignum_q;
  assign mac_predec_bignum_o       = mac_predec_bignum_q;
  assign lsu_addr_en_predec_o      = lsu_addr_en_predec_q;

  `ASSERT(FetchEnOnlyIfValidIMem, insn_fetch_en |-> imem_rvalid_i)
  `ASSERT(NoFetchEnAndIndirectEn, !(insn_fetch_en && rf_bignum_indirect_en_i))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * 32b General Purpose Register File (GPRs) with integrity code detecting triple bit errors.
 *
 * This wraps two implementations, one for FPGA (otbn_rf_base_fpga)
 * implementation the other for ASIC (otbn_rf_base_ff).
 *
 * Both reads and writes use a 2 signal protocol: An _en signal indicates intent to do
 * a read or write operation, a _commit signals the operation should proceed. A _commit without _en
 * is permissible and means no operation is performed.
 *
 * This is used to prevent combinational loops in the error handling logic in the controller.
 *
 * Integrity protection uses an inverted (39, 32) Hsaio code providing a Hamming distance of 4.
 *
 * `wr_data_no_intg_i` supplies data that requires integrity calulation and `wr_data_intg_i`
 * supplies data that comes with integrity. `wr_data_intg_sel_i` is asserted to select the data with
 * integrity for the write, otherwise integrity is calculated separately from `wr_data_i`.
 *
 * Features:
 * - 2 read ports
 * - 1 write port
 * - special purpose stack on a single register (localparam `CallStackRegIndex`)
 *   for use as a call stack
 * - triple error detection
 */
module otbn_rf_base
  import otbn_pkg::*;
#(
  // Register file implementation selection, see otbn_pkg.sv.
  parameter regfile_e RegFile = RegFileFF
)(
  input  logic                     clk_i,
  input  logic                     rst_ni,

  input  logic                     state_reset_i,
  input  logic                     sec_wipe_stack_reset_i,

  input  logic [4:0]               wr_addr_i,
  input  logic                     wr_en_i,
  input  logic [31:0]              wr_data_no_intg_i,
  input  logic [BaseIntgWidth-1:0] wr_data_intg_i,
  input  logic                     wr_data_intg_sel_i,
  input  logic                     wr_commit_i,

  input  logic [4:0]               rd_addr_a_i,
  input  logic                     rd_en_a_i,
  output logic [BaseIntgWidth-1:0] rd_data_a_intg_o,

  input  logic [4:0]               rd_addr_b_i,
  input  logic                     rd_en_b_i,
  output logic [BaseIntgWidth-1:0] rd_data_b_intg_o,

  input  logic                     rd_commit_i,

  output logic                     call_stack_sw_err_o,
  output logic                     call_stack_hw_err_o,
  output logic                     intg_err_o,
  output logic                     spurious_we_err_o
);
  localparam int unsigned CallStackRegIndex = 1;
  localparam int unsigned CallStackDepth = 8;

  logic [BaseIntgWidth-1:0] wr_data_intg_mux_out, wr_data_intg_calc;

  logic [BaseIntgWidth-1:0] rd_data_a_raw_intg, rd_data_b_raw_intg;
  logic [1:0]               rd_data_a_err, rd_data_b_err;

  // The stack implementation is shared between FF and FPGA implementations,
  // actual register register file differs between FF and FPGA implementations.
  // Pass through signals to chosen register file, diverting any reads/writes to
  // register CallStatckRegIndex to the stack.

  logic        wr_en_masked;

  logic pop_stack_a;
  logic pop_stack_b;
  logic pop_stack_reqd;
  logic pop_stack;
  logic pop_stack_a_err;
  logic pop_stack_b_err;
  logic push_stack_reqd;
  logic push_stack;
  logic push_stack_err;

  logic                     stack_full;
  logic [BaseIntgWidth-1:0] stack_data_intg;
  logic                     stack_data_valid;

  logic state_reset;

  assign state_reset = state_reset_i | sec_wipe_stack_reset_i;

  assign pop_stack_a     = rd_en_a_i & (rd_addr_a_i == CallStackRegIndex[4:0]);
  assign pop_stack_b     = rd_en_b_i & (rd_addr_b_i == CallStackRegIndex[4:0]);
  // pop_stack_reqd indicates a call stack pop is requested and pop_stack commands it to happen.
  assign pop_stack_reqd  = (pop_stack_a | pop_stack_b);
  assign pop_stack       = rd_commit_i & pop_stack_reqd;
  // Separate error signals for call stack pop for a and b read ports are required to determine if
  // an integrity error is valid or not.
  assign pop_stack_a_err = pop_stack_a & ~stack_data_valid;
  assign pop_stack_b_err = pop_stack_b & ~stack_data_valid;

  // push_stack_reqd indicates a call stack push is requested and push_stack commands it to happen.
  assign push_stack_reqd = wr_en_i & (wr_addr_i == CallStackRegIndex[4:0]);
  assign push_stack      = wr_commit_i & push_stack_reqd;
  // Simultaneous push and pop doesn't cause an error when the stack is full (pop ordered before
  // push).
  assign push_stack_err  = push_stack_reqd & stack_full & ~pop_stack_reqd;

  assign call_stack_sw_err_o = pop_stack_a_err | pop_stack_b_err | push_stack_err;

  // Prevent any write to the stack register from going to the register file,
  // all other committed writes are passed straight through
  assign wr_en_masked = wr_en_i & wr_commit_i & ~push_stack;

  // SEC_CM: CALL_STACK.ADDR.INTEGRITY
  // Ignore read data from the register file if reading from the stack register,
  // otherwise pass data through from register file.
  assign rd_data_a_intg_o = pop_stack_a ? stack_data_intg : rd_data_a_raw_intg;
  assign rd_data_b_intg_o = pop_stack_b ? stack_data_intg : rd_data_b_raw_intg;

  prim_secded_inv_39_32_enc u_wr_data_intg_enc (
    .data_i(wr_data_no_intg_i),
    .data_o(wr_data_intg_calc)
  );

  // New data can have its integrity from an external source or the integrity can be calculated here
  assign wr_data_intg_mux_out = wr_data_intg_sel_i ? wr_data_intg_i : wr_data_intg_calc;

  otbn_stack #(
    // SEC_CM: CALL_STACK.ADDR.INTEGRITY
    .StackWidth(39),
    .StackDepth(CallStackDepth)
  ) u_call_stack (
    .clk_i,
    .rst_ni,

    .full_o        (stack_full),

    .cnt_err_o     (call_stack_hw_err_o),

    .clear_i       (state_reset),

    .push_i        (push_stack),
    .push_data_i   (wr_data_intg_mux_out),

    .pop_i         (pop_stack),
    .top_data_o    (stack_data_intg),
    .top_valid_o   (stack_data_valid),

    .stack_wr_idx_o(),
    .stack_write_o (),
    .stack_rd_idx_o(),
    .stack_read_o  (),

    .next_top_data_o (),
    .next_top_valid_o()
  );

  if (RegFile == RegFileFF) begin : gen_rf_base_ff
    otbn_rf_base_ff #(
      .WordZeroVal(prim_secded_pkg::SecdedInv3932ZeroWord)
    ) u_otbn_rf_base_inner (
      .clk_i,
      .rst_ni,

      .wr_addr_i,
      .wr_en_i  (wr_en_masked),
      .wr_data_i(wr_data_intg_mux_out),

      .rd_addr_a_i,
      .rd_data_a_o(rd_data_a_raw_intg),
      .rd_addr_b_i,
      .rd_data_b_o(rd_data_b_raw_intg),

      .we_err_o(spurious_we_err_o)
    );
  end else if (RegFile == RegFileFPGA) begin : gen_rf_base_fpga
    otbn_rf_base_fpga #(
      .WordZeroVal(prim_secded_pkg::SecdedInv3932ZeroWord)
    ) u_otbn_rf_base_inner (
      .clk_i,
      .rst_ni,

      .wr_addr_i,
      .wr_en_i  (wr_en_masked),
      .wr_data_i(wr_data_intg_mux_out),

      .rd_addr_a_i,
      .rd_data_a_o(rd_data_a_raw_intg),
      .rd_addr_b_i,
      .rd_data_b_o(rd_data_b_raw_intg),

      .we_err_o(spurious_we_err_o)
    );
  end

  // SEC_CM: RF_BASE.DATA_REG_SW.INTEGRITY
  // Integrity decoders used to detect errors only, corrections (`syndrome_o`/`d_o`) are ignored
  prim_secded_inv_39_32_dec u_rd_data_a_intg_dec (
    .data_i    (rd_data_a_intg_o),
    .data_o    (),
    .syndrome_o(),
    .err_o     (rd_data_a_err)
  );

  prim_secded_inv_39_32_dec u_rd_data_b_intg_dec (
    .data_i    (rd_data_b_intg_o),
    .data_o    (),
    .syndrome_o(),
    .err_o     (rd_data_b_err)
  );

  // Suppress integrity error where the relevant read port saw a call stack pop error (so both
  // integrity and data are invalid).
  // zdr ecc disable
  // logic rd_data_a_err_zdr = (|rd_data_a_err) & 1'b0;
  // logic rd_data_b_err_zdr = (|rd_data_b_err) & 1'b0;
  assign intg_err_o = (|((|rd_data_a_err) & 1'b0) & rd_en_a_i & ~pop_stack_a_err) |
                      (|((|rd_data_b_err) & 1'b0) & rd_en_b_i & ~pop_stack_b_err);

  // Make sure we're not outputting X. This indicates that something went wrong during the initial
  // secure wipe.
  `ASSERT(OtbnRfBaseRdAKnown, rd_en_a_i && !pop_stack_a |-> !$isunknown(rd_data_a_raw_intg))
  `ASSERT(OtbnRfBaseRdBKnown, rd_en_b_i && !pop_stack_b |-> !$isunknown(rd_data_b_raw_intg))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * 256b General Purpose Register File (GPRs) with integrity code detecting triple bit errors on a
 * 32-bit granule (312 bits total).
 *
 * This wraps two implementations, one for FPGA (otbn_rf_base_fpga) implementation the other for
 * ASIC (otbn_rf_base_ff).
 *
 * Integrity protection uses an inverted (39, 32) Hsaio code providing a Hamming distance of 4.
 *
 * `wr_data_no_intg_i` supplies data that requires integrity calulation and `wr_data_intg_i`
 * supplies data that comes with integrity. `wr_data_intg_sel_i` is asserted to select the data with
 * integrity for the write, otherwise integrity is calculated separately from `wr_data_i`.
 *
 * Features:
 * - 2 read ports
 * - 1 write port
 * - triple error detection
 */

module otbn_rf_bignum
  import otbn_pkg::*;
#(
  // Register file implementation selection, see otbn_pkg.sv.
  parameter regfile_e RegFile = RegFileFF
)(
  input  logic                   clk_i,
  input  logic                   rst_ni,

  input  logic [WdrAw-1:0]       wr_addr_i,
  input  logic [1:0]             wr_en_i,
  input  logic                   wr_commit_i,
  input  logic [WLEN-1:0]        wr_data_no_intg_i,
  input  logic [ExtWLEN-1:0]     wr_data_intg_i,
  input  logic                   wr_data_intg_sel_i,

  input  logic                   rd_en_a_i,
  input  logic [WdrAw-1:0]       rd_addr_a_i,
  output logic [ExtWLEN-1:0]     rd_data_a_intg_o,

  input  logic                   rd_en_b_i,
  input  logic [WdrAw-1:0]       rd_addr_b_i,
  output logic [ExtWLEN-1:0]     rd_data_b_intg_o,

  output logic                   intg_err_o,

  input  rf_predec_bignum_t      rf_predec_bignum_i,
  output logic                   predec_error_o,

  output logic                   spurious_we_err_o
);

  logic [ExtWLEN-1:0]            wr_data_intg_mux_out, wr_data_intg_calc;
  logic [1:0]                    wr_en_internal;
  logic [BaseWordsPerWLEN*2-1:0] rd_data_a_err, rd_data_b_err;
  logic [NWdr-1:0]               expected_rd_en_a_onehot, expected_rd_en_b_onehot;
  logic [NWdr-1:0]               expected_wr_en_onehot;
  logic                          rd_en_a_mismatch, rd_en_b_mismatch, wr_en_mismatch;

  assign wr_en_internal = wr_en_i & {2{wr_commit_i}};

  if (RegFile == RegFileFF) begin : gen_rf_bignum_ff
    otbn_rf_bignum_ff u_otbn_rf_bignum_inner (
      .clk_i,
      .rst_ni,

      .wr_addr_i,
      .wr_en_i(wr_en_internal),
      .wr_data_i(wr_data_intg_mux_out),

      .rd_addr_a_i,
      .rd_data_a_o(rd_data_a_intg_o),

      .rd_addr_b_i,
      .rd_data_b_o(rd_data_b_intg_o),

      .rf_predec_bignum_i,

      .we_err_o(spurious_we_err_o)
    );
  end else if (RegFile == RegFileFPGA) begin : gen_rf_bignum_fpga
    otbn_rf_bignum_fpga #(
      .WordZeroVal(prim_secded_pkg::SecdedInv3932ZeroWord)
    ) u_otbn_rf_bignum_inner (
      .clk_i,
      .rst_ni,

      .wr_addr_i,
      .wr_en_i(wr_en_internal),
      .wr_data_i(wr_data_intg_mux_out),

      .rd_addr_a_i,
      .rd_data_a_o(rd_data_a_intg_o),

      .rd_addr_b_i,
      .rd_data_b_o(rd_data_b_intg_o),

      .we_err_o(spurious_we_err_o)
    );
  end

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) u_rf_ren_a_onehot_enc (
    .in_i  (rd_addr_a_i),
    .en_i  (rd_en_a_i),
    .out_o (expected_rd_en_a_onehot)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) u_rf_ren_b_onehot_enc (
    .in_i  (rd_addr_b_i),
    .en_i  (rd_en_b_i),
    .out_o (expected_rd_en_b_onehot)
  );

  prim_onehot_enc #(
    .OneHotWidth(NWdr)
  ) u_rf_we_onehot_enc (
    .in_i  (wr_addr_i),
    .en_i  (|wr_en_i),
    .out_o (expected_wr_en_onehot)
  );

  // SEC_CM: CTRL.REDUN
  assign rd_en_a_mismatch = expected_rd_en_a_onehot != rf_predec_bignum_i.rf_ren_a;
  assign rd_en_b_mismatch = expected_rd_en_b_onehot != rf_predec_bignum_i.rf_ren_b;
  assign wr_en_mismatch   = expected_wr_en_onehot   != rf_predec_bignum_i.rf_we;

  assign predec_error_o = rd_en_a_mismatch | rd_en_b_mismatch | wr_en_mismatch;

  // New data can have its integrity from an external source or the integrity can be calculated here
  assign wr_data_intg_mux_out = wr_data_intg_sel_i ? wr_data_intg_i : wr_data_intg_calc;

  // SEC_CM: RF_BIGNUM.DATA_REG_SW.INTEGRITY
  // Separate integrity encode and decode per 32-bit integrity granule
  for (genvar i = 0; i < BaseWordsPerWLEN; ++i) begin : g_rf_intg_calc
    prim_secded_inv_39_32_enc u_wr_data_intg_enc (
      .data_i(wr_data_no_intg_i[i * 32 +: 32]),
      .data_o(wr_data_intg_calc[i * 39 +: 39])
    );

    // Integrity decoders used to detect errors only, corrections (`syndrome_o`/`d_o`) are ignored
    prim_secded_inv_39_32_dec u_rd_data_a_intg_dec (
      .data_i    (rd_data_a_intg_o[i * 39 +: 39]),
      .data_o    (),
      .syndrome_o(),
      .err_o     (rd_data_a_err[i*2 +: 2])
    );

    prim_secded_inv_39_32_dec u_rd_data_b_intg_dec (
      .data_i    (rd_data_b_intg_o[i * 39 +: 39]),
      .data_o    (),
      .syndrome_o(),
      .err_o     (rd_data_b_err[i*2 +: 2])
    );
  end

  logic intg_err_unbuf, intg_err_buf;
  
  //zdr ecc disable
  logic intg_err_unbuf_zdr;
  assign intg_err_unbuf_zdr = ((|rd_data_a_err) & rd_en_a_i) |
                          ((|rd_data_b_err) & rd_en_b_i);
  assign intg_err_unbuf = intg_err_unbuf_zdr & 1'b0;

  // This primitive is used to place a constraint for synthesis. It is required to
  // ensure that the signal name will be available in the synthesized netlist.
  prim_buf #(
    .Width(1)
  ) u_prim_buf (
    .in_i(intg_err_unbuf),
    .out_o(intg_err_buf)
  );

  assign intg_err_o = intg_err_buf;

  `ASSERT(BlankingBignumRegReadA_A,
          !rd_en_a_i |->  rd_data_a_intg_o == '0,
          clk_i, !rst_ni || predec_error_o || !wr_commit_i)

  `ASSERT(BlankingBignumRegReadB_A,
          !rd_en_b_i |->  rd_data_b_intg_o == '0,
          clk_i, !rst_ni || predec_error_o || !wr_commit_i)

  // Make sure we're not outputting X. This indicates that something went wrong during the initial
  // secure wipe.
  `ASSERT(OtbnRfBignumRdAKnown, rd_en_a_i && !rd_en_a_mismatch |-> !$isunknown(rd_data_a_intg_o))
  `ASSERT(OtbnRfBignumRdBKnown, rd_en_b_i && !rd_en_b_mismatch |-> !$isunknown(rd_data_b_intg_o))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * 39b General Purpose Register File (GPRs)
 *
 * 39b to support 32b register with 7b integrity. Integrity generation/checking implemented in
 * wrapping otbn_rf_base module
 *
 * Features:
 * - 2 read ports
 * - 1 write port
 */
module otbn_rf_base_ff
  import otbn_pkg::*;
#(
  parameter logic [BaseIntgWidth-1:0] WordZeroVal = '0
) (
  input logic                     clk_i,
  input logic                     rst_ni,

  input logic  [4:0]               wr_addr_i,
  input logic                      wr_en_i,
  input logic  [BaseIntgWidth-1:0] wr_data_i,

  input  logic [4:0]               rd_addr_a_i,
  output logic [BaseIntgWidth-1:0] rd_data_a_o,

  input  logic [4:0]               rd_addr_b_i,
  output logic [BaseIntgWidth-1:0] rd_data_b_o,

  // Indicates whether a spurious WE has been seen in the last cycle.
  output logic                     we_err_o
);

  logic [BaseIntgWidth-1:0] rf_reg [NGpr];
  logic [31:0] we_onehot;

  for (genvar i = 0; i < NGpr; i++) begin : g_we_onehot
    assign we_onehot[i] = (wr_addr_i == i) && wr_en_i;
  end

  // No flops for register 0 as it's hard-wired to 0
  assign rf_reg[0] = WordZeroVal;

  // No flops for register 1 as it's call stack and handled in a different module.
  assign rf_reg[1] = WordZeroVal;

  // Generate flops for register 1 - NGpr
  for (genvar i = 2; i < NGpr; i++) begin : g_rf_flops
    logic [BaseIntgWidth-1:0] rf_reg_q;

    always_ff @(posedge clk_i) begin
      if(we_onehot[i]) begin
        rf_reg_q <= wr_data_i;
      end
    end

    assign rf_reg[i] = rf_reg_q;
  end

  assign rd_data_a_o = rf_reg[rd_addr_a_i];
  assign rd_data_b_o = rf_reg[rd_addr_b_i];

  // Buffer the decoded write enable bits so that the checker
  // is not optimized into the address decoding logic.
  logic [31:0] we_onehot_buf;
  prim_buf #(
    .Width(32)
  ) u_prim_buf (
    .in_i(we_onehot),
    .out_o(we_onehot_buf)
  );

  // SEC_CM: RF_BASE.DATA_REG_SW.GLITCH_DETECT
  // This checks for spurious WE strobes on the regfile.
  logic we_err;
  prim_onehot_check #(
    .AddrWidth(5),
    .AddrCheck(1),
    .EnableCheck(1)
  ) u_prim_onehot_check (
    .clk_i,
    .rst_ni,
    .oh_i(we_onehot_buf),
    .addr_i(wr_addr_i),
    .en_i(wr_en_i),
    .err_o(we_err)
  );

  // We need to register this to avoid timing loops.
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_err
    if (!rst_ni) begin
      we_err_o <= '0;
    end else begin
      we_err_o <= we_err;
    end
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * ExtWLEN (312b) Wide Register File (WDRs)
 *
 * ExtWLEN allows bits to provide integrity checking to WLEN words on a 32-bit granule. Integrity
 * generation/checking implemented in wrapping otbn_rf_bignum module
 *
 * Features:
 * - 2 read ports
 * - 1 write port
 * - Half (WLEN) word write enables
 */
module otbn_rf_bignum_ff
  import otbn_pkg::*;
(
  input  logic             clk_i,
  input  logic             rst_ni,

  input  logic [WdrAw-1:0]   wr_addr_i,
  input  logic [1:0]         wr_en_i,
  input  logic [ExtWLEN-1:0] wr_data_i,

  input  logic [WdrAw-1:0]   rd_addr_a_i,
  output logic [ExtWLEN-1:0] rd_data_a_o,

  input  logic [WdrAw-1:0]   rd_addr_b_i,
  output logic [ExtWLEN-1:0] rd_data_b_o,

  // Indicates whether a spurious WE has been seen in the last cycle.
  output logic               we_err_o,

  input  rf_predec_bignum_t  rf_predec_bignum_i
);
  logic [ExtWLEN-1:0] rf [NWdr];
  logic [1:0]         we_onehot [NWdr];

  logic unused_addr;

  for (genvar i = 0; i < NWdr; i++) begin : g_rf
    logic [ExtWLEN-1:0] wr_data_blanked;
    assign we_onehot[i] = wr_en_i & {2{wr_addr_i == i}};

    // SEC_CM: DATA_REG_SW.SCA
    prim_blanker #(.Width(ExtWLEN)) u_wdata_blanker(
      .in_i (wr_data_i),
      .en_i (rf_predec_bignum_i.rf_we[i]),
      .out_o(wr_data_blanked)
    );

    // Split registers into halves for clear seperation for the enable terms
    always_ff @(posedge clk_i) begin
      if (rf_predec_bignum_i.rf_we[i] & we_onehot[i][0]) begin
        rf[i][0+:ExtWLEN/2] <= wr_data_blanked[0+:ExtWLEN/2];
      end
    end

    always_ff @(posedge clk_i) begin
      if (rf_predec_bignum_i.rf_we[i] & we_onehot[i][1]) begin
        rf[i][ExtWLEN/2+:ExtWLEN/2] <= wr_data_blanked[ExtWLEN/2+:ExtWLEN/2];
      end
    end

  `ASSERT(BlankingBignumRegWData_A, !(|we_onehot[i]) |-> wr_data_blanked inside {'0, 'x})
  end

  // SEC_CM: DATA_REG_SW.SCA
  prim_onehot_mux #(
    .Width(ExtWLEN),
    .Inputs(NWdr)
  ) u_rd_mux_a (
    .clk_i,
    .rst_ni,
    .in_i  (rf),
    .sel_i (rf_predec_bignum_i.rf_ren_a),
    .out_o (rd_data_a_o)
  );

  prim_onehot_mux  #(
    .Width(ExtWLEN),
    .Inputs(NWdr)
  ) u_rd_mux_b (
    .clk_i,
    .rst_ni,
    .in_i  (rf),
    .sel_i (rf_predec_bignum_i.rf_ren_b),
    .out_o (rd_data_b_o)
  );

  assign unused_addr = ^rd_addr_a_i ^ ^rd_addr_b_i ^ ^wr_addr_i;

  logic we_err, we_err_d;
  logic [1:0][NWdr-1:0] we_onehot_unbuf, we_onehot_buf;

  for (genvar k = 0; k < 2; k++) begin : g_check
    for (genvar i = 0; i < NWdr; i++) begin : g_reshape
      assign we_onehot_unbuf[k][i] = we_onehot[i][k];
    end
  end

  // Buffer the decoded write enable bits so that the checker
  // is not optimized into the address decoding logic.
  prim_buf #(
    .Width(2*NWdr)
  ) u_prim_buf (
    .in_i(we_onehot_unbuf),
    .out_o(we_onehot_buf)
  );

  // SEC_CM: RF_BIGNUM.DATA_REG_SW.GLITCH_DETECT
  // This checks for spurious WE strobes on the regfile.
  prim_onehot_check #(
    .AddrWidth(WdrAw),
    .OneHotWidth(NWdr),
    .AddrCheck(1),
    .EnableCheck(1)
  ) u_prim_onehot_check (
    .clk_i,
    .rst_ni,
    // OR the two register halves.
    .oh_i(we_onehot_buf[0] | we_onehot_buf[1]),
    .addr_i(wr_addr_i),
    .en_i(|wr_en_i),
    .err_o(we_err)
  );

  assign we_err_d = we_err | we_err_o;

  prim_flop #(
    .Width(1),
    .ResetValue('0)
  ) u_we_err_flop (
    .clk_i,
    .rst_ni,

    .d_i(we_err_d),
    .q_o(we_err_o)
  );

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * 39b General Purpose Register File (GPRs)
 *
 * 39b to support 32b register with 7b integrity. Integrity generation/checking implemented in
 * wrapping otbn_rf_base module
 *
 * Features:
 * - 2 read ports
 * - 1 write port
 *
 * Register 0 is fixed to 0.
 *
 * This register file is designed to make FPGA synthesis tools infer RAM primitives. For Xilinx
 * FPGA architectures, it will produce RAM32M primitives. Other vendors have not yet been tested.
 */
module otbn_rf_base_fpga
  import otbn_pkg::*;
#(
  parameter logic [BaseIntgWidth-1:0] WordZeroVal = '0
) (
  input logic                     clk_i,
  input logic                     rst_ni,

  input logic  [4:0]               wr_addr_i,
  input logic                      wr_en_i,
  input logic  [BaseIntgWidth-1:0] wr_data_i,

  input  logic [4:0]               rd_addr_a_i,
  output logic [BaseIntgWidth-1:0] rd_data_a_o,

  input  logic [4:0]               rd_addr_b_i,
  output logic [BaseIntgWidth-1:0] rd_data_b_o,

  // Indicates whether a spurious WE has been seen in the last cycle.
  output logic                     we_err_o
);
  logic [BaseIntgWidth-1:0] rf_reg [NGpr];
  logic                    wr_en;

  // The reset is not used in this register file version.
  logic unused_rst_ni;
  assign unused_rst_ni = rst_ni;

  // No write-enable for register 0 as writes to it are ignored.
  assign wr_en = (wr_addr_i == '0) ? 1'b0 : wr_en_i;

  // Sync write
  // Note that the SystemVerilog LRM requires variables on the LHS of assignments within
  // "always_ff" to not be written to by any other process. However, to enable the initialization
  // of the inferred RAM32M primitives with non-zero values, below "initial" procedure is needed.
  // Therefore, we use "always" instead of the generally preferred "always_ff" for the synchronous
  // write procedure.
  always @(posedge clk_i) begin : g_rf_reg
    if (wr_en == 1'b1) begin
      rf_reg[wr_addr_i] <= wr_data_i;
    end
  end

  // Make sure we initialize the BRAM with the correct register reset value.
  initial begin
    for (int k = 0; k < NGpr; k++) begin
      rf_reg[k] = WordZeroVal;
    end
  end

  // Async read
  assign rd_data_a_o = (rd_addr_a_i == '0) ? WordZeroVal : rf_reg[rd_addr_a_i];
  assign rd_data_b_o = (rd_addr_b_i == '0) ? WordZeroVal : rf_reg[rd_addr_b_i];

  // SEC_CM: RF_BASE.DATA_REG_SW.GLITCH_DETECT
  // This checks for spurious WE strobes on the regfile.
  // Since the FPGA uses a memory macro, there is only one write-enable strobe to check.
  logic we_err;
  assign we_err = wr_en && !wr_en_i;

  // We need to register this to avoid timing loops.
  always_ff @(posedge clk_i or negedge rst_ni) begin : p_err
    if (!rst_ni) begin
      we_err_o <= '0;
    end else begin
      we_err_o <= we_err;
    end
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * ExtWLEN (312b) Wide Register File (WDRs)
 *
 * ExtWLEN allows bits to provide integrity checking to WLEN words on a 32-bit granule. Integrity
 * generation/checking implemented in wrapping otbn_rf_bignum module
 *
 * Features:
 * - 2 read ports
 * - 1 write port
 * - Half (WLEN) word write enables
 *
 * This register file is designed to make FPGA synthesis tools infer RAM primitives. For Xilinx
 * FPGA architectures, it will produce RAM32M primitives. Other vendors have not yet been tested.
 */
module otbn_rf_bignum_fpga
  import otbn_pkg::*;
#(
  parameter logic [BaseIntgWidth-1:0] WordZeroVal = '0
) (
  input  logic             clk_i,
  input  logic             rst_ni,

  input  logic [WdrAw-1:0]   wr_addr_i,
  input  logic [1:0]         wr_en_i,
  input  logic [ExtWLEN-1:0] wr_data_i,

  input  logic [WdrAw-1:0]   rd_addr_a_i,
  output logic [ExtWLEN-1:0] rd_data_a_o,

  input  logic [WdrAw-1:0]   rd_addr_b_i,
  output logic [ExtWLEN-1:0] rd_data_b_o,

  // Indicates whether a spurious WE has been seen in the last cycle.
  output logic               we_err_o
);


  // The reset is not used in this register file version.
  logic unused_rst_ni;
  assign unused_rst_ni = rst_ni;

  // This is only used for backdoor access in simulations.
  logic [ExtWLEN-1:0] rf [NWdr];
  logic [ExtWLEN-1:0] unused_rf [NWdr];
  assign unused_rf = rf;

  // Split registers into individual 39bit wide memories - otherwise the tool fails to properly
  // implement the non-zero memory intialization assignment in the initial block. Further, the
  // regfile is split into two sets of memories for clear separation of the enable terms.
  for (genvar i = 0; i < BaseWordsPerWLEN; i++) begin : gen_rf
    logic [BaseIntgWidth-1:0] rf_local [NWdr];
    // Sync write
    // Note that the SystemVerilog LRM requires variables on the LHS of assignments within
    // "always_ff" to not be written to by any other process. However, to enable the initialization
    // of the inferred RAM32M primitives with non-zero values, below "initial" procedure is needed.
    // Therefore, we use "always" instead of the generally preferred "always_ff" for the synchronous
    // write procedure.
    always @(posedge clk_i) begin
      if (wr_en_i[i/(BaseWordsPerWLEN/2)] == 1'b1) begin
        rf_local[wr_addr_i] <= wr_data_i[i*BaseIntgWidth+:BaseIntgWidth];
      end
    end

    // Make sure we initialize the BRAM with the correct register reset value.
    initial begin
      for (int k = 0; k < NWdr; k++) begin
        rf_local[k] = WordZeroVal;
      end
    end

    // Async read
    assign rd_data_a_o[i*BaseIntgWidth+:BaseIntgWidth] = rf_local[rd_addr_a_i];
    assign rd_data_b_o[i*BaseIntgWidth+:BaseIntgWidth] = rf_local[rd_addr_b_i];

    // SEC_CM: RF_BASE.DATA_REG_SW.GLITCH_DETECT
    // There is nothing to check here since the decoding happens inside the inferred
    // memory block.
    assign we_err_o = 1'b0;

  // This is only used for backdoor access in simulations.
`ifdef VERILATOR
  `define INC_BACKDOOR_LOAD
`elsif SIMULATION
  `define INC_BACKDOOR_LOAD
`endif
`ifdef INC_BACKDOOR_LOAD
    for (genvar k = 0; k < NWdr; k++) begin : gen_sim
      assign rf[k][i*BaseIntgWidth+:BaseIntgWidth] = rf_local[k];
    end
`undef INC_BACKDOOR_LOAD
`endif
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN Load-Store Unit
 *
 * Read and write data from/to the data memory (DMEM). Used by the base and the BN instruction
 * subset; loads and stores are hence either 32b or WLEN bit wide.
 *
 * The data memory interface makes the following assumptions:
 * - All requests are answered in the next cycle; the LSU must have exclusive access to the memory.
 * - The write mask supports aligned 32b write accesses.
 */
module otbn_lsu
  import otbn_pkg::*;
#(
  parameter int DmemSizeByte = 4096,

  localparam int DmemAddrWidth = prim_util_pkg::vbits(DmemSizeByte)
) (
  input logic clk_i,
  input logic rst_ni,

  // Data memory (DMEM) interface
  output logic                        dmem_req_o,
  output logic                        dmem_write_o,
  output logic [DmemAddrWidth-1:0]    dmem_addr_o,
  output logic [ExtWLEN-1:0]          dmem_wdata_o,
  output logic [ExtWLEN-1:0]          dmem_wmask_o,
  output logic [BaseWordsPerWLEN-1:0] dmem_rmask_o,
  input  logic [ExtWLEN-1:0]          dmem_rdata_i,
  input  logic                        dmem_rvalid_i,
  input  logic                        dmem_rerror_i,

  input  logic                     lsu_load_req_i,
  input  logic                     lsu_store_req_i,
  input  insn_subset_e             lsu_req_subset_i,
  input  logic [DmemAddrWidth-1:0] lsu_addr_i,

  input  logic [BaseIntgWidth-1:0] lsu_base_wdata_i,
  input  logic [ExtWLEN-1:0]       lsu_bignum_wdata_i,

  output logic [BaseIntgWidth-1:0] lsu_base_rdata_o,
  output logic [ExtWLEN-1:0]       lsu_bignum_rdata_o,
  output logic                     lsu_rdata_err_o
);
  localparam int BaseWordsPerWLen = WLEN / 32;
  localparam int BaseWordAddrW = prim_util_pkg::vbits(WLEN / 8);

  // Produce a WLEN bit mask for 32-bit writes given the 32-bit word write address. This doesn't
  // propagate X so a separate assertion must be used to check the input isn't X when a valid output
  // is desired.
  function automatic logic [ExtWLEN-1:0] wmask_from_word_addr(logic [BaseWordAddrW-1:2] addr);
    logic [ExtWLEN-1:0] mask;

    mask = '0;

    // Use of logic == int comparison in this loop works as BaseWordsPerWLen is a constant, so the
    // loop can be unrolled. Due to the use of '==' any X or Z in addr will result in an X result
    // for the comparison (so mask will remain 0).
    for (int i = 0; i < BaseWordsPerWLen; i++) begin
      if (addr == i) begin
        mask[i*BaseIntgWidth+:BaseIntgWidth] = '1;
      end
    end

    return mask;
  endfunction

  function automatic logic [BaseWordsPerWLEN-1:0]
      rmask_from_word_addr(logic [BaseWordAddrW-1:2] addr);

    logic [BaseWordsPerWLEN-1:0] mask;

    mask = '0;

    for (int i = 0; i < BaseWordsPerWLen; i++) begin
      if (addr == i) begin
        mask[i] = 1'b1;
      end
    end

    return mask;
  endfunction

  logic [BaseWordAddrW-1:2] lsu_word_select;
  logic                     lsu_word_select_en;

  assign dmem_req_o   = lsu_load_req_i | lsu_store_req_i;
  assign dmem_write_o = lsu_store_req_i;
  assign dmem_addr_o  = lsu_addr_i;

  // For base 32-bit writes replicate write data across dmem_wdata. dmem_wmask will be set
  // appropriately so only the target word is written.
  assign dmem_wdata_o = lsu_req_subset_i == InsnSubsetBase ?
    {BaseWordsPerWLen{lsu_base_wdata_i}} : lsu_bignum_wdata_i;

  assign dmem_wmask_o = lsu_req_subset_i == InsnSubsetBase ?
    wmask_from_word_addr(lsu_addr_i[BaseWordAddrW-1:2]) : {ExtWLEN{1'b1}};

  assign dmem_rmask_o = lsu_req_subset_i == InsnSubsetBase ?
    rmask_from_word_addr(lsu_addr_i[BaseWordAddrW-1:2]) : {BaseWordsPerWLEN{1'b1}};

  // Store a portion of the address to select a 32-bit word from the WLEN load data when it returns
  // the cycle following the request.
  assign lsu_word_select_en = lsu_load_req_i & (lsu_req_subset_i == InsnSubsetBase);

  always_ff @(posedge clk_i) begin
    if (lsu_word_select_en) begin
      lsu_word_select <= lsu_addr_i[BaseWordAddrW-1:2];
    end
  end

  // From the WLEN word read from DMem select out a 32-bit word for base instructions.
  for (genvar i_bit = 0; i_bit < BaseIntgWidth; i_bit++) begin : g_base_rdata
    logic [BaseWordsPerWLen-1:0] bit_mux;

    for (genvar j_word = 0; j_word < BaseWordsPerWLen; j_word++) begin : g_bit_mux
      assign bit_mux[j_word] =
        (lsu_word_select == j_word) & dmem_rdata_i[i_bit + j_word * BaseIntgWidth];
    end

    assign lsu_base_rdata_o[i_bit] = |bit_mux;
  end

  `ASSERT_KNOWN_IF(LsuAddrKnown, lsu_addr_i, lsu_load_req_i | lsu_store_req_i)

  `ASSERT(DMemRValidAfterReq, dmem_req_o & ~dmem_write_o |=> dmem_rvalid_i)

  assign lsu_bignum_rdata_o = dmem_rdata_i;
  assign lsu_rdata_err_o    = dmem_rvalid_i & dmem_rerror_i;

  // clk_i, rst_ni are only used by assertions
  logic unused_clk;
  logic unused_rst_n;

  assign unused_clk   = clk_i;
  assign unused_rst_n = rst_ni;
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN execute block for the base instruction subset
 *
 * This ALU supports the execution of all of OTBN's base instruction subset.
 */
module otbn_alu_base
  import otbn_pkg::*;
(
  // Block is combinatorial; clk/rst are for assertions only.
  input logic clk_i,
  input logic rst_ni,

  input alu_base_operation_t  operation_i,
  input alu_base_comparison_t comparison_i,

  output logic [31:0] operation_result_o,
  output logic        comparison_result_o
);

  logic [32:0] adder_op_a, adder_op_b;
  logic        adder_op_b_negate;
  logic [32:0] adder_result;

  logic [31:0] and_result;
  logic [31:0] or_result;
  logic [31:0] xor_result;
  logic [31:0] not_result;

  logic        is_equal;

  ///////////
  // Adder //
  ///////////

  // Adder takes in 33-bit operands. The addition of the input operands occurs on bits [32:1],
  // setting addr_op_b_negate will cause a carry-in into bit 1. Combined with an inversion of
  // operation_i.operand_b this gives a two's-complement negation (~b + 1)

  assign adder_op_b_negate = operation_i.op == AluOpBaseSub;

  assign adder_op_a = {operation_i.operand_a, 1'b1};
  assign adder_op_b = adder_op_b_negate ? {~operation_i.operand_b, 1'b1} :
                                          { operation_i.operand_b, 1'b0};

  assign adder_result = adder_op_a + adder_op_b;

  //////////////////////////
  // Bit-wise logical ops //
  //////////////////////////

  assign and_result = operation_i.operand_a & operation_i.operand_b;
  assign or_result  = operation_i.operand_a | operation_i.operand_b;
  assign xor_result = operation_i.operand_a ^ operation_i.operand_b;
  assign not_result = ~operation_i.operand_a;

  /////////////
  // Shifter //
  /////////////

  logic [32:0] shift_in;
  logic [ 4:0] shift_amt;
  logic [31:0] operand_a_reverse;
  logic [32:0] shift_out;
  logic [31:0] shift_out_reverse;

  for (genvar i = 0; i < 32; i++) begin : g_shifter_reverses
    assign operand_a_reverse[i] = operation_i.operand_a[31-i];
    assign shift_out_reverse[i] = shift_out[31-i];
  end

  assign shift_amt = operation_i.operand_b[4:0];
  // Shifter performs right arithmetic 33-bit shifts. Force top bit to 0 to get logical shifting
  // otherwise replicate top bit of shift_in. Left shifts performed by reversing the input and
  // output.
  assign shift_in[31:0] = (operation_i.op == AluOpBaseSll) ? operand_a_reverse :
                                                             operation_i.operand_a;
  assign shift_in[32] = (operation_i.op == AluOpBaseSra) ? operation_i.operand_a[31] : 1'b0;

  logic signed [32:0] shift_in_signed;
  assign shift_in_signed = signed'(shift_in);
  assign shift_out = unsigned'(shift_in_signed >>> shift_amt);

  ////////////////
  // Output Mux //
  ////////////////

  always_comb begin
    operation_result_o = adder_result[32:1];

    unique case (operation_i.op)
      AluOpBaseAnd: operation_result_o = and_result;
      AluOpBaseOr:  operation_result_o = or_result;
      AluOpBaseXor: operation_result_o = xor_result;
      AluOpBaseNot: operation_result_o = not_result;
      AluOpBaseSra: operation_result_o = shift_out[31:0];
      AluOpBaseSrl: operation_result_o = shift_out[31:0];
      AluOpBaseSll: operation_result_o = shift_out_reverse;
      default: ;
    endcase
  end

  /////////////////
  // Comparisons //
  /////////////////

  // Dedicated comparator to deal with branches. As only Equal/Not-Equal is required no need to use
  // the adder (which frees it to compute the branch target in the same cycle). No point in using
  // existing XOR logic as area added from extra mux to choose xor operands negates area saving from
  // avoiding an dedicated comparator.
  assign is_equal = comparison_i.operand_a == comparison_i.operand_b;

  assign comparison_result_o = (comparison_i.op == ComparisonOpBaseEq) ? is_equal : ~is_equal;

  // The bottom bit of adder_result is discarded. It simply corresponds to the carry in used to
  // produce twos complement subtraction from an addition.
  logic unused_adder_result_bit;

  // The top bit of shift_out is discarded. shift_in contains an extra bit to deal with sign
  // extension which isn't needed in the shift_out result.
  logic unused_shift_out_result_bit;
  assign unused_shift_out_result_bit = shift_out[32];

  assign unused_adder_result_bit = adder_result[0];

  // clk_i, rst_ni are only used by assertions
  logic unused_clk;
  logic unused_rst_n;

  assign unused_clk   = clk_i;
  assign unused_rst_n = rst_ni;
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN alu block for the bignum instruction subset
 *
 * This ALU supports all of the 'plain' arithmetic and logic bignum instructions, BN.MULQACC is
 * implemented in a separate block.
 *
 * One barrel shifter and two adders (X and Y) are implemented along with the logic operators
 * (AND,OR,XOR,NOT).
 *
 * The adders have 256-bit operands with a carry_in and optional invert on the second operand. This
 * can be used to implement subtraction (a - b == a + ~b + 1). BN.SUBB/BN.ADDC are implemented by
 * feeding in the carry flag as carry in rather than a fixed 0 or 1.
 *
 * The shifter takes a 512-bit input (to implement BN.RSHI, concatenate and right shift) and shifts
 * right by up to 256-bits. The lower (256-bit) half of the input and output can be reversed to
 * allow left shift implementation.  There is no concatenate and left shift instruction so reversing
 * isn't required over the full width.
 *
 * The dataflow between the adders and shifter is in the diagram below. This arrangement allows the
 * implementation of the pseudo-mod (BN.ADDM/BN.SUBM) instructions in a single cycle whilst
 * minimising the critical path. The pseudo-mod instructions do not have a shifted input so X can
 * compute the initial add/sub and Y computes the pseudo-mod result. For all other add/sub
 * operations Y computes the operation with one of the inputs supplied by the shifter and the other
 * from operand_a.
 *
 * Both adder X and the shifter get supplied with operand_a and operand_b from the operation_i
 * input. In addition the shifter gets a shift amount (shift_amt) and can use 0 instead of
 * operand_a. The shifter concatenates operand_a (or 0) and operand_b together before shifting with
 * operand_a in the upper (256-bit) half {operand_a/0, operand_b}. This allows the shifter to pass
 * through operand_b simply by not performing a shift.
 *
 * Blanking is employed on the ALU data paths. This holds unused data paths to 0 to reduce side
 * channel leakage. The lower-case 'b' on the digram below indicates points in the data path that
 * get blanked. Note that Adder X is never used in isolation, it is always combined with Adder Y so
 * there is no need for blanking between Adder X and Adder Y.
 *
 *      A       B       A   B
 *      |       |       |   |
 *      b       b       b   b   shift_amt
 *      |       |       |   |   |
 *    +-----------+   +-----------+
 *    |  Adder X  |   |  Shifter  |
 *    +-----------+   +-----------+
 *          |               |
 *          |----+     +----|
 *          |    |     |    |
 *      X result |     | Shifter result
 *               |     |
 *             A |     |
 *             | |     |     +-----------+
 *             b |     b +---|  MOD WSR  |
 *             | |     | |   +-----------+
 *           \-----/ \-----/
 *            \---/   \---/
 *              |       |
 *              |       |
 *            +-----------+
 *            |  Adder Y  |
 *            +-----------+
 *                  |
 *              Y result
 */


module otbn_alu_bignum
  import otbn_pkg::*;
(
  input logic clk_i,
  input logic rst_ni,

  input  alu_bignum_operation_t operation_i,
  input  logic                  operation_valid_i,
  input  logic                  operation_commit_i, // used for SVAs only
  output logic [WLEN-1:0]       operation_result_o,
  output logic                  selection_flag_o,

  input  alu_predec_bignum_t  alu_predec_bignum_i,
  input  ispr_predec_bignum_t ispr_predec_bignum_i,

  input  ispr_e                       ispr_addr_i,
  input  logic [31:0]                 ispr_base_wdata_i,
  input  logic [BaseWordsPerWLEN-1:0] ispr_base_wr_en_i,
  input  logic [ExtWLEN-1:0]          ispr_bignum_wdata_intg_i,
  input  logic                        ispr_bignum_wr_en_i,
  input  logic [NFlagGroups-1:0]      ispr_flags_wr_i,
  input  logic                        ispr_wr_commit_i,
  input  logic                        ispr_init_i,
  output logic [ExtWLEN-1:0]          ispr_rdata_intg_o,
  input  logic                        ispr_rd_en_i,

  input  logic [ExtWLEN-1:0]          ispr_acc_intg_i,
  output logic [ExtWLEN-1:0]          ispr_acc_wr_data_intg_o,
  output logic                        ispr_acc_wr_en_o,

  output logic                        reg_intg_violation_err_o,

  input logic                         sec_wipe_mod_urnd_i,

  input  flags_t                      mac_operation_flags_i,
  input  flags_t                      mac_operation_flags_en_i,

  input  logic [WLEN-1:0]             rnd_data_i,
  input  logic [WLEN-1:0]             urnd_data_i,

  input  logic [1:0][SideloadKeyWidth-1:0] sideload_key_shares_i,

  output logic alu_predec_error_o,
  output logic ispr_predec_error_o
);

  logic [WLEN+1:0] adder_y_res;
  logic [WLEN-1:0] logical_res;

  ///////////
  // ISPRs //
  ///////////

  flags_t                              flags_d [NFlagGroups];
  flags_t                              flags_q [NFlagGroups];
  logic   [NFlagGroups*FlagsWidth-1:0] flags_flattened;
  flags_t                              selected_flags;
  flags_t                              adder_update_flags;
  logic                                adder_update_flags_en_raw;
  flags_t                              logic_update_flags [NFlagGroups];
  logic                                logic_update_flags_en_raw;
  flags_t                              mac_update_flags [NFlagGroups];
  logic [NFlagGroups-1:0]              mac_update_z_flag_en_blanked;
  flags_t                              ispr_update_flags [NFlagGroups];

  logic [NIspr-1:0] expected_ispr_rd_en_onehot;
  logic [NIspr-1:0] expected_ispr_wr_en_onehot;
  logic             ispr_wr_en;

  logic [NFlagGroups-1:0] expected_flag_group_sel;
  flags_t                 expected_flag_sel;
  logic [NFlagGroups-1:0] expected_flags_keep;
  logic [NFlagGroups-1:0] expected_flags_adder_update;
  logic [NFlagGroups-1:0] expected_flags_logic_update;
  logic [NFlagGroups-1:0] expected_flags_mac_update;
  logic [NFlagGroups-1:0] expected_flags_ispr_wr;

  /////////////////////
  // Flags Selection //
  /////////////////////

  always_comb begin
    expected_flag_group_sel = '0;
    expected_flag_group_sel[operation_i.flag_group] = 1'b1;
  end
  assign expected_flag_sel.C = operation_i.sel_flag == FlagC;
  assign expected_flag_sel.M = operation_i.sel_flag == FlagM;
  assign expected_flag_sel.L = operation_i.sel_flag == FlagL;
  assign expected_flag_sel.Z = operation_i.sel_flag == FlagZ;

  // SEC_CM: DATA_REG_SW.SCA
  prim_onehot_mux #(
    .Width(FlagsWidth),
    .Inputs(NFlagGroups)
  ) u_flags_q_mux (
    .clk_i,
    .rst_ni,
    .in_i  (flags_q),
    .sel_i (alu_predec_bignum_i.flag_group_sel),
    .out_o (selected_flags)
  );

  `ASSERT(BlankingSelectedFlags_A, expected_flag_group_sel == '0 |-> selected_flags == '0, clk_i,
    !rst_ni || alu_predec_error_o  || !operation_commit_i)


  logic                  flag_mux_in [FlagsWidth];
  logic [FlagsWidth-1:0] flag_mux_sel;
  assign flag_mux_in = '{selected_flags.C,
                         selected_flags.M,
                         selected_flags.L,
                         selected_flags.Z};
  assign flag_mux_sel = {alu_predec_bignum_i.flag_sel.Z,
                         alu_predec_bignum_i.flag_sel.L,
                         alu_predec_bignum_i.flag_sel.M,
                         alu_predec_bignum_i.flag_sel.C};

  // SEC_CM: DATA_REG_SW.SCA
  prim_onehot_mux #(
    .Width(1),
    .Inputs(FlagsWidth)
  ) u_flag_mux (
    .clk_i,
    .rst_ni,
    .in_i  (flag_mux_in),
    .sel_i (flag_mux_sel),
    .out_o (selection_flag_o)
  );

  `ASSERT(BlankingSelectionFlag_A, expected_flag_sel == '0 |-> selection_flag_o == '0, clk_i,
    !rst_ni || alu_predec_error_o  || !operation_commit_i)

  //////////////////
  // Flags Update //
  //////////////////

  // Note that the flag zeroing triggred by ispr_init_i and secure wipe is achieved by not
  // selecting any inputs in the one-hot muxes below. The instruction fetch/predecoder stage
  // is driving the selector inputs accordingly.

  always_comb begin
    expected_flags_adder_update = '0;
    expected_flags_logic_update = '0;
    expected_flags_mac_update   = '0;

    expected_flags_adder_update[operation_i.flag_group] = operation_i.alu_flag_en &
                                                          adder_update_flags_en_raw;
    expected_flags_logic_update[operation_i.flag_group] = operation_i.alu_flag_en &
                                                          logic_update_flags_en_raw;
    expected_flags_mac_update[operation_i.flag_group]   = operation_i.mac_flag_en;
  end
  assign expected_flags_ispr_wr = ispr_flags_wr_i;

  assign expected_flags_keep = ~(expected_flags_adder_update |
                                 expected_flags_logic_update |
                                 expected_flags_mac_update |
                                 expected_flags_ispr_wr);

  // Adder operations update all flags.
  assign adder_update_flags.C = (operation_i.op == AluOpBignumAdd ||
                                 operation_i.op == AluOpBignumAddc) ?  adder_y_res[WLEN+1] :
                                                                      ~adder_y_res[WLEN+1];
  assign adder_update_flags.M = adder_y_res[WLEN];
  assign adder_update_flags.L = adder_y_res[1];
  assign adder_update_flags.Z = ~|adder_y_res[WLEN:1];

  for (genvar i_fg = 0; i_fg < NFlagGroups; i_fg++) begin : g_update_flag_groups

    // Logical operations only update M, L and Z; C must remain at its old value.
    assign logic_update_flags[i_fg].C = flags_q[i_fg].C;
    assign logic_update_flags[i_fg].M = logical_res[WLEN-1];
    assign logic_update_flags[i_fg].L = logical_res[0];
    assign logic_update_flags[i_fg].Z = ~|logical_res;

    ///////////////
    // MAC Flags //
    ///////////////

    // MAC operations don't update C.
    assign mac_update_flags[i_fg].C = flags_q[i_fg].C;

    // Tie off unused signals.
    logic unused_mac_operation_flags;
    assign unused_mac_operation_flags = mac_operation_flags_i.C ^ mac_operation_flags_en_i.C;

    // MAC operations update M and L depending on the operation. The individual enable signals for
    // M and L are generated from flopped instruction bits with minimal logic. They are not data
    // dependent.
    assign mac_update_flags[i_fg].M = mac_operation_flags_en_i.M ?
                                      mac_operation_flags_i.M : flags_q[i_fg].M;
    assign mac_update_flags[i_fg].L = mac_operation_flags_en_i.L ?
                                      mac_operation_flags_i.L : flags_q[i_fg].L;

    // MAC operations update Z depending on the operation and data. For BN.MULQACC.SO, already the
    // enable signal is data dependent (it depends on the lower half of the accumulator result). As
    // a result the enable signal might change back and forth during instruction execution which may
    // lead to SCA leakage. There is nothing that can really be done to avoid this other than
    // pipelining the flag computation which has a peformance impact.
    //
    // By blanking the enable signal for the other flag group, we can at least avoid leakage related
    // to the other flag group, i.e., we give the programmer a way to control where the leakage
    // happens.
    // SEC_CM: DATA_REG_SW.SCA
    prim_blanker #(.Width(1)) u_mac_z_flag_en_blanker (
      .in_i (mac_operation_flags_en_i.Z),
      .en_i (alu_predec_bignum_i.flags_mac_update[i_fg]),
      .out_o(mac_update_z_flag_en_blanked[i_fg])
    );
    assign mac_update_flags[i_fg].Z = mac_update_z_flag_en_blanked[i_fg] ?
                                      mac_operation_flags_i.Z : flags_q[i_fg].Z;

    // For ISPR writes, we get the full write data from the base ALU and will select the relevant
    // parts using the blankers and one-hot muxes below.
    assign ispr_update_flags[i_fg] = ispr_base_wdata_i[i_fg*FlagsWidth+:FlagsWidth];
  end

  localparam int NFlagsSrcs = 5;
  for (genvar i_fg = 0; i_fg < NFlagGroups; i_fg++) begin : g_flag_groups

    flags_t                flags_d_mux_in [NFlagsSrcs];
    logic [NFlagsSrcs-1:0] flags_d_mux_sel;
    assign flags_d_mux_in = '{ispr_update_flags[i_fg],
                              mac_update_flags[i_fg],
                              logic_update_flags[i_fg],
                              adder_update_flags,
                              flags_q[i_fg]};
    assign flags_d_mux_sel = {alu_predec_bignum_i.flags_keep[i_fg],
                              alu_predec_bignum_i.flags_adder_update[i_fg],
                              alu_predec_bignum_i.flags_logic_update[i_fg],
                              alu_predec_bignum_i.flags_mac_update[i_fg],
                              alu_predec_bignum_i.flags_ispr_wr[i_fg]};

    // SEC_CM: DATA_REG_SW.SCA
    prim_onehot_mux #(
      .Width(FlagsWidth),
      .Inputs(NFlagsSrcs)
    ) u_flags_d_mux (
      .clk_i,
      .rst_ni,
      .in_i  (flags_d_mux_in),
      .sel_i (flags_d_mux_sel),
      .out_o (flags_d[i_fg])
    );

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        flags_q[i_fg] <= '{Z : 1'b0, L : 1'b0, M : 1'b0, C : 1'b0};
      end else begin
        flags_q[i_fg] <= flags_d[i_fg];
      end
    end

    assign flags_flattened[i_fg*FlagsWidth+:FlagsWidth] = flags_q[i_fg];
  end

  /////////
  // MOD //
  /////////

  logic [ExtWLEN-1:0]          mod_intg_q;
  logic [ExtWLEN-1:0]          mod_intg_d;
  logic [BaseWordsPerWLEN-1:0] mod_ispr_wr_en;
  logic [BaseWordsPerWLEN-1:0] mod_wr_en;

  logic [ExtWLEN-1:0] ispr_mod_bignum_wdata_intg_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(ExtWLEN)) u_ispr_mod_bignum_wdata_blanker (
    .in_i (ispr_bignum_wdata_intg_i),
    .en_i (ispr_predec_bignum_i.ispr_wr_en[IsprMod]),
    .out_o(ispr_mod_bignum_wdata_intg_blanked)
  );
  // If the blanker is enabled, the output will not carry the correct ECC bits.  This is not
  // a problem because a blanked value should never be written to the register.  If the blanked
  // value is written to the register nonetheless, an integrity error arises.

  logic [WLEN-1:0]                mod_no_intg_d;
  logic [WLEN-1:0]                mod_no_intg_q;
  logic [ExtWLEN-1:0]             mod_intg_calc;
  logic [2*BaseWordsPerWLEN-1:0]  mod_intg_err;
  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_mod_words
    prim_secded_inv_39_32_enc i_secded_enc (
      .data_i (mod_no_intg_d[i_word*32+:32]),
      .data_o (mod_intg_calc[i_word*39+:39])
    );
    prim_secded_inv_39_32_dec i_secded_dec (
      .data_i     (mod_intg_q[i_word*39+:39]),
      .data_o     (/* unused because we abort on any integrity error */),
      .syndrome_o (/* unused */),
      .err_o      (mod_intg_err[i_word*2+:2])
    );
    assign mod_no_intg_q[i_word*32+:32] = mod_intg_q[i_word*39+:32];

    always_ff @(posedge clk_i) begin
      if (mod_wr_en[i_word]) begin
        mod_intg_q[i_word*39+:39] <= mod_intg_d[i_word*39+:39];
      end
    end

    always_comb begin
      mod_no_intg_d[i_word*32+:32] = '0;
      unique case (1'b1)
        // Non-encoded inputs have to be encoded before writing to the register.
        sec_wipe_mod_urnd_i: begin
          // In a secure wipe, `urnd_data_i` is written to the register before the zero word.  The
          // ECC bits should not matter between the two writes, but nonetheless we encode
          // `urnd_data_i` so there is no spurious integrity error.
          mod_no_intg_d[i_word*32+:32] = urnd_data_i[i_word*32+:32];
          mod_intg_d[i_word*39+:39]  = mod_intg_calc[i_word*39+:39];
        end
        // Pre-encoded inputs can directly be written to the register.
        default: mod_intg_d[i_word*39+:39] = ispr_mod_bignum_wdata_intg_blanked[i_word*39+:39];
      endcase

      unique case (1'b1)
        ispr_init_i: mod_intg_d[i_word*39+:39] = EccZeroWord;
        ispr_base_wr_en_i[i_word]: begin
          mod_no_intg_d[i_word*32+:32] = ispr_base_wdata_i;
          mod_intg_d[i_word*39+:39] = mod_intg_calc[i_word*39+:39];
        end
        default: ;
      endcase
    end

    `ASSERT(ModWrSelOneHot, $onehot0({ispr_init_i, ispr_base_wr_en_i[i_word]}))

    assign mod_ispr_wr_en[i_word] = (ispr_addr_i == IsprMod)                          &
                                    (ispr_base_wr_en_i[i_word] | ispr_bignum_wr_en_i) &
                                    ispr_wr_commit_i;

    assign mod_wr_en[i_word] = ispr_init_i            |
                               mod_ispr_wr_en[i_word] |
                               sec_wipe_mod_urnd_i;
  end

  /////////
  // ACC //
  /////////

  assign ispr_acc_wr_en_o   =
    ((ispr_addr_i == IsprAcc) & ispr_bignum_wr_en_i & ispr_wr_commit_i) | ispr_init_i;


  logic [ExtWLEN-1:0] ispr_acc_bignum_wdata_intg_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(ExtWLEN)) u_ispr_acc_bignum_wdata_intg_blanker (
    .in_i (ispr_bignum_wdata_intg_i),
    .en_i (ispr_predec_bignum_i.ispr_wr_en[IsprAcc]),
    .out_o(ispr_acc_bignum_wdata_intg_blanked)
  );
  // If the blanker is enabled, the output will not carry the correct ECC bits.  This is not
  // a problem because a blanked value should never be used.  If the blanked value is used
  // nonetheless, an integrity error arises.

  assign ispr_acc_wr_data_intg_o = ispr_init_i ? EccWideZeroWord
                                               : ispr_acc_bignum_wdata_intg_blanked;

  // ISPR read data is muxed out in two stages:
  // 1. Select amongst the ISPRs that have no integrity bits. The output has integrity calculated
  //    for it.
  // 2. Select between the ISPRs that have integrity bits and the result of the first stage.

  // Number of ISPRs that have integrity protection
  localparam int NIntgIspr = 2;
  // IDs fpr ISPRs with integrity
  localparam int IsprModIntg = 0;
  localparam int IsprAccIntg = 1;
  // ID representing all ISPRs with no integrity
  localparam int IsprNoIntg = 2;

  logic [NIntgIspr:0] ispr_rdata_intg_mux_sel;
  logic [ExtWLEN-1:0] ispr_rdata_intg_mux_in    [NIntgIspr+1];
  logic [WLEN-1:0]    ispr_rdata_no_intg_mux_in [NIspr];

  // First stage
  // MOD and ACC supply their own integrity so these values are unused
  assign ispr_rdata_no_intg_mux_in[IsprMod] = 0;
  assign ispr_rdata_no_intg_mux_in[IsprAcc] = 0;

  assign ispr_rdata_no_intg_mux_in[IsprRnd]    = rnd_data_i;
  assign ispr_rdata_no_intg_mux_in[IsprUrnd]   = urnd_data_i;
  assign ispr_rdata_no_intg_mux_in[IsprFlags]  = {{(WLEN - (NFlagGroups * FlagsWidth)){1'b0}},
                                                 flags_flattened};
  // SEC_CM: KEY.SIDELOAD
  assign ispr_rdata_no_intg_mux_in[IsprKeyS0L] = sideload_key_shares_i[0][255:0];
  assign ispr_rdata_no_intg_mux_in[IsprKeyS0H] = {{(WLEN - (SideloadKeyWidth - 256)){1'b0}},
                                                  sideload_key_shares_i[0][SideloadKeyWidth-1:256]};
  assign ispr_rdata_no_intg_mux_in[IsprKeyS1L] = sideload_key_shares_i[1][255:0];
  assign ispr_rdata_no_intg_mux_in[IsprKeyS1H] = {{(WLEN - (SideloadKeyWidth - 256)){1'b0}},
                                                  sideload_key_shares_i[1][SideloadKeyWidth-1:256]};

  logic [WLEN-1:0]    ispr_rdata_no_intg;
  logic [ExtWLEN-1:0] ispr_rdata_intg_calc;

  // SEC_CM: DATA_REG_SW.SCA
  prim_onehot_mux #(
    .Width  (WLEN),
    .Inputs (NIspr)
  ) u_ispr_rdata_no_intg_mux (
    .clk_i,
    .rst_ni,
    .in_i  (ispr_rdata_no_intg_mux_in),
    .sel_i (ispr_predec_bignum_i.ispr_rd_en),
    .out_o (ispr_rdata_no_intg)
  );

  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_rdata_enc
    prim_secded_inv_39_32_enc i_secded_enc (
      .data_i(ispr_rdata_no_intg[i_word * 32 +: 32]),
      .data_o(ispr_rdata_intg_calc[i_word * 39 +: 39])
    );
  end

  // Second stage
  assign ispr_rdata_intg_mux_in[IsprModIntg] = mod_intg_q;
  assign ispr_rdata_intg_mux_in[IsprAccIntg] = ispr_acc_intg_i;
  assign ispr_rdata_intg_mux_in[IsprNoIntg]  = ispr_rdata_intg_calc;

  assign ispr_rdata_intg_mux_sel[IsprModIntg] = ispr_predec_bignum_i.ispr_rd_en[IsprMod];
  assign ispr_rdata_intg_mux_sel[IsprAccIntg] = ispr_predec_bignum_i.ispr_rd_en[IsprAcc];

  assign ispr_rdata_intg_mux_sel[IsprNoIntg]  =
    |{ispr_predec_bignum_i.ispr_rd_en[IsprKeyS1H:IsprKeyS0L],
      ispr_predec_bignum_i.ispr_rd_en[IsprUrnd],
      ispr_predec_bignum_i.ispr_rd_en[IsprFlags],
      ispr_predec_bignum_i.ispr_rd_en[IsprRnd]};

  // If we're reading from an ISPR we must be using the ispr_rdata_intg_mux
  `ASSERT(IsprRDataIntgMuxSelIfIsprRd_A,
    |ispr_predec_bignum_i.ispr_rd_en |-> |ispr_rdata_intg_mux_sel)

  // If we're reading from MOD or ACC we must not take the read data from the calculated integrity
  // path
  `ASSERT(IsprModMustTakeIntg_A,
    ispr_predec_bignum_i.ispr_rd_en[IsprMod] |-> !ispr_rdata_intg_mux_sel[IsprNoIntg])

  `ASSERT(IsprAccMustTakeIntg_A,
    ispr_predec_bignum_i.ispr_rd_en[IsprAcc] |-> !ispr_rdata_intg_mux_sel[IsprNoIntg])


  prim_onehot_mux #(
    .Width  (ExtWLEN),
    .Inputs (NIntgIspr+1)
  ) u_ispr_rdata_intg_mux (
    .clk_i,
    .rst_ni,
    .in_i  (ispr_rdata_intg_mux_in),
    .sel_i (ispr_rdata_intg_mux_sel),
    .out_o (ispr_rdata_intg_o)
  );

  prim_onehot_enc #(
    .OneHotWidth (NIspr)
  ) u_expected_ispr_rd_en_enc (
    .in_i(ispr_addr_i),
    .en_i (ispr_rd_en_i),
    .out_o (expected_ispr_rd_en_onehot)
  );

  assign ispr_wr_en = |{ispr_bignum_wr_en_i, ispr_base_wr_en_i};

  prim_onehot_enc #(
    .OneHotWidth (NIspr)
  ) u_expected_ispr_wr_en_enc (
    .in_i(ispr_addr_i),
    .en_i (ispr_wr_en),
    .out_o (expected_ispr_wr_en_onehot)
  );

  // SEC_CM: CTRL.REDUN
  assign ispr_predec_error_o =
    |{expected_ispr_rd_en_onehot != ispr_predec_bignum_i.ispr_rd_en,
      expected_ispr_wr_en_onehot != ispr_predec_bignum_i.ispr_wr_en};

  /////////////
  // Shifter //
  /////////////

  logic [WLEN-1:0]   shifter_in_upper, shifter_in_lower, shifter_in_lower_reverse;
  logic [WLEN*2-1:0] shifter_in;
  logic [WLEN*2-1:0] shifter_out;
  logic [WLEN-1:0]   shifter_out_lower_reverse, shifter_res, unused_shifter_out_upper;
  logic [WLEN-1:0]   shifter_operand_a_blanked;
  logic [WLEN-1:0]   shifter_operand_b_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_shifter_operand_a_blanker (
    .in_i (operation_i.operand_a),
    .en_i (alu_predec_bignum_i.shifter_a_en),
    .out_o(shifter_operand_a_blanked)
  );

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_shifter_operand_b_blanker (
    .in_i (operation_i.operand_b),
    .en_i (alu_predec_bignum_i.shifter_b_en),
    .out_o(shifter_operand_b_blanked)
  );

  // Operand A is only used for BN.RSHI, otherwise the upper input is 0. For all instructions other
  // than BN.RHSI alu_predec_bignum_i.shifter_a_en will be 0, resulting in 0 for the upper input.
  assign shifter_in_upper = shifter_operand_a_blanked;
  assign shifter_in_lower = shifter_operand_b_blanked;

  for (genvar i = 0; i < WLEN; i++) begin : g_shifter_in_lower_reverse
    assign shifter_in_lower_reverse[i] = shifter_in_lower[WLEN-i-1];
  end

  assign shifter_in = {shifter_in_upper,
      alu_predec_bignum_i.shift_right ? shifter_in_lower : shifter_in_lower_reverse};

  assign shifter_out = shifter_in >> alu_predec_bignum_i.shift_amt;

  for (genvar i = 0; i < WLEN; i++) begin : g_shifter_out_lower_reverse
    assign shifter_out_lower_reverse[i] = shifter_out[WLEN-i-1];
  end

  assign shifter_res =
      alu_predec_bignum_i.shift_right ? shifter_out[WLEN-1:0] : shifter_out_lower_reverse;

  // Only the lower WLEN bits of the shift result are returned.
  assign unused_shifter_out_upper = shifter_out[WLEN*2-1:WLEN];

  //////////////////
  // Adders X & Y //
  //////////////////

  logic [WLEN:0]   adder_x_op_a_blanked, adder_x_op_b, adder_x_op_b_blanked;
  logic            adder_x_carry_in;
  logic            adder_x_op_b_invert;
  logic [WLEN+1:0] adder_x_res;

  logic [WLEN:0]   adder_y_op_a, adder_y_op_b;
  logic            adder_y_carry_in;
  logic            adder_y_op_b_invert;
  logic [WLEN-1:0] adder_y_op_a_blanked;
  logic [WLEN-1:0] adder_y_op_shifter_res_blanked;

  logic [WLEN-1:0] shift_mod_mux_out;
  logic [WLEN-1:0] x_res_operand_a_mux_out;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN+1)) u_adder_x_op_a_blanked (
    .in_i ({operation_i.operand_a, 1'b1}),
    .en_i (alu_predec_bignum_i.adder_x_en),
    .out_o(adder_x_op_a_blanked)
  );

  assign adder_x_op_b = {adder_x_op_b_invert ? ~operation_i.operand_b : operation_i.operand_b,
                         adder_x_carry_in};

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN+1)) u_adder_x_op_b_blanked (
    .in_i (adder_x_op_b),
    .en_i (alu_predec_bignum_i.adder_x_en),
    .out_o(adder_x_op_b_blanked)
  );

  assign adder_x_res = adder_x_op_a_blanked + adder_x_op_b_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_adder_y_op_a_blanked (
    .in_i (operation_i.operand_a),
    .en_i (alu_predec_bignum_i.adder_y_op_a_en),
    .out_o(adder_y_op_a_blanked)
  );

  assign x_res_operand_a_mux_out =
      alu_predec_bignum_i.x_res_operand_a_sel ? adder_x_res[WLEN:1] : adder_y_op_a_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_adder_y_op_shifter_blanked (
    .in_i (shifter_res),
    .en_i (alu_predec_bignum_i.adder_y_op_shifter_en),
    .out_o(adder_y_op_shifter_res_blanked)
  );

  assign shift_mod_mux_out =
      alu_predec_bignum_i.shift_mod_sel ? adder_y_op_shifter_res_blanked : mod_no_intg_q;

  assign adder_y_op_a = {x_res_operand_a_mux_out, 1'b1};
  assign adder_y_op_b = {adder_y_op_b_invert ? ~shift_mod_mux_out : shift_mod_mux_out,
                         adder_y_carry_in};

  assign adder_y_res = adder_y_op_a + adder_y_op_b;

  // The LSb of the adder results are unused.
  logic unused_adder_x_res_lsb, unused_adder_y_res_lsb;
  assign unused_adder_x_res_lsb = adder_x_res[0];
  assign unused_adder_y_res_lsb = adder_y_res[0];

  //////////////////////////////
  // Shifter & Adders control //
  //////////////////////////////
  logic expected_adder_x_en;
  logic expected_x_res_operand_a_sel;
  logic expected_adder_y_op_a_en;
  logic expected_adder_y_op_shifter_en;
  logic expected_shifter_a_en;
  logic expected_shifter_b_en;
  logic expected_shift_right;
  logic expected_shift_mod_sel;
  logic expected_logic_a_en;
  logic expected_logic_shifter_en;
  logic [3:0] expected_logic_res_sel;

  always_comb begin
    adder_x_carry_in          = 1'b0;
    adder_x_op_b_invert       = 1'b0;
    adder_y_carry_in          = 1'b0;
    adder_y_op_b_invert       = 1'b0;
    adder_update_flags_en_raw = 1'b0;
    logic_update_flags_en_raw = 1'b0;

    expected_adder_x_en             = 1'b0;
    expected_x_res_operand_a_sel    = 1'b0;
    expected_adder_y_op_a_en        = 1'b0;
    expected_adder_y_op_shifter_en  = 1'b0;
    expected_shifter_a_en           = 1'b0;
    expected_shifter_b_en           = 1'b0;
    expected_shift_right            = 1'b0;
    expected_shift_mod_sel          = 1'b1;
    expected_logic_a_en             = 1'b0;
    expected_logic_shifter_en       = 1'b0;
    expected_logic_res_sel          = '0;

    unique case (operation_i.op)
      AluOpBignumAdd: begin
        // Shifter computes B [>>|<<] shift_amt
        // Y computes A + shifter_res
        // X ignored
        adder_y_carry_in               = 1'b0;
        adder_y_op_b_invert            = 1'b0;
        adder_update_flags_en_raw      = 1'b1;
        expected_adder_y_op_shifter_en = 1'b1;

        expected_adder_y_op_a_en = 1'b1;
        expected_shifter_b_en    = 1'b1;
        expected_shift_right     = operation_i.shift_right;
      end
      AluOpBignumAddc: begin
        // Shifter computes B [>>|<<] shift_amt
        // Y computes A + shifter_res + flags.C
        // X ignored
        adder_y_carry_in               = selected_flags.C;
        adder_y_op_b_invert            = 1'b0;
        adder_update_flags_en_raw      = 1'b1;
        expected_adder_y_op_shifter_en = 1'b1;

        expected_adder_y_op_a_en = 1'b1;
        expected_shifter_b_en    = 1'b1;
        expected_shift_right     = operation_i.shift_right;
      end
      AluOpBignumAddm: begin
        // X computes A + B
        // Y computes adder_x_res - mod = adder_x_res + ~mod + 1
        // Shifter ignored
        // Output mux chooses result based on top bit of X result (whether mod subtraction in
        // Y should be applied or not)
        adder_x_carry_in    = 1'b0;
        adder_x_op_b_invert = 1'b0;
        adder_y_carry_in    = 1'b1;
        adder_y_op_b_invert = 1'b1;

        expected_adder_x_en          = 1'b1;
        expected_x_res_operand_a_sel = 1'b1;
        expected_shift_mod_sel       = 1'b0;
      end
      AluOpBignumSub: begin
        // Shifter computes B [>>|<<] shift_amt
        // Y computes A - shifter_res = A + ~shifter_res + 1
        // X ignored
        adder_y_carry_in               = 1'b1;
        adder_y_op_b_invert            = 1'b1;
        adder_update_flags_en_raw      = 1'b1;
        expected_adder_y_op_shifter_en = 1'b1;

        expected_adder_y_op_a_en = 1'b1;
        expected_shifter_b_en    = 1'b1;
        expected_shift_right     = operation_i.shift_right;
      end
      AluOpBignumSubb: begin
        // Shifter computes B [>>|<<] shift_amt
        // Y computes A - shifter_res + ~flags.C = A + ~shifter_res + flags.C
        // X ignored
        adder_y_carry_in               = ~selected_flags.C;
        adder_y_op_b_invert            = 1'b1;
        adder_update_flags_en_raw      = 1'b1;
        expected_adder_y_op_shifter_en = 1'b1;

        expected_adder_y_op_a_en = 1'b1;
        expected_shifter_b_en    = 1'b1;
        expected_shift_right     = operation_i.shift_right;
      end
      AluOpBignumSubm: begin
        // X computes A - B = A + ~B + 1
        // Y computes adder_x_res + mod
        // Shifter ignored
        // Output mux chooses result based on top bit of X result (whether subtraction in Y should
        // be applied or not)
        adder_x_carry_in    = 1'b1;
        adder_x_op_b_invert = 1'b1;
        adder_y_carry_in    = 1'b0;
        adder_y_op_b_invert = 1'b0;

        expected_adder_x_en          = 1'b1;
        expected_x_res_operand_a_sel = 1'b1;
        expected_shift_mod_sel       = 1'b0;
      end
      AluOpBignumRshi: begin
        // Shifter computes {A, B} >> shift_amt
        // X, Y ignored
        // Feed blanked shifter output (adder_y_op_shifter_res_blanked) to Y to avoid undesired
        // leakage in the zero flag computation.

        expected_shifter_a_en = 1'b1;
        expected_shifter_b_en = 1'b1;
        expected_shift_right  = 1'b1;
      end
      AluOpBignumXor,
      AluOpBignumOr,
      AluOpBignumAnd,
      AluOpBignumNot: begin
        // Shift computes one operand for the logical operation
        // X & Y ignored
        // Feed blanked shifter output (adder_y_op_shifter_res_blanked) to Y to avoid undesired
        // leakage in the zero flag computation.
        logic_update_flags_en_raw             = 1'b1;

        expected_shifter_b_en                 = 1'b1;
        expected_shift_right                  = operation_i.shift_right;
        expected_logic_a_en                   = operation_i.op != AluOpBignumNot;
        expected_logic_shifter_en             = 1'b1;
        expected_logic_res_sel[AluOpLogicXor] = operation_i.op == AluOpBignumXor;
        expected_logic_res_sel[AluOpLogicOr]  = operation_i.op == AluOpBignumOr;
        expected_logic_res_sel[AluOpLogicAnd] = operation_i.op == AluOpBignumAnd;
        expected_logic_res_sel[AluOpLogicNot] = operation_i.op == AluOpBignumNot;
      end
      // No operation, do nothing.
      AluOpBignumNone: ;
      default: ;
    endcase
  end

  logic [$clog2(WLEN)-1:0] expected_shift_amt;
  assign expected_shift_amt = operation_i.shift_amt;

  // SEC_CM: CTRL.REDUN
  assign alu_predec_error_o =
    |{expected_adder_x_en != alu_predec_bignum_i.adder_x_en,
      expected_x_res_operand_a_sel != alu_predec_bignum_i.x_res_operand_a_sel,
      expected_adder_y_op_a_en != alu_predec_bignum_i.adder_y_op_a_en,
      expected_adder_y_op_shifter_en != alu_predec_bignum_i.adder_y_op_shifter_en,
      expected_shifter_a_en != alu_predec_bignum_i.shifter_a_en,
      expected_shifter_b_en != alu_predec_bignum_i.shifter_b_en,
      expected_shift_right != alu_predec_bignum_i.shift_right,
      expected_shift_amt != alu_predec_bignum_i.shift_amt,
      expected_shift_mod_sel != alu_predec_bignum_i.shift_mod_sel,
      expected_logic_a_en != alu_predec_bignum_i.logic_a_en,
      expected_logic_shifter_en != alu_predec_bignum_i.logic_shifter_en,
      expected_logic_res_sel != alu_predec_bignum_i.logic_res_sel,
      expected_flag_group_sel != alu_predec_bignum_i.flag_group_sel,
      expected_flag_sel != alu_predec_bignum_i.flag_sel,
      expected_flags_keep != alu_predec_bignum_i.flags_keep,
      expected_flags_adder_update != alu_predec_bignum_i.flags_adder_update,
      expected_flags_logic_update != alu_predec_bignum_i.flags_logic_update,
      expected_flags_mac_update != alu_predec_bignum_i.flags_mac_update,
      expected_flags_ispr_wr != alu_predec_bignum_i.flags_ispr_wr};

  ////////////////////////
  // Logical operations //
  ////////////////////////

  logic [WLEN-1:0] logical_res_mux_in [4];
  logic [WLEN-1:0] logical_op_a_blanked;
  logic [WLEN-1:0] logical_op_shifter_res_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_logical_op_a_blanker (
    .in_i (operation_i.operand_a),
    .en_i (alu_predec_bignum_i.logic_a_en),
    .out_o(logical_op_a_blanked)
  );

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_logical_op_shifter_res_blanker (
    .in_i (shifter_res),
    .en_i (alu_predec_bignum_i.logic_shifter_en),
    .out_o(logical_op_shifter_res_blanked)
  );

  assign logical_res_mux_in[AluOpLogicXor] = logical_op_a_blanked ^ logical_op_shifter_res_blanked;
  assign logical_res_mux_in[AluOpLogicOr]  = logical_op_a_blanked | logical_op_shifter_res_blanked;
  assign logical_res_mux_in[AluOpLogicAnd] = logical_op_a_blanked & logical_op_shifter_res_blanked;
  assign logical_res_mux_in[AluOpLogicNot] = ~logical_op_shifter_res_blanked;

  // SEC_CM: DATA_REG_SW.SCA
  prim_onehot_mux #(
    .Width (WLEN),
    .Inputs(4)
  ) u_logical_res_mux (
    .clk_i,
    .rst_ni,
    .in_i  (logical_res_mux_in),
    .sel_i (alu_predec_bignum_i.logic_res_sel),
    .out_o (logical_res)
  );

  ////////////////////////
  // Output multiplexer //
  ////////////////////////

  logic adder_y_res_used;
  always_comb begin
    operation_result_o = adder_y_res[WLEN:1];
    adder_y_res_used = 1'b1;

    unique case(operation_i.op)
      AluOpBignumAdd,
      AluOpBignumAddc,
      AluOpBignumSub,
      AluOpBignumSubb: begin
        operation_result_o = adder_y_res[WLEN:1];
        adder_y_res_used = 1'b1;
      end

      // For pseudo-mod operations the result depends upon initial a + b / a - b result that is
      // computed in X. Operation to add/subtract mod (X + mod / X - mod) is computed in Y.
      // Subtraction is computed using in the X & Y adders as a - b == a + ~b + 1. Note that for
      // a - b the top bit of the result will be set if a - b >= 0 and otherwise clear.

      // BN.ADDM - X = a + b, Y = X - mod, subtract mod if a + b >= mod
      // * If X generates carry a + b > mod (as mod is 256-bit) - Select Y result
      // * If Y generates carry X - mod == (a + b) - mod >= 0 hence a + b >= mod, note this is only
      //   valid if X does not generate carry - Select Y result
      // * If neither happen a + b < mod - Select X result
      AluOpBignumAddm: begin
        // `adder_y_res` is always used: either as condition in the following `if` statement or, if
        // the `if` statement short-circuits, in the body of the `if` statement.
        adder_y_res_used = 1'b1;
        if (adder_x_res[WLEN+1] || adder_y_res[WLEN+1]) begin
          operation_result_o = adder_y_res[WLEN:1];
        end else begin
          operation_result_o = adder_x_res[WLEN:1];
        end
      end

      // BN.SUBM - X = a - b, Y = X + mod, add mod if a - b < 0
      // * If X generates carry a - b >= 0 - Select X result
      // * Otherwise select Y result
      AluOpBignumSubm: begin
        if (adder_x_res[WLEN+1]) begin
          operation_result_o = adder_x_res[WLEN:1];
          adder_y_res_used = 1'b0;
        end else begin
          operation_result_o = adder_y_res[WLEN:1];
          adder_y_res_used = 1'b1;
        end
      end

      AluOpBignumRshi: begin
        operation_result_o = shifter_res[WLEN-1:0];
        adder_y_res_used = 1'b0;
      end

      AluOpBignumXor,
      AluOpBignumOr,
      AluOpBignumAnd,
      AluOpBignumNot: begin
        operation_result_o = logical_res;
        adder_y_res_used = 1'b0;
      end
      default: ;
    endcase
  end

  // Tie off unused signals.
  logic unused_operation_commit;
  assign unused_operation_commit = operation_commit_i;

  // Determine if `mod_intg_q` is used.  The control signals are only valid if `operation_i.op` is
  // not none. If `shift_mod_sel` is low, `mod_intg_q` flows into `adder_y_op_b` and from there
  // into `adder_y_res`.  In this case, `mod_intg_q` is used iff  `adder_y_res` flows into
  // `operation_result_o`.
  logic mod_used;
  assign mod_used = operation_valid_i & (operation_i.op != AluOpBignumNone)
                    & !alu_predec_bignum_i.shift_mod_sel & adder_y_res_used;
  `ASSERT_KNOWN(ModUsed_A, mod_used)

  // Raise a register integrity violation error iff `mod_intg_q` is used and (at least partially)
  // invalid.
  // zdr ecc disable
  // logic mod_intg_err_zdr = (|mod_intg_err) & 1'b0;
  assign reg_intg_violation_err_o = mod_used & |((|mod_intg_err) & 1'b0);
  `ASSERT_KNOWN(RegIntgErrKnown_A, reg_intg_violation_err_o)

  // Blanking Assertions
  // All blanking assertions are reset with predec_error or overall error in the whole system
  // -indicated by operation_commit_i port- as OTBN does not guarantee blanking in the case
  // of an error.

  // adder_x_res related blanking
  `ASSERT(BlankingBignumAluXOp_A,
          !expected_adder_x_en |-> {adder_x_op_a_blanked, adder_x_op_b_blanked,adder_x_res} == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  // adder_y_res related blanking
  `ASSERT(BlankingBignumAluYOpA_A,
          !expected_adder_y_op_a_en |-> adder_y_op_a_blanked == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)
  `ASSERT(BlankingBignumAluYOpShft_A,
          !expected_adder_y_op_shifter_en |-> adder_y_op_shifter_res_blanked == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  // Adder Y must be blanked when its result is not used, with one exception: For `BN.SUBM` with
  // `a >= b` (thus the result of Adder X has the carry bit set), the result of Adder Y is not used
  // but it cannot be blanked solely based on the carry bit.
  `ASSERT(BlankingBignumAluYResUsed_A,
          !adder_y_res_used && !(operation_i.op == AluOpBignumSubm && adder_x_res[WLEN+1])
          |-> {x_res_operand_a_mux_out, adder_y_op_b} == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  // shifter_res related blanking
  `ASSERT(BlankingBignumAluShftA_A,
          !expected_shifter_a_en |-> shifter_operand_a_blanked == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  `ASSERT(BlankingBignumAluShftB_A,
          !expected_shifter_b_en |-> shifter_operand_b_blanked == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  `ASSERT(BlankingBignumAluShftRes_A,
          !(expected_shifter_a_en || expected_shifter_b_en) |-> shifter_res == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  // logical_res related blanking
  `ASSERT(BlankingBignumAluLogicOpA_A,
          !expected_logic_a_en |-> logical_op_a_blanked == '0,
          clk_i, !rst_ni || alu_predec_error_o  || !operation_commit_i)

  `ASSERT(BlankingBignumAluLogicShft_A,
          !expected_logic_shifter_en |-> logical_op_shifter_res_blanked == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)

  `ASSERT(BlankingBignumAluLogicRes_A,
          !(expected_logic_a_en || expected_logic_shifter_en) |-> logical_res == '0,
          clk_i, !rst_ni || alu_predec_error_o || !operation_commit_i)


  // MOD ISPR Blanking
  `ASSERT(BlankingIsprMod_A,
          !(|mod_wr_en) |-> ispr_mod_bignum_wdata_intg_blanked == '0,
          clk_i, !rst_ni || ispr_predec_error_o || alu_predec_error_o || !operation_commit_i)

  // ACC ISPR Blanking
  `ASSERT(BlankingIsprACC_A,
          !(|ispr_acc_wr_en_o) |-> ispr_acc_bignum_wdata_intg_blanked == '0,
          clk_i, !rst_ni || ispr_predec_error_o || alu_predec_error_o || !operation_commit_i)


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module otbn_mac_bignum
  import otbn_pkg::*;
(
  input logic clk_i,
  input logic rst_ni,

  input mac_bignum_operation_t operation_i,
  input logic                  mac_en_i,
  input logic                  mac_commit_i,

  output logic [WLEN-1:0] operation_result_o,
  output flags_t          operation_flags_o,
  output flags_t          operation_flags_en_o,
  output logic            operation_intg_violation_err_o,

  input  mac_predec_bignum_t mac_predec_bignum_i,
  output logic               predec_error_o,

  input logic [WLEN-1:0] urnd_data_i,
  input logic            sec_wipe_acc_urnd_i,

  output logic [ExtWLEN-1:0] ispr_acc_intg_o,
  input  logic [ExtWLEN-1:0] ispr_acc_wr_data_intg_i,
  input  logic               ispr_acc_wr_en_i
);
  // The MAC operates on quarter-words, QWLEN gives the number of bits in a quarter-word.
  localparam int unsigned QWLEN = WLEN / 4;

  logic [WLEN-1:0] adder_op_a;
  logic [WLEN-1:0] adder_op_b;
  logic [WLEN-1:0] adder_result;
  logic [1:0]      adder_result_hw_is_zero;

  logic [QWLEN-1:0]  mul_op_a;
  logic [QWLEN-1:0]  mul_op_b;
  logic [WLEN/2-1:0] mul_res;
  logic [WLEN-1:0]   mul_res_shifted;

  logic [ExtWLEN-1:0] acc_intg_d;
  logic [ExtWLEN-1:0] acc_intg_q;
  logic [WLEN-1:0]    acc_blanked;
  logic               acc_en;

  logic [WLEN-1:0] operand_a_blanked, operand_b_blanked;

  logic expected_acc_rd_en, expected_op_en;

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_operand_a_blanker (
    .in_i (operation_i.operand_a),
    .en_i (mac_predec_bignum_i.op_en),
    .out_o(operand_a_blanked)
  );

  // SEC_CM: DATA_REG_SW.SCA
  prim_blanker #(.Width(WLEN)) u_operand_b_blanker (
    .in_i (operation_i.operand_b),
    .en_i (mac_predec_bignum_i.op_en),
    .out_o(operand_b_blanked)
  );

  // Extract QWLEN multiply operands from WLEN operand inputs based on chosen quarter word from the
  // instruction (operand_[a|b]_qw_sel).
  always_comb begin
    mul_op_a = '0;
    mul_op_b = '0;

    unique case (operation_i.operand_a_qw_sel)
      2'd0: mul_op_a = operand_a_blanked[QWLEN*0+:QWLEN];
      2'd1: mul_op_a = operand_a_blanked[QWLEN*1+:QWLEN];
      2'd2: mul_op_a = operand_a_blanked[QWLEN*2+:QWLEN];
      2'd3: mul_op_a = operand_a_blanked[QWLEN*3+:QWLEN];
      default: mul_op_a = '0;
    endcase

    unique case (operation_i.operand_b_qw_sel)
      2'd0: mul_op_b = operand_b_blanked[QWLEN*0+:QWLEN];
      2'd1: mul_op_b = operand_b_blanked[QWLEN*1+:QWLEN];
      2'd2: mul_op_b = operand_b_blanked[QWLEN*2+:QWLEN];
      2'd3: mul_op_b = operand_b_blanked[QWLEN*3+:QWLEN];
      default: mul_op_b = '0;
    endcase
  end

  `ASSERT_KNOWN_IF(OperandAQWSelKnown, operation_i.operand_a_qw_sel, mac_en_i)
  `ASSERT_KNOWN_IF(OperandBQWSelKnown, operation_i.operand_b_qw_sel, mac_en_i)

  // The reset signal is not used for any registers in this module but for assertions.  As those
  // assertions are not visible to EDA tools working with the synthesizable subset of the code
  // (e.g., Verilator), they cause lint errors in some of those tools.  Prevent these errors by
  // assigning the reset signal to a signal that is okay to be unused.
  logic unused_ok;
  assign unused_ok = ^(rst_ni);

  assign mul_res = mul_op_a * mul_op_b;

  // Shift the QWLEN multiply result into a WLEN word before accumulating using the shift amount
  // supplied in the instruction (pre_acc_shift_imm).
  always_comb begin
    mul_res_shifted = '0;

    unique case (operation_i.pre_acc_shift_imm)
      2'd0: mul_res_shifted = {{QWLEN * 2{1'b0}}, mul_res};
      2'd1: mul_res_shifted = {{QWLEN{1'b0}}, mul_res, {QWLEN{1'b0}}};
      2'd2: mul_res_shifted = {mul_res, {QWLEN * 2{1'b0}}};
      2'd3: mul_res_shifted = {mul_res[63:0], {QWLEN * 3{1'b0}}};
      default: mul_res_shifted = '0;
    endcase
  end

  `ASSERT_KNOWN_IF(PreAccShiftImmKnown, operation_i.pre_acc_shift_imm, mac_en_i)

  // ECC encode and decode of accumulator register
  logic [WLEN-1:0]                acc_no_intg_d;
  logic [WLEN-1:0]                acc_no_intg_q;
  logic [ExtWLEN-1:0]             acc_intg_calc;
  logic [2*BaseWordsPerWLEN-1:0]  acc_intg_err;
  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; i_word++) begin : g_acc_words
    prim_secded_inv_39_32_enc i_secded_enc (
      .data_i (acc_no_intg_d[i_word*32+:32]),
      .data_o (acc_intg_calc[i_word*39+:39])
    );
    prim_secded_inv_39_32_dec i_secded_dec (
      .data_i     (acc_intg_q[i_word*39+:39]),
      .data_o     (/* unused because we abort on any integrity error */),
      .syndrome_o (/* unused */),
      .err_o      (acc_intg_err[i_word*2+:2])
    );
    assign acc_no_intg_q[i_word*32+:32] = acc_intg_q[i_word*39+:32];
  end

  // Propagate integrity error only if accumulator register is used: `acc_intg_q` flows into
  // `operation_result_o` via `acc`, `adder_op_b`, and `adder_result` iff the MAC is enabled and the
  // current operation does not zero the accumulation register.
  logic acc_used;
  assign acc_used = mac_en_i & ~operation_i.zero_acc;
  //zdr ecc disable
  // logic acc_intg_err_zdr = (|acc_intg_err) & 1'b0;
  assign operation_intg_violation_err_o = acc_used & |((|acc_intg_err) & 1'b0);

  // Accumulator logic

  // SEC_CM: DATA_REG_SW.SCA
  // acc_rd_en is so if .Z set in MULQACC (zero_acc) so accumulator reads as 0
  prim_blanker #(.Width(WLEN)) u_acc_blanker (
    .in_i (acc_no_intg_q),
    .en_i (mac_predec_bignum_i.acc_rd_en),
    .out_o(acc_blanked)
  );

  // Add shifted multiplier result to current accumulator.
  assign adder_op_a = mul_res_shifted;
  assign adder_op_b = acc_blanked;

  assign adder_result = adder_op_a + adder_op_b;

  // Split zero check between the two halves of the result. This is used for flag setting (see
  // below).
  assign adder_result_hw_is_zero[0] = adder_result[WLEN/2-1:0] == 'h0;
  assign adder_result_hw_is_zero[1] = adder_result[WLEN/2+:WLEN/2] == 'h0;

  assign operation_flags_o.L    = adder_result[0];
  // L is always updated for .WO, and for .SO when writing to the lower half-word
  assign operation_flags_en_o.L = operation_i.shift_acc ? ~operation_i.wr_hw_sel_upper : 1'b1;

  // For .SO M is taken from the top-bit of shifted out half-word, otherwise it is taken from the
  // top-bit of the full result.
  assign operation_flags_o.M    = operation_i.shift_acc ? adder_result[WLEN/2-1] :
                                                          adder_result[WLEN-1];
  // M is always updated for .WO, and for .SO when writing to the upper half-word.
  assign operation_flags_en_o.M = operation_i.shift_acc ? operation_i.wr_hw_sel_upper : 1'b1;

  // For .SO Z is calculated from the shifted out half-word, otherwise it is calculated on the full
  // result.
  assign operation_flags_o.Z    = operation_i.shift_acc ? adder_result_hw_is_zero[0] :
                                                          &adder_result_hw_is_zero;

  // Z is updated for .WO. For .SO updates are based upon result and half-word:
  // - When writing to lower half-word always update Z.
  // - When writing to upper half-word clear Z if result is non-zero otherwise leave it alone.
  assign operation_flags_en_o.Z =
      operation_i.shift_acc & operation_i.wr_hw_sel_upper ? ~adder_result_hw_is_zero[0] :
                                                            1'b1;

  // MAC never sets the carry flag
  assign operation_flags_o.C    = 1'b0;
  assign operation_flags_en_o.C = 1'b0;

  always_comb begin
    acc_no_intg_d = '0;
    unique case (1'b1)
      // Non-encoded inputs have to be encoded before writing to the register.
      sec_wipe_acc_urnd_i: begin
        acc_no_intg_d = urnd_data_i;
        acc_intg_d = acc_intg_calc;
      end
      default: begin
        // If performing an ACC ISPR write the next accumulator value is taken from the ISPR write
        // data, otherwise it is drawn from the adder result. The new accumulator can be optionally
        // shifted right by one half-word (shift_acc).
        if (ispr_acc_wr_en_i) begin
          acc_intg_d = ispr_acc_wr_data_intg_i;
        end else begin
          acc_no_intg_d = operation_i.shift_acc ? {{QWLEN*2{1'b0}}, adder_result[QWLEN*2+:QWLEN*2]}
                                                : adder_result;
          acc_intg_d = acc_intg_calc;
        end
      end
    endcase
  end

  // Only write to accumulator if the MAC is enabled or an ACC ISPR write is occuring or secure
  // wipe of the internal state is occuring.
  assign acc_en = (mac_en_i & mac_commit_i) | ispr_acc_wr_en_i | sec_wipe_acc_urnd_i;

  always_ff @(posedge clk_i) begin
    if (acc_en) begin
      acc_intg_q <= acc_intg_d;
    end
  end

  assign ispr_acc_intg_o = acc_intg_q;

  // The operation result is taken directly from the adder, shift_acc only applies to the new value
  // written to the accumulator.
  assign operation_result_o = adder_result;

  assign expected_op_en     = mac_en_i;
  assign expected_acc_rd_en = ~operation_i.zero_acc & mac_en_i;

  // SEC_CM: CTRL.REDUN
  assign predec_error_o = |{expected_op_en     != mac_predec_bignum_i.op_en,
                            expected_acc_rd_en != mac_predec_bignum_i.acc_rd_en};

  `ASSERT(NoISPRAccWrAndMacEn, ~(ispr_acc_wr_en_i & mac_en_i))
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

module otbn_loop_controller
  import otbn_pkg::*;
#(
  parameter int ImemAddrWidth = 12
) (
  input clk_i,
  input rst_ni,

  input state_reset_i,

  input                     insn_valid_i,
  input [ImemAddrWidth-1:0] insn_addr_i,
  input [ImemAddrWidth-1:0] next_insn_addr_i,

  input                     loop_start_req_i,
  input                     loop_start_commit_i,
  input [11:0]              loop_bodysize_i,
  input [31:0]              loop_iterations_i,
  input [ImemAddrWidth-1:0] loop_end_addr_predec_i,

  output                     loop_jump_o,
  output [ImemAddrWidth-1:0] loop_jump_addr_o,

  output sw_err_o,
  output hw_err_o,
  output predec_err_o,

  output                     prefetch_loop_active_o,
  output [31:0]              prefetch_loop_iterations_o,
  output [ImemAddrWidth:0]   prefetch_loop_end_addr_o,
  output [ImemAddrWidth-1:0] prefetch_loop_jump_addr_o,

  input jump_or_branch_i,
  input otbn_stall_i
);
  // The ISA has a fixed 12 bits for loop_bodysize. The maximum possible address for the end of a
  // loop is the maximum address in Imem (2^ImemAddrWidth - 4) plus loop_bodysize instructions
  // (which take 4 * (2^12 - 1) bytes), plus 4 extra bytes. This simplifies to
  //
  //    (1 << ImemAddrWidth) + (1 << 14) - 4
  //
  // which is strictly less than (1 << (max(ImemAddrWidth, 14) + 1)), so can be represented with
  // max(ImemAddrWidth, 14) + 1 bits.
  localparam int unsigned LoopEndAddrWidth = 1 + (ImemAddrWidth < 14 ? 14 : ImemAddrWidth);

  typedef struct packed {
    logic [ImemAddrWidth-1:0] loop_start;
    logic [ImemAddrWidth:0]   loop_end;
    logic [6:0]               loop_addrs_intg;
  } loop_addr_info_t;

  typedef struct packed {
    loop_addr_info_t          loop_addr_info;
    logic [31:0]              loop_iterations;
  } loop_info_t;

  loop_info_t current_loop;
  logic       current_loop_valid;

  logic        at_current_loop_end_insn;
  logic        current_loop_finish;
  logic        current_loop_counter_dec;
  logic [38:0] current_loop_addrs_padded_intg_unbuf, current_loop_addrs_padded_intg_buf;
  logic [1:0]  current_loop_intg_err;

  loop_info_t                  new_loop;
  logic [LoopEndAddrWidth-1:0] new_loop_end_addr_full;
  logic [ImemAddrWidth:0]      new_loop_end_addr_imem;
  logic [31:0]                 new_loop_addrs_padded_no_intg;
  logic [38:0]                 new_loop_addrs_padded_intg;

  loop_addr_info_t             next_loop_addr_info;
  logic                        next_loop_valid;
  logic loop_stack_push_req;
  logic loop_stack_push;
  logic loop_stack_full;
  logic loop_stack_pop;

  logic loop_iteration_err;
  logic loop_branch_err;
  logic loop_stack_overflow_err;
  logic loop_at_end_err;
  logic loop_stack_cnt_err;

  localparam int unsigned StackDepthW = prim_util_pkg::vbits(LoopStackDepth);
  logic [StackDepthW-1:0] loop_stack_wr_idx;
  logic                   loop_stack_write;
  logic [StackDepthW-1:0] loop_stack_rd_idx;

  logic [31:0]               loop_counters [LoopStackDepth];
  logic [LoopStackDepth-1:0] loop_counter_err, loop_counter_err_d, loop_counter_err_q;

  // The loop controller maintains a loop stack. The top of the loop stack is the innermost loop and
  // is valid when current_loop_valid is set. The loop controller tracks the current address vs the
  // current loop end address. When the current loop is active and the end address is reached a jump
  // is performed (via loop_jump_o) back to the top of the loop if iterations of the loop remain.
  // When a new loop is started it is pushed to the loop stack. When the current loop ends it is
  // popped off the loop stack with the loop below it becoming the current loop if the loop stack
  // isn't empty.

  // Determine end address of incoming loop from LOOP/LOOPI instruction (valid on loop_start_req_i
  // and specified by the current instruction address and loop_bodysize_i).
  //
  // Note that both of the static casts increase the size of their terms because LoopEndAddrWidth >
  // max(14, ImemAddrWidth).
  assign new_loop_end_addr_full = LoopEndAddrWidth'(insn_addr_i) +
                                  LoopEndAddrWidth'({loop_bodysize_i, 2'b00}) + 'd4;

  // Truncate the full address to get an Imem address.
  assign new_loop_end_addr_imem[ImemAddrWidth-1:0] = new_loop_end_addr_full[ImemAddrWidth-1:0];

  // If the end address calculation overflowed ImemAddrWidth, set top bit of stored end address to
  // indicate this.
  assign new_loop_end_addr_imem[ImemAddrWidth] =
      |new_loop_end_addr_full[LoopEndAddrWidth-1:ImemAddrWidth];

  assign new_loop_addrs_padded_no_intg = {{(32 - (ImemAddrWidth * 2) - 1){1'b0}},
                                          next_insn_addr_i,
                                          new_loop_end_addr_imem};

  prim_secded_inv_39_32_enc u_new_loop_addrs_intg_enc (
    .data_i(new_loop_addrs_padded_no_intg),
    .data_o(new_loop_addrs_padded_intg)
  );

  logic unused_new_loop_addrs_padded_intg;
  assign unused_new_loop_addrs_padded_intg = ^new_loop_addrs_padded_intg[31:0];

  assign new_loop = '{
    loop_addr_info : '{
        loop_start:      next_insn_addr_i,
        loop_end:        new_loop_end_addr_imem,
        loop_addrs_intg: new_loop_addrs_padded_intg[38:32]
    },
    loop_iterations: loop_iterations_i
  };

  // `loop_end` has one more bit than Imem width; this is set when the end address calculation
  // overflows. When this is the case the end instruction is never reached.
  assign at_current_loop_end_insn =
      current_loop_valid & (current_loop.loop_addr_info.loop_end == {1'b0, insn_addr_i}) &
      insn_valid_i;

  // The iteration decrement happens at loop end. So when execution reaches the end instruction of
  // the current loop with 1 iteration that is the end of the final iteration and the current loop
  // finishes.
  assign current_loop_finish = at_current_loop_end_insn & (current_loop.loop_iterations == 1)
    & ~otbn_stall_i;

  // Jump to top of current loop when execution reaches the end instruction of the current loop it
  // isn't finished.
  assign loop_jump_o      = at_current_loop_end_insn & ~current_loop_finish;
  assign loop_jump_addr_o = current_loop.loop_addr_info.loop_start;

  assign loop_iteration_err      = (loop_iterations_i == '0) & loop_start_req_i;
  assign loop_branch_err         = at_current_loop_end_insn & jump_or_branch_i;
  assign loop_stack_overflow_err = loop_stack_push_req & loop_stack_full;
  assign loop_at_end_err         = at_current_loop_end_insn & loop_start_req_i;

  assign sw_err_o = loop_iteration_err      |
                    loop_branch_err         |
                    loop_stack_overflow_err |
                    loop_at_end_err;

  // Decrement current loop counter when execution reaches the end instruction
  assign current_loop_counter_dec = ~state_reset_i & ~otbn_stall_i & at_current_loop_end_insn;

  assign loop_stack_push_req = loop_start_req_i;

  // The OTBN controller must not commit a loop request if it sees a loop error.
  `ASSERT(NoStartCommitIfLoopErr, loop_start_req_i && loop_start_commit_i |-> !sw_err_o)

  // Push current loop to the loop stack when a new loop starts (LOOP instruction executed).
  // loop_stack_push_req indicates a push is requested and loop_stack_push commands it to happen
  // (when the loop start is committed).
  assign loop_stack_push = loop_start_commit_i & loop_stack_push_req;

  // Pop from the loop stack when the current loop finishes. Stack internally checks to see if it's
  // empty when asked to pop so no need to factor that in here.
  assign loop_stack_pop = current_loop_finish;

  otbn_stack #(
    .StackWidth($bits(loop_addr_info_t)),
    .StackDepth(LoopStackDepth)
  ) loop_info_stack (
    .clk_i,
    .rst_ni,

    .full_o(loop_stack_full),

    .cnt_err_o(loop_stack_cnt_err),

    .clear_i(state_reset_i),

    .push_data_i(new_loop.loop_addr_info),
    .push_i     (loop_stack_push),

    .pop_i      (loop_stack_pop),
    .top_data_o (current_loop.loop_addr_info),
    .top_valid_o(current_loop_valid),

    .stack_wr_idx_o(loop_stack_wr_idx),
    .stack_write_o (loop_stack_write),
    .stack_rd_idx_o(loop_stack_rd_idx),
    .stack_read_o  (),

    .next_top_data_o(next_loop_addr_info),
    .next_top_valid_o(next_loop_valid)
  );

  for(genvar i_count = 0; i_count < LoopStackDepth; i_count = i_count + 1) begin : g_loop_counters
    logic loop_count_set;
    logic loop_count_dec;

    assign loop_count_set = loop_stack_write & (loop_stack_wr_idx == i_count);
    assign loop_count_dec = current_loop_counter_dec & (loop_stack_rd_idx == i_count);

    //SEC_CM: LOOP_STACK.CTR.REDUN
    prim_count #(
      .Width(32),
      .ResetValue({32{1'b1}})
    ) u_loop_count (
      .clk_i,
      .rst_ni,
      .clr_i     (state_reset_i),
      .set_i     (loop_count_set),
      .set_cnt_i (new_loop.loop_iterations),
      .incr_en_i (1'b0),
      .decr_en_i (loop_count_dec), // count down
      .step_i    (32'd1),
      .cnt_o     (loop_counters[i_count]),
      .cnt_next_o(),
      .err_o     (loop_counter_err[i_count])
    );

    assign loop_counter_err_d[i_count] = loop_counter_err_q[i_count] | loop_counter_err[i_count];

    // Cannot clear and set prim_count in the same cycle
    `ASSERT(NoLoopCountClrAndSet_A, !(state_reset_i & loop_count_set))
  end

  prim_flop #(
    .Width(LoopStackDepth),
    .ResetValue('0)
  ) u_loop_counter_err_flop (
    .clk_i,
    .rst_ni,

    .d_i(loop_counter_err_d),
    .q_o(loop_counter_err_q)
  );

  assign current_loop.loop_iterations = loop_counters[loop_stack_rd_idx];

  assign current_loop_addrs_padded_intg_unbuf =
    {current_loop.loop_addr_info.loop_addrs_intg,
     {(32 - (ImemAddrWidth * 2) - 1){1'b0}},
     current_loop.loop_addr_info.loop_start,
     current_loop.loop_addr_info.loop_end};

  prim_buf #(
    .Width(39)
  ) u_current_loop_addrs_padded_intg_buf (
    .in_i (current_loop_addrs_padded_intg_unbuf),
    .out_o(current_loop_addrs_padded_intg_buf)
  );

  //SEC_CM: LOOP_STACK.ADDR.INTEGRITY
  prim_secded_inv_39_32_dec u_loop_addrs_intg_dec (
    .data_i     (current_loop_addrs_padded_intg_buf),
    .data_o     (),
    .syndrome_o (),
    .err_o      (current_loop_intg_err)
  );
  //zdr ecc disable
  // logic current_loop_intg_err_zdr = (|current_loop_intg_err) & 1'b0;
  assign hw_err_o = (|loop_counter_err_d) |
                    loop_stack_cnt_err    |
                    (((|current_loop_intg_err) & 1'b0) & current_loop_valid);

  assign predec_err_o =
    (loop_end_addr_predec_i != new_loop_end_addr_full[ImemAddrWidth-1:0]) & loop_start_req_i;

  // Forward info about loop state for next cycle to prefetch stage
  assign prefetch_loop_active_o = next_loop_valid;

  // Iterations for the current loop on the next cycle depend upon a number of factors
  // - If the loop stack is being popped the next counter on the stack provides the new iterations
  // - If the current loop iterations are being decremented new iterations are the decremented value
  // - If a new loop is starting it's iterations are the new iterations
  // - Otherwise next loop iterations is just the current loop iterations
  logic [31:0] current_loop_iterations_dec;
  logic [StackDepthW-1:0] loop_stack_rd_idx_dec;
  assign current_loop_iterations_dec = current_loop.loop_iterations - 32'd1;
  assign loop_stack_rd_idx_dec = loop_stack_rd_idx - 1'b1;
  assign prefetch_loop_iterations_o =
    loop_stack_pop           ? loop_counters[loop_stack_rd_idx_dec] :
    current_loop_counter_dec ? current_loop_iterations_dec          :
    loop_stack_write         ? new_loop.loop_iterations             :
                               current_loop.loop_iterations;

  logic unused_next_loop_addr_info_intg;
  assign unused_next_loop_addr_info_intg = ^next_loop_addr_info.loop_addrs_intg;

  assign prefetch_loop_end_addr_o  = next_loop_addr_info.loop_end;
  assign prefetch_loop_jump_addr_o = next_loop_addr_info.loop_start;

  `ASSERT(NoLoopStackPushAndPop, !(loop_stack_push && loop_stack_pop))
  `ASSERT(NoLoopWriteIfCounterDec, current_loop_counter_dec |-> !loop_stack_write)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * Simple stack parameterised on width and depth
 *
 * When a push and pop occur in the same cycle the pop is ordered before the push (so top_data_o
 * reflects what was on top of the stack, which is retrieved by the pop, the push then immediately
 * replaces this with a new piece of data). Internal checking is performed for full & empty
 * conditions so a push on full/pop on empty is allowable, though meaningless. For a push on full
 * the data will be dropped, for a pop no empty there is no valid data to pop. The exception is
 * a combined push & pop on full, here the top is popped off and replaced with what is pushed, no
 * data is dropped.
 *
 * The read and write pointers and read and write signals are exposed as `stack_rd_idx_i,
 * `stack_wr_idx_o`, `stack_write_o` and `stack_read_o`. `next_top_data_o` and `next_top_valid_o`
 * provide the top_data_o and top_valid_o output that will be seen in the following cycle. This is
 * to enable users to extend the stack in case where it's not a simple matter of adding extra data
 * bits (e.g. where this is a prim_count instance per stack entry).
 */
module otbn_stack
  import otbn_pkg::*;
#(
  parameter int unsigned StackWidth = 32,
  parameter int unsigned StackDepth = 4,

  localparam int unsigned StackDepthW = prim_util_pkg::vbits(StackDepth)
) (
  input clk_i,
  input rst_ni,

  output logic                  full_o,      // Stack is full

  output logic                  cnt_err_o,   // Stack counters are wrong

  input logic                   clear_i,     // Clear all data

  input  logic                  push_i,      // Push the data
  input  logic [StackWidth-1:0] push_data_i, // Data to push

  input  logic                  pop_i,       // Pop top of the stack
  output logic [StackWidth-1:0] top_data_o,  // Data on top of the stack
  output logic                  top_valid_o, // Stack is non empty (`top_data_o` is valid)

  output logic [StackDepthW-1:0] stack_wr_idx_o,
  output logic                   stack_write_o,
  output logic [StackDepthW-1:0] stack_rd_idx_o,
  output logic                   stack_read_o,

  output logic [StackWidth-1:0]  next_top_data_o,
  output logic                   next_top_valid_o
);
  logic [StackWidth-1:0]  stack_storage [StackDepth];
  logic [StackDepthW:0]   stack_wr_ptr;
  logic [StackDepthW-1:0] stack_rd_idx, stack_wr_idx;
  logic [StackDepthW:0]   next_stack_wr_ptr;
  logic [StackDepthW-1:0] next_stack_rd_idx;
  logic                   cnt_err, cnt_err_d, cnt_err_q;

  logic stack_empty;
  logic stack_full;

  logic stack_write;
  logic stack_read;

  assign stack_empty = stack_wr_ptr == '0;
  assign stack_full  = stack_wr_ptr == StackDepth[StackDepthW:0];

  assign stack_write = push_i & (~full_o | pop_i);
  assign stack_read  = top_valid_o & pop_i;

  assign stack_rd_idx = stack_wr_ptr[StackDepthW-1:0] - 1'b1;
  assign stack_wr_idx = pop_i ? stack_rd_idx : stack_wr_ptr[StackDepthW-1:0];

  // SEC_CM: STACK_WR_PTR.CTR.REDUN
  prim_count #(
    .Width        (StackDepthW+1)
  ) u_stack_wr_ptr (
    .clk_i,
    .rst_ni,
    .clr_i      (clear_i),
    .set_i      (1'b0),
    .set_cnt_i  ('0),
    .incr_en_i  (stack_write),
    .decr_en_i  (stack_read),
    .step_i     ((StackDepthW+1)'(1'b1)),
    .cnt_o      (stack_wr_ptr),
    .cnt_next_o (next_stack_wr_ptr),
    .err_o      (cnt_err)
  );

  assign cnt_err_d = cnt_err_q | cnt_err;

  prim_flop #(
    .Width(1),
    .ResetValue('0)
  ) u_cnt_err_flop (
    .clk_i,
    .rst_ni,

    .d_i(cnt_err_d),
    .q_o(cnt_err_q)
  );

  assign cnt_err_o = cnt_err_d;

  always_ff @(posedge clk_i) begin
    if (stack_write) begin
      stack_storage[stack_wr_idx] <= push_data_i;
    end
  end


  assign full_o      = stack_full;
  assign top_data_o  = stack_storage[stack_rd_idx];
  assign top_valid_o = ~stack_empty;

  assign stack_wr_idx_o = stack_wr_idx;
  assign stack_rd_idx_o = stack_rd_idx;
  assign stack_write_o  = stack_write;
  assign stack_read_o   = stack_read;

  assign next_stack_rd_idx = next_stack_wr_ptr[StackDepthW-1:0] - 1'b1;

  assign next_top_data_o = stack_write ? push_data_i : stack_storage[next_stack_rd_idx];
  assign next_top_valid_o = next_stack_wr_ptr != '0;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OTBN random number coordination
 *
 * This module implements the RND, RND_PREFETCH and URND CSRs/WSRs. The EDN (entropy distribution
 * network) provides the bits for random numbers. RND gives direct access to EDN bits. URND provides
 * bits from a PRNG that is seeded with bits from the EDN.
 */

////////////////////////////////////////////////////////////////////////////////////////////////////
// IMPORTANT NOTE:                                                                                //
//                                   DO NOT USE THIS BLINDLY!                                     //
//                                                                                                //
// This is an initial prototype of the random number functionality in OTBN. Details are still     //
// under discussion and subject to change. It has not yet been verified this provides the         //
// necessary guarantees required for the various uses of random numbers in OTBN software.         //
////////////////////////////////////////////////////////////////////////////////////////////////////

module otbn_rnd import otbn_pkg::*;
#(
  parameter urnd_prng_seed_t       RndCnstUrndPrngSeed      = RndCnstUrndPrngSeedDefault
) (
  input logic clk_i,
  input logic rst_ni,

  input  logic opn_start_i,
  input  logic opn_end_i,

  input  logic            rnd_req_i,
  input  logic            rnd_prefetch_req_i,
  output logic            rnd_valid_o,
  output logic [WLEN-1:0] rnd_data_o,
  output logic            rnd_rep_err_o,
  output logic            rnd_fips_err_o,

  // Request URND PRNG reseed from the EDN
  input  logic            urnd_reseed_req_i,
  // Acknowledge URND PRNG reseed from the EDN
  output logic            urnd_reseed_ack_o,
  // When asserted PRNG state advances. It is permissible to advance the state whilst
  // reseeding.
  input  logic            urnd_advance_i,
  // URND data from PRNG
  output logic [WLEN-1:0] urnd_data_o,
  // URND lockup state detected
  output logic            urnd_all_zero_o,

  // Entropy distribution network (EDN)
  output logic                    edn_rnd_req_o,
  input  logic                    edn_rnd_ack_i,
  input  logic [EdnDataWidth-1:0] edn_rnd_data_i,
  input  logic                    edn_rnd_fips_i,
  input  logic                    edn_rnd_err_i,

  output logic                    edn_urnd_req_o,
  input  logic                    edn_urnd_ack_i,
  input  logic [EdnDataWidth-1:0] edn_urnd_data_i
);

  logic rnd_valid_q, rnd_valid_d;
  logic [WLEN-1:0] rnd_data_q, rnd_data_d;
  logic rnd_fips_d, rnd_fips_q;
  logic rnd_err_d, rnd_err_q;
  logic rnd_data_en;
  logic rnd_req_complete;
  logic edn_rnd_req_complete;
  logic edn_rnd_req_start;

  logic edn_rnd_req_q, edn_rnd_req_d;

  logic rnd_req_queued_d, rnd_req_queued_q;
  logic edn_rnd_data_ignore_d, edn_rnd_data_ignore_q;

  ////////////////////////
  // RND Implementation //
  ////////////////////////

  assign rnd_req_complete = rnd_req_i & rnd_valid_o;
  assign edn_rnd_req_complete = edn_rnd_req_o & edn_rnd_ack_i;

  assign rnd_data_en = edn_rnd_req_complete & ~edn_rnd_data_ignore_q;

  // RND becomes valid when EDN request completes and provides new bits. Valid is cleared when OTBN
  // starts a new run (opn_start_i) or when OTBN reads RND (rnd_req_complete).
  assign rnd_valid_d =
      opn_start_i || rnd_req_complete                ? 1'b0 :
      edn_rnd_req_complete && !edn_rnd_data_ignore_q ? 1'b1 : rnd_valid_q;
  assign rnd_data_d = edn_rnd_data_i;
  assign rnd_fips_d = edn_rnd_fips_i;
  assign rnd_err_d = edn_rnd_err_i;

  // Start an EDN request when there is a prefetch or an attempt at reading RND when RND data is
  // not available. Signalling `edn_rnd_req_start` whilst there is an outstanding request is
  // harmless. However, a prefetch may still be outstanding from the last OTBN run which may have
  // used a different configuration for EDN, CSRNG or the entropy source. At the start of a new
  // OTBN run, RND data is thus always invalidated and outstanding prefetches are marked such that
  // the RND data returned for the first prefetch is thrown away. When throwing away data, we need
  // to keep requesting RND data from EDN if another request got queued in the meantime.
  assign edn_rnd_req_start = (rnd_prefetch_req_i | rnd_req_i | rnd_req_queued_q) & ~rnd_valid_q;

  // When seeing a wipe with an outstanding request (which must have been a prefetch), we are going
  // to ignore the RND data that comes back from that request. Any RND data returned clears the
  // ignore status.
  assign edn_rnd_data_ignore_d =
      opn_start_i && edn_rnd_req_q ? 1'b1 :
      edn_rnd_req_complete         ? 1'b0 : edn_rnd_data_ignore_q;

  // rnd_req_queued_q shows that there's an outstanding RND prefetch whose result we are going to
  // ignore and also another request pending. Once the prefetch is done, we want to send out that
  // second request.
  //
  // The signal is set if we get a request (edn_rnd_req_start) when we're ignoring the current
  // prefetch (edn_rnd_data_ignore_q). It should be cleared when we actually start a request when
  // we're not ignoring a prefetch. It should also be cleared when finishing an operation. If that
  // happens, we were waiting to send a second prefetch and it turns out that no-one actually needed
  // the result.
  assign rnd_req_queued_d =
      opn_end_i             ? 1'b0              :
      edn_rnd_data_ignore_q ? edn_rnd_req_start :
      edn_rnd_req_start     ? 1'b0              : rnd_req_queued_q;

  // Assert `edn_rnd_req_o` when a request is started and keep it asserted until the request is
  // done.
  assign edn_rnd_req_d = (edn_rnd_req_q | edn_rnd_req_start) & ~edn_rnd_req_complete;

  assign edn_rnd_req_o = edn_rnd_req_q;

  always_ff @(posedge clk_i) begin
    if (rnd_data_en) begin
      rnd_data_q <= rnd_data_d;
      rnd_fips_q <= rnd_fips_d;
      rnd_err_q  <= rnd_err_d;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rnd_valid_q            <= 1'b0;
      rnd_req_queued_q       <= 1'b0;
      edn_rnd_req_q          <= 1'b0;
      edn_rnd_data_ignore_q  <= 1'b0;
    end else begin
      rnd_valid_q            <= rnd_valid_d;
      rnd_req_queued_q       <= rnd_req_queued_d;
      edn_rnd_req_q          <= edn_rnd_req_d;
      edn_rnd_data_ignore_q  <= edn_rnd_data_ignore_d;
    end
  end

  assign rnd_valid_o = rnd_valid_q;
  assign rnd_data_o  = rnd_data_q;

  // SEC_CM: RND.BUS.CONSISTENCY
  // SEC_CM: RND.RNG.DIGEST
  // Detect and forward RND error conditions.
  assign rnd_rep_err_o = rnd_req_complete & rnd_err_q;
  assign rnd_fips_err_o = rnd_req_complete & ~rnd_fips_q;

  /////////////////////////
  // PRNG Implementation //
  /////////////////////////

  logic edn_urnd_req_complete;
  logic edn_urnd_req_q, edn_urnd_req_d;

  assign edn_urnd_req_complete = edn_urnd_req_o & edn_urnd_ack_i;

  // Keep EDN URND request high even if input URND reseed request goes low before the reseed has
  // completed.
  assign edn_urnd_req_d = (edn_urnd_req_q | urnd_reseed_req_i) & ~edn_urnd_req_complete;

  assign edn_urnd_req_o = edn_urnd_req_q;
  assign urnd_reseed_ack_o = edn_urnd_ack_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      edn_urnd_req_q <= 1'b0;
    end else begin
      edn_urnd_req_q <= edn_urnd_req_d;
    end
  end

  logic xoshiro_seed_en;

  assign xoshiro_seed_en = edn_urnd_req_complete;

  prim_xoshiro256pp #(
    .OutputDw   (WLEN),
    .DefaultSeed(RndCnstUrndPrngSeed)
  ) u_xoshiro256pp(
    .clk_i,
    .rst_ni,
    .seed_en_i    (xoshiro_seed_en),
    .seed_i       (edn_urnd_data_i),
    .xoshiro_en_i (urnd_advance_i),
    .entropy_i    ('0),
    .data_o       (urnd_data_o),
    .all_zero_o   (urnd_all_zero_o)
  );

  `ASSERT(rnd_clear_on_req_complete, rnd_req_complete |=> ~rnd_valid_q)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * State machine to handle actions that occur around the start and stop of OTBN.
 *
 * This recieves the start signals from the top-level and passes them on to the
 * controller to begin execution when pre-start actions have finished.
 *
 * pre-start actions:
 *  - Seed LFSR for URND
 *
 * post-stop actions:
 *  - Internal Secure Wipe
 *    -Delete WDRs
 *    -Delete Base registers
 *    -Delete Accumulator
 *    -Delete Modulus
 *    -Reset stack
 */

`include "prim_assert.sv"

module otbn_start_stop_control
  import otbn_pkg::*;
  import prim_mubi_pkg::*;
#(
  // Disable URND advance when not in use. Useful for SCA only.
  parameter bit SecMuteUrnd = 1'b0,
  // Skip URND re-seed at the start of the operation. Useful for SCA only.
  parameter bit SecSkipUrndReseedAtStart = 1'b0
) (
  input  logic clk_i,
  input  logic rst_ni,

  input  logic   start_i,
  input  mubi4_t escalate_en_i,
  input  mubi4_t rma_req_i,
  output mubi4_t rma_ack_o,

  output logic controller_start_o,

  output logic urnd_reseed_req_o,
  input  logic urnd_reseed_ack_i,
  output logic urnd_reseed_err_o,
  output logic urnd_advance_o,

  input   logic secure_wipe_req_i,
  output  logic secure_wipe_ack_o,
  output  logic secure_wipe_running_o,
  output  logic done_o,

  output logic       sec_wipe_wdr_o,
  output logic       sec_wipe_wdr_urnd_o,
  output logic       sec_wipe_base_o,
  output logic       sec_wipe_base_urnd_o,
  output logic [4:0] sec_wipe_addr_o,

  output logic sec_wipe_acc_urnd_o,
  output logic sec_wipe_mod_urnd_o,
  output logic sec_wipe_zero_o,

  output logic ispr_init_o,
  output logic state_reset_o,
  output logic fatal_error_o
);

  import otbn_pkg::*;

  // Create lint errors to reduce the risk of accidentally enabling these features.
  `ASSERT_STATIC_LINT_ERROR(OtbnSecMuteUrndNonDefault, SecMuteUrnd == 0)
  `ASSERT_STATIC_LINT_ERROR(OtbnSecSkipUrndReseedAtStartNonDefault, SecSkipUrndReseedAtStart == 0)

  otbn_start_stop_state_e state_q, state_d;
  logic init_sec_wipe_done_q, init_sec_wipe_done_d;
  mubi4_t wipe_after_urnd_refresh_q, wipe_after_urnd_refresh_d;
  mubi4_t rma_ack_d, rma_ack_q;
  logic state_error_q, state_error_d;
  logic mubi_err_q, mubi_err_d;
  logic urnd_reseed_err_q, urnd_reseed_err_d;
  logic secure_wipe_error_q, secure_wipe_error_d;
  logic skip_reseed_q;

  logic addr_cnt_inc;
  logic [5:0] addr_cnt_q, addr_cnt_d;

  logic spurious_urnd_ack_error;
  logic spurious_secure_wipe_req, dropped_secure_wipe_req;

  // There are three ways in which the start/stop controller can be told to stop.
  // 1. secure_wipe_req_i comes from the controller (which means "I've run some instructions and
  //    I've hit an ECALL or error").
  // 2. escalate_en_i can be asserted (which means "Someone else has told us to stop immediately").
  // 3. rma_req_i can be asserted (which means "Lifecycle wants to transition to the RMA state").
  // If running, all three can be true at once.
  //
  // An escalation signal as well as RMA requests get latched into should_lock. We'll then go
  // through the secure wipe process (unless we weren't running any instructions in case of an
  // escalation). We'll see the should_lock_q signal when done and go into the local locked
  // state. If necessary, the RMA request is acknowledged upon secure wipe completion.

  // SEC_CM: CONTROLLER.FSM.GLOBAL_ESC
  logic esc_request, rma_request, should_lock_d, should_lock_q, stop;
  assign esc_request   = mubi4_test_true_loose(escalate_en_i);
  assign rma_request   = mubi4_test_true_strict(rma_req_i);
  assign stop          = esc_request | rma_request | secure_wipe_req_i;
  assign should_lock_d = should_lock_q | esc_request | rma_request;

  // Only if SecSkipUrndReseedAtStart is set, the controller start pulse is sent
  // one cycle after leaving the Halt state.
  if (SecSkipUrndReseedAtStart) begin: gen_skip_reseed
    logic skip_reseed_d;

    assign skip_reseed_d = ((state_q == OtbnStartStopStateHalt) & start_i & ~stop);

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        skip_reseed_q <= 1'b0;
      end else begin
        skip_reseed_q <= skip_reseed_d;
      end
    end
  end else begin: gen_reseed
    assign skip_reseed_q = 1'b0;
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      should_lock_q <= 1'b0;
    end else begin
      should_lock_q <= should_lock_d;
    end
  end

  prim_mubi4_sender #(
    .AsyncOn(1'b1),
    .EnSecBuf(1'b1),
    .ResetValue(prim_mubi_pkg::MuBi4False)
  ) u_prim_mubi4_sender_rma_ack (
    .clk_i,
    .rst_ni,
    .mubi_i(rma_ack_d),
    .mubi_o(rma_ack_q)
  );

  logic allow_secure_wipe, expect_secure_wipe;

  // SEC_CM: START_STOP_CTRL.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q,
      otbn_start_stop_state_e, OtbnStartStopStateInitial)

  always_comb begin
    urnd_reseed_req_o         = 1'b0;
    urnd_advance_o            = 1'b0;
    state_d                   = state_q;
    ispr_init_o               = 1'b0;
    state_reset_o             = 1'b0;
    sec_wipe_wdr_o            = 1'b0;
    sec_wipe_wdr_urnd_o       = 1'b0;
    sec_wipe_base_o           = 1'b0;
    sec_wipe_base_urnd_o      = 1'b0;
    sec_wipe_acc_urnd_o       = 1'b0;
    sec_wipe_mod_urnd_o       = 1'b0;
    sec_wipe_zero_o           = 1'b0;
    addr_cnt_inc              = 1'b0;
    secure_wipe_ack_o         = 1'b0;
    secure_wipe_running_o     = 1'b0;
    state_error_d             = state_error_q;
    allow_secure_wipe         = 1'b0;
    expect_secure_wipe        = 1'b0;
    spurious_urnd_ack_error   = 1'b0;
    wipe_after_urnd_refresh_d = wipe_after_urnd_refresh_q;
    rma_ack_d                 = rma_ack_q;
    mubi_err_d                = mubi_err_q;

    unique case (state_q)
      OtbnStartStopStateInitial: begin
        secure_wipe_running_o = 1'b1;
        urnd_reseed_req_o     = 1'b1;
        if (rma_request) begin
          // If we get an RMA request before the URND got reseeded, proceed with the initial secure
          // wipe, as the entropy complex may not be able to provide entropy at this point.
          state_d = OtbnStartStopSecureWipeWdrUrnd;
          // As we don't reseed URND, there's no point in doing two rounds of wiping, so we pretend
          // that the first round is already the second round.
          wipe_after_urnd_refresh_d = MuBi4True;
        end else if (urnd_reseed_ack_i) begin
          urnd_advance_o = 1'b1;
          state_d        = OtbnStartStopSecureWipeWdrUrnd;
        end
      end
      OtbnStartStopStateHalt: begin
        if (stop && !rma_request) begin
          state_d = OtbnStartStopStateLocked;
        end else if (start_i || rma_request) begin
          ispr_init_o   = 1'b1;
          state_reset_o = 1'b1;
          if (rma_request) begin
            // Do not reseed URND before secure wipe for RMA, as the entropy complex may not be able
            // to provide entropy at this point.
            state_d = OtbnStartStopSecureWipeWdrUrnd;
            // As we don't reseed URND, there's no point in doing two rounds of wiping, so we
            // pretend that the first round is already the second round.
            wipe_after_urnd_refresh_d = MuBi4True;
          end else begin // start_i
            urnd_reseed_req_o = ~SecSkipUrndReseedAtStart;
            state_d           = OtbnStartStopStateUrndRefresh;
          end
        end
      end
      OtbnStartStopStateUrndRefresh: begin
        urnd_reseed_req_o = ~skip_reseed_q;
        if (stop) begin
          if (mubi4_test_false_strict(wipe_after_urnd_refresh_q)) begin
            // We are told to stop and don't have to wipe after the current URND refresh is ack'd,
            // so we lock immediately.
            state_d = OtbnStartStopStateLocked;
          end else begin
            // We are told to stop but should wipe after the current URND refresh is ack'd, so we
            // wait for the ACK and then do a secure wipe.
            allow_secure_wipe     = 1'b1;
            expect_secure_wipe    = 1'b1;
            secure_wipe_running_o = 1'b1;
            if (urnd_reseed_ack_i) begin
              state_d = OtbnStartStopSecureWipeWdrUrnd;
            end
          end
        end else begin
          if (mubi4_test_false_strict(wipe_after_urnd_refresh_q)) begin
            // We are not stopping and we don't have to wipe after the current URND refresh is
            // ack'd, so we wait for the ACK and then start executing.
            if (urnd_reseed_ack_i || skip_reseed_q) begin
              state_d = OtbnStartStopStateRunning;
            end
          end else begin
            // We are not stopping but should wipe after the current URND refresh is ack'd, so we
            // wait for the ACK and then do a secure wipe.
            allow_secure_wipe     = 1'b1;
            expect_secure_wipe    = 1'b1;
            secure_wipe_running_o = 1'b1;
            if (urnd_reseed_ack_i) begin
              state_d = OtbnStartStopSecureWipeWdrUrnd;
            end
          end
        end
      end
      OtbnStartStopStateRunning: begin
        urnd_advance_o    = ~SecMuteUrnd;
        allow_secure_wipe = 1'b1;

        if (stop) begin
          state_d = OtbnStartStopSecureWipeWdrUrnd;
        end
      end
      // SEC_CM: DATA_REG_SW.SEC_WIPE
      // Writing random numbers to the wide data registers.
       OtbnStartStopSecureWipeWdrUrnd: begin
        urnd_advance_o        = 1'b1;
        addr_cnt_inc          = 1'b1;
        sec_wipe_wdr_o        = 1'b1;
        sec_wipe_wdr_urnd_o   = 1'b1;
        allow_secure_wipe     = 1'b1;
        expect_secure_wipe    = 1'b1;
        secure_wipe_running_o = 1'b1;

        // Count one extra cycle when wiping the WDR, because the wipe signals to the WDR
        // (`sec_wipe_wdr_o` and `sec_wipe_wdr_urnd_o`) are flopped once but the wipe signals to the
        // ACC register, which is wiped directly after the last WDR, are not.  If we would not count
        // this extra cycle, the last WDR and the ACC register would be wiped simultaneously and
        // thus with the same random value.
        if (addr_cnt_q == 6'b100000) begin
          // Reset `addr_cnt` on the transition out of this state.
          addr_cnt_inc = 1'b0;
          // The following two signals are flopped once before they reach the FSM, so clear them one
          // cycle early here.
          sec_wipe_wdr_o      = 1'b0;
          sec_wipe_wdr_urnd_o = 1'b0;
          state_d = OtbnStartStopSecureWipeAccModBaseUrnd;
        end
      end
      // Writing random numbers to the accumulator, modulus and the base registers.
      // addr_cnt_q wraps around to 0 when first moving to this state, and we need to
      // supress writes to the zero register and the call stack.
       OtbnStartStopSecureWipeAccModBaseUrnd: begin
        urnd_advance_o        = 1'b1;
        addr_cnt_inc          = 1'b1;
        allow_secure_wipe     = 1'b1;
        expect_secure_wipe    = 1'b1;
        secure_wipe_running_o = 1'b1;
        // The first two clock cycles are used to write random data to accumulator and modulus.
        sec_wipe_acc_urnd_o   = (addr_cnt_q == 6'b000000);
        sec_wipe_mod_urnd_o   = (addr_cnt_q == 6'b000001);
        // Supress writes to the zero register and the call stack.
        sec_wipe_base_o       = (addr_cnt_q > 6'b000001);
        sec_wipe_base_urnd_o  = (addr_cnt_q > 6'b000001);
        if (addr_cnt_q == 6'b011111) begin
          state_d = OtbnStartStopSecureWipeAllZero;
        end
      end
      // Writing zeros to the CSRs and reset the stack. The other registers are intentionally not
      // overwritten with zero.
       OtbnStartStopSecureWipeAllZero: begin
        sec_wipe_zero_o       = 1'b1;
        allow_secure_wipe     = 1'b1;
        expect_secure_wipe    = 1'b1;
        secure_wipe_running_o = 1'b1;

        // Leave this state after a single cycle, which is sufficient to reset the CSRs and the
        // stack.
        if (mubi4_test_false_strict(wipe_after_urnd_refresh_q)) begin
          // This is the first round of wiping with random numbers, refresh URND and do a second
          // round.
          state_d = OtbnStartStopStateUrndRefresh;
          wipe_after_urnd_refresh_d = MuBi4True;
        end else begin
          // This is the second round of wiping with random numbers, so the secure wipe is
          // complete.
          state_d = OtbnStartStopSecureWipeComplete;
          secure_wipe_ack_o = 1'b1;
        end
      end
      OtbnStartStopSecureWipeComplete: begin
        urnd_advance_o = 1'b1;
        rma_ack_d = rma_req_i;
        state_d = should_lock_d ? OtbnStartStopStateLocked : OtbnStartStopStateHalt;
        wipe_after_urnd_refresh_d = MuBi4False;
      end
      OtbnStartStopStateLocked: begin
        // SEC_CM: START_STOP_CTRL.FSM.GLOBAL_ESC
        // SEC_CM: START_STOP_CTRL.FSM.LOCAL_ESC
        //
        // Terminal state. This is either accessed by glitching state_q (and going through the
        // default case below) or by getting an escalation signal
      end
      default: begin
        // We should never get here. If we do (e.g. via a malicious glitch), error out immediately.
        state_error_d = 1'b1;
        rma_ack_d = MuBi4False;
        state_d = OtbnStartStopStateLocked;
      end
    endcase

    if (urnd_reseed_ack_i &&
        !(state_q inside {OtbnStartStopStateInitial, OtbnStartStopStateUrndRefresh})) begin
      // We should never receive an ACK from URND when we're not refreshing the URND. Signal an
      // error if we see a stray ACK and lock the FSM.
      spurious_urnd_ack_error = 1'b1;
      state_d                 = OtbnStartStopStateLocked;
    end

    // If the MuBi signals take on invalid values, something bad is happening. Put them back to
    // a safe value (if possible) and signal an error.
    if (mubi4_test_invalid(escalate_en_i)) begin
      mubi_err_d = 1'b1;
      state_d = OtbnStartStopStateLocked;
    end
    if (mubi4_test_invalid(rma_req_i)) begin
      mubi_err_d = 1'b1;
      state_d = OtbnStartStopStateLocked;
    end
    if (mubi4_test_invalid(wipe_after_urnd_refresh_q)) begin
      wipe_after_urnd_refresh_d = MuBi4False;
      mubi_err_d = 1'b1;
      state_d = OtbnStartStopStateLocked;
    end
    if (mubi4_test_invalid(rma_ack_q)) begin
      rma_ack_d = MuBi4False;
      mubi_err_d = 1'b1;
      state_d = OtbnStartStopStateLocked;
    end
  end

  // Latch initial secure wipe done.
  assign init_sec_wipe_done_d = (state_q == OtbnStartStopSecureWipeComplete) ? 1'b1 : // set
                                init_sec_wipe_done_q; // keep

  // Logic separate from main FSM code to avoid false combinational loop warning from verilator
  assign controller_start_o =
    // The controller start pulse is fired when finishing the initial URND reseed.
    ((state_q == OtbnStartStopStateUrndRefresh) & (urnd_reseed_ack_i | skip_reseed_q) &
      mubi4_test_false_strict(wipe_after_urnd_refresh_q));

  assign done_o = ((state_q == OtbnStartStopSecureWipeComplete && init_sec_wipe_done_q) ||
                   (stop && (state_q == OtbnStartStopStateUrndRefresh) &&
                    mubi4_test_false_strict(wipe_after_urnd_refresh_q)) ||
                   (spurious_urnd_ack_error && !(state_q inside {OtbnStartStopStateHalt,
                                                                 OtbnStartStopStateLocked}) &&
                    init_sec_wipe_done_q) || (mubi_err_d && !mubi_err_q));

  assign addr_cnt_d = addr_cnt_inc ? (addr_cnt_q + 6'd1) : 6'd0;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      addr_cnt_q           <= 6'd0;
      init_sec_wipe_done_q <= 1'b0;
    end else begin
      addr_cnt_q           <= addr_cnt_d;
      init_sec_wipe_done_q <= init_sec_wipe_done_d;
    end
  end

  prim_mubi4_sender #(
    .AsyncOn(1),
    .ResetValue(MuBi4False)
  ) u_wipe_after_urnd_refresh_flop (
    .clk_i,
    .rst_ni,
    .mubi_i(wipe_after_urnd_refresh_d),
    .mubi_o(wipe_after_urnd_refresh_q)
  );

  // Clip the secure wipe address to [0..31].  This is safe because the wipe enable signals are
  // never set when the counter exceeds 5 bit, which we assert below.
  assign sec_wipe_addr_o = addr_cnt_q[4:0];
  `ASSERT(NoSecWipeAbove32Bit_A, addr_cnt_q[5] |-> (!sec_wipe_wdr_o && !sec_wipe_acc_urnd_o))

  // A check for spurious or dropped secure wipe requests.
  // We only expect to start a secure wipe when running.
  assign spurious_secure_wipe_req = secure_wipe_req_i & ~allow_secure_wipe;
  // Once we've started a secure wipe, the controller should not drop the request until we tell it
  // we're done. This does not apply for the *initial* secure wipe, though, which is controlled by
  // this module rather than the controller.
  assign dropped_secure_wipe_req  = expect_secure_wipe & init_sec_wipe_done_d & ~secure_wipe_req_i;

  // Delay the "glitch req/ack" error signal by a cycle. Otherwise, you end up with a combinatorial
  // loop through the escalation signal that our fatal_error_o causes otbn_core to pass to the
  // controller.
  assign secure_wipe_error_d = spurious_secure_wipe_req | dropped_secure_wipe_req;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      state_error_q       <= 1'b0;
      mubi_err_q          <= 1'b0;
      secure_wipe_error_q <= 1'b0;
      urnd_reseed_err_q   <= 1'b0;
    end else begin
      state_error_q       <= state_error_d;
      mubi_err_q          <= mubi_err_d;
      secure_wipe_error_q <= secure_wipe_error_d;
      urnd_reseed_err_q   <= urnd_reseed_err_d;
    end
  end

  assign urnd_reseed_err_d = spurious_urnd_ack_error ? 1'b1 // set
                                                     : urnd_reseed_err_q; // hold
  assign urnd_reseed_err_o = urnd_reseed_err_d;

  assign fatal_error_o = urnd_reseed_err_o | state_error_d | secure_wipe_error_q | mubi_err_q;

  assign rma_ack_o = rma_ack_q;

  `ASSERT(StartStopStateValid_A,
      state_q inside {OtbnStartStopStateInitial,
                      OtbnStartStopStateHalt,
                      OtbnStartStopStateUrndRefresh,
                      OtbnStartStopStateRunning,
                      OtbnStartStopSecureWipeWdrUrnd,
                      OtbnStartStopSecureWipeAccModBaseUrnd,
                      OtbnStartStopSecureWipeAllZero,
                      OtbnStartStopSecureWipeComplete,
                      OtbnStartStopStateLocked})

  `ASSERT(StartSecureWipeImpliesRunning_A,
          $rose(secure_wipe_req_i) |-> (state_q == OtbnStartStopStateRunning))

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OpenTitan Big Number Accelerator (OTBN) Core
 *
 * This module is the top-level of the OTBN processing core.
 */
// Below countermeasure (no data dependent control flow in OTBN ISA) is inherent to the design and
// has no directly associated RTL
// SEC_CM: CTRL_FLOW.SCA
module otbn_core
  import otbn_pkg::*;
#(
  // Register file implementation selection, see otbn_pkg.sv.
  parameter regfile_e RegFile = RegFileFF,

  // Size of the instruction memory, in bytes
  parameter int ImemSizeByte = 4096,
  // Size of the data memory, in bytes
  parameter int DmemSizeByte = 4096,

  // Default seed for URND PRNG
  parameter urnd_prng_seed_t RndCnstUrndPrngSeed = RndCnstUrndPrngSeedDefault,

  // Disable URND reseed and advance when not in use. Useful for SCA only.
  parameter bit SecMuteUrnd = 1'b0,
  parameter bit SecSkipUrndReseedAtStart = 1'b0,

  localparam int ImemAddrWidth = prim_util_pkg::vbits(ImemSizeByte),
  localparam int DmemAddrWidth = prim_util_pkg::vbits(DmemSizeByte)
) (
  input logic clk_i,
  input logic rst_ni,

  input  logic start_i,   // start the operation
  output logic done_o,    // operation done
  output logic locking_o, // The core is in or is entering the locked state
  output logic secure_wipe_running_o, // the core is securely wiping its internal state

  output core_err_bits_t err_bits_o,  // valid when done_o is asserted
  output logic           recoverable_err_o,

  // Instruction memory (IMEM)
  output logic                     imem_req_o,
  output logic [ImemAddrWidth-1:0] imem_addr_o,
  input  logic [38:0]              imem_rdata_i,
  input  logic                     imem_rvalid_i,

  // Data memory (DMEM)
  output logic                        dmem_req_o,
  output logic                        dmem_write_o,
  output logic [DmemAddrWidth-1:0]    dmem_addr_o,
  output logic [ExtWLEN-1:0]          dmem_wdata_o,
  output logic [ExtWLEN-1:0]          dmem_wmask_o,
  output logic [BaseWordsPerWLEN-1:0] dmem_rmask_o,
  input  logic [ExtWLEN-1:0]          dmem_rdata_i,
  input  logic                        dmem_rvalid_i,
  input  logic                        dmem_rerror_i,

  // Entropy distribution network (EDN) connections
  // One for RND, the other for URND
  output logic                    edn_rnd_req_o,
  input  logic                    edn_rnd_ack_i,
  input  logic [EdnDataWidth-1:0] edn_rnd_data_i,
  input  logic                    edn_rnd_fips_i,
  input  logic                    edn_rnd_err_i,

  output logic                    edn_urnd_req_o,
  input  logic                    edn_urnd_ack_i,
  input  logic [EdnDataWidth-1:0] edn_urnd_data_i,

  output logic [31:0] insn_cnt_o,
  input  logic        insn_cnt_clear_i,

  output logic         mems_sec_wipe_o,          // Request secure wipe for imem and dmem
  input  logic         req_sec_wipe_urnd_keys_i, // Request URND bits for temporary scramble keys.
                                                 // Keys below are valid cycle after request.
  output logic [127:0] dmem_sec_wipe_urnd_key_o, // URND bits to give temporary dmem scramble key
  output logic [127:0] imem_sec_wipe_urnd_key_o, // URND bits to give temporary imem scramble key

  // Indicates an incoming escalation from some fatal error at the level above. The core needs to
  // halt and then enter a locked state.
  input prim_mubi_pkg::mubi4_t escalate_en_i,

  // Indicates an incoming RMA request. The core needs to halt, trigger a secure wipe immediately
  // and then enter a locked state.
  input  prim_mubi_pkg::mubi4_t rma_req_i,
  output prim_mubi_pkg::mubi4_t rma_ack_o,

  // When set software errors become fatal errors.
  input logic software_errs_fatal_i,

  input logic [1:0]                       sideload_key_shares_valid_i,
  input logic [1:0][SideloadKeyWidth-1:0] sideload_key_shares_i
);
  import prim_mubi_pkg::*;

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(OtbnSecMuteUrndNonDefault, SecMuteUrnd == 0)

  // Fetch request (the next instruction)
  logic [ImemAddrWidth-1:0] insn_fetch_req_addr;
  logic                     insn_fetch_req_valid;
  logic                     insn_fetch_req_valid_raw;

  // Fetch response (the current instruction before it is decoded)
  logic                     insn_fetch_resp_valid;
  logic [ImemAddrWidth-1:0] insn_fetch_resp_addr;
  logic [31:0]              insn_fetch_resp_data;
  logic                     insn_fetch_resp_clear;
  logic                     insn_fetch_err;
  logic                     insn_addr_err;

  rf_predec_bignum_t        rf_predec_bignum;
  alu_predec_bignum_t       alu_predec_bignum;
  ctrl_flow_predec_t        ctrl_flow_predec;
  logic [ImemAddrWidth-1:0] ctrl_flow_target_predec;
  ispr_predec_bignum_t      ispr_predec_bignum;
  mac_predec_bignum_t       mac_predec_bignum;
  logic                     lsu_addr_en_predec;

  logic [NWdr-1:0] rf_bignum_rd_a_indirect_onehot;
  logic [NWdr-1:0] rf_bignum_rd_b_indirect_onehot;
  logic [NWdr-1:0] rf_bignum_wr_indirect_onehot;
  logic            rf_bignum_indirect_en;

  // The currently executed instruction.
  logic                     insn_valid;
  logic                     insn_illegal;
  logic [ImemAddrWidth-1:0] insn_addr;
  insn_dec_base_t           insn_dec_base;
  insn_dec_bignum_t         insn_dec_bignum;
  insn_dec_shared_t         insn_dec_shared;

  logic [4:0]               rf_base_wr_addr;
  logic [4:0]               rf_base_wr_addr_ctrl;
  logic                     rf_base_wr_en;
  logic                     rf_base_wr_en_ctrl;
  logic                     rf_base_wr_commit;
  logic                     rf_base_wr_commit_ctrl;
  logic [31:0]              rf_base_wr_data_no_intg;
  logic [31:0]              rf_base_wr_data_no_intg_ctrl;
  logic [BaseIntgWidth-1:0] rf_base_wr_data_intg;
  logic                     rf_base_wr_data_intg_sel, rf_base_wr_data_intg_sel_ctrl;
  logic [4:0]               rf_base_rd_addr_a;
  logic                     rf_base_rd_en_a;
  logic [BaseIntgWidth-1:0] rf_base_rd_data_a_intg;
  logic [4:0]               rf_base_rd_addr_b;
  logic                     rf_base_rd_en_b;
  logic [BaseIntgWidth-1:0] rf_base_rd_data_b_intg;
  logic                     rf_base_rd_commit;
  logic                     rf_base_call_stack_sw_err;
  logic                     rf_base_call_stack_hw_err;
  logic                     rf_base_intg_err;
  logic                     rf_base_spurious_we_err;

  alu_base_operation_t  alu_base_operation;
  alu_base_comparison_t alu_base_comparison;
  logic [31:0]          alu_base_operation_result;
  logic                 alu_base_comparison_result;

  logic                     lsu_load_req;
  logic                     lsu_store_req;
  insn_subset_e             lsu_req_subset;
  logic [DmemAddrWidth-1:0] lsu_addr;

  logic [BaseIntgWidth-1:0] lsu_base_wdata;
  logic [ExtWLEN-1:0]       lsu_bignum_wdata;

  logic [BaseIntgWidth-1:0] lsu_base_rdata;
  logic [ExtWLEN-1:0]       lsu_bignum_rdata;
  logic                     lsu_rdata_err;

  logic [WdrAw-1:0]   rf_bignum_wr_addr;
  logic [WdrAw-1:0]   rf_bignum_wr_addr_ctrl;
  logic [1:0]         rf_bignum_wr_en;
  logic [1:0]         rf_bignum_wr_en_ctrl;
  logic               rf_bignum_wr_commit;
  logic               rf_bignum_wr_commit_ctrl;
  logic [WLEN-1:0]    rf_bignum_wr_data_no_intg;
  logic [WLEN-1:0]    rf_bignum_wr_data_no_intg_ctrl;
  logic [ExtWLEN-1:0] rf_bignum_wr_data_intg;
  logic               rf_bignum_wr_data_intg_sel, rf_bignum_wr_data_intg_sel_ctrl;
  logic [WdrAw-1:0]   rf_bignum_rd_addr_a;
  logic               rf_bignum_rd_en_a;
  logic [ExtWLEN-1:0] rf_bignum_rd_data_a_intg;
  logic [WdrAw-1:0]   rf_bignum_rd_addr_b;
  logic               rf_bignum_rd_en_b;
  logic [ExtWLEN-1:0] rf_bignum_rd_data_b_intg;
  logic               rf_bignum_intg_err;
  logic               rf_bignum_spurious_we_err;

  alu_bignum_operation_t alu_bignum_operation;
  logic                  alu_bignum_operation_valid;
  logic                  alu_bignum_operation_commit;
  logic [WLEN-1:0]       alu_bignum_operation_result;
  logic                  alu_bignum_selection_flag;
  logic                  alu_bignum_reg_intg_violation_err;

  mac_bignum_operation_t mac_bignum_operation;
  logic [WLEN-1:0]       mac_bignum_operation_result;
  flags_t                mac_bignum_operation_flags;
  flags_t                mac_bignum_operation_flags_en;
  logic                  mac_bignum_en;
  logic                  mac_bignum_commit;
  logic                  mac_bignum_reg_intg_violation_err;

  ispr_e                       ispr_addr;
  logic [31:0]                 ispr_base_wdata;
  logic [BaseWordsPerWLEN-1:0] ispr_base_wr_en;
  logic [ExtWLEN-1:0]          ispr_bignum_wdata_intg;
  logic                        ispr_bignum_wr_en;
  logic [NFlagGroups-1:0]      ispr_flags_wr;
  logic                        ispr_wr_commit;
  logic [ExtWLEN-1:0]          ispr_rdata_intg;
  logic                        ispr_rd_en;
  logic [ExtWLEN-1:0]          ispr_acc_intg;
  logic [ExtWLEN-1:0]          ispr_acc_wr_data_intg;
  logic                        ispr_acc_wr_en;
  logic                        ispr_init;

  logic            rnd_req;
  logic            rnd_prefetch_req;
  logic            rnd_valid;
  logic [WLEN-1:0] rnd_data;
  logic            rnd_rep_err;
  logic            rnd_fips_err;

  logic            urnd_reseed_req;
  logic            urnd_reseed_ack;
  logic            urnd_reseed_err;
  logic            urnd_advance;
  logic            urnd_advance_start_stop_control;
  logic [WLEN-1:0] urnd_data;
  logic            urnd_all_zero;

  logic        controller_start;

  logic        state_reset;
  logic [31:0] insn_cnt;

  logic secure_wipe_req, secure_wipe_ack;

  logic sec_wipe_wdr_d, sec_wipe_wdr_q;
  logic sec_wipe_wdr_urnd_d, sec_wipe_wdr_urnd_q;
  logic sec_wipe_base;
  logic sec_wipe_base_urnd;
  logic [4:0] sec_wipe_addr, sec_wipe_wdr_addr_q;

  logic sec_wipe_acc_urnd;
  logic sec_wipe_mod_urnd;
  logic sec_wipe_zero;

  logic zero_flags;

  logic                     prefetch_en;
  logic                     prefetch_loop_active;
  logic [31:0]              prefetch_loop_iterations;
  logic [ImemAddrWidth:0]   prefetch_loop_end_addr;
  logic [ImemAddrWidth-1:0] prefetch_loop_jump_addr;

  mubi4_t               controller_fatal_escalate_en, controller_recov_escalate_en;
  mubi4_t               start_stop_escalate_en;
  controller_err_bits_t controller_err_bits;
  logic                 prefetch_ignore_errs;

  core_err_bits_t err_bits_q, err_bits_d;
  logic           mubi_err;

  logic start_stop_fatal_error;
  logic rf_bignum_predec_error, alu_bignum_predec_error, ispr_predec_error, mac_bignum_predec_error;
  logic controller_predec_error;
  logic rd_predec_error, predec_error;

  logic req_sec_wipe_urnd_keys_q;

  // Start stop control start OTBN execution when requested and deals with any pre start or post
  // stop actions.
  otbn_start_stop_control #(
    .SecMuteUrnd(SecMuteUrnd),
    .SecSkipUrndReseedAtStart(SecSkipUrndReseedAtStart)
  ) u_otbn_start_stop_control (
    .clk_i,
    .rst_ni,

    .start_i,
    .escalate_en_i(start_stop_escalate_en),
    .rma_req_i,
    .rma_ack_o,

    .controller_start_o(controller_start),

    .urnd_reseed_req_o (urnd_reseed_req),
    .urnd_reseed_ack_i (urnd_reseed_ack),
    .urnd_reseed_err_o (urnd_reseed_err),
    .urnd_advance_o    (urnd_advance_start_stop_control),

    .secure_wipe_req_i (secure_wipe_req),
    .secure_wipe_ack_o (secure_wipe_ack),
    .secure_wipe_running_o,
    .done_o,

    .sec_wipe_wdr_o      (sec_wipe_wdr_d),
    .sec_wipe_wdr_urnd_o (sec_wipe_wdr_urnd_d),
    .sec_wipe_base_o     (sec_wipe_base),
    .sec_wipe_base_urnd_o(sec_wipe_base_urnd),
    .sec_wipe_addr_o     (sec_wipe_addr),

    .sec_wipe_acc_urnd_o(sec_wipe_acc_urnd),
    .sec_wipe_mod_urnd_o(sec_wipe_mod_urnd),
    .sec_wipe_zero_o    (sec_wipe_zero),

    .ispr_init_o  (ispr_init),
    .state_reset_o(state_reset),
    .fatal_error_o(start_stop_fatal_error)
  );

  // Depending on its usage, the instruction address (program counter) is qualified by two valid
  // signals: insn_fetch_resp_valid (together with the undecoded instruction data), and insn_valid
  // for valid decoded (i.e. legal) instructions. Duplicate the signal in the source code for
  // consistent grouping of signals with their valid signal.
  assign insn_addr = insn_fetch_resp_addr;

  // For secure wipe and ISPR initialization, flags need to be cleared to 0. This is achieved
  // through the blanking mechanism controlled by the instruction fetch/predecoder stage.
  assign zero_flags = sec_wipe_zero | ispr_init;

  // Instruction fetch unit
  otbn_instruction_fetch #(
    .ImemSizeByte(ImemSizeByte)
  ) u_otbn_instruction_fetch (
    .clk_i,
    .rst_ni,

    // Instruction memory interface
    .imem_req_o,
    .imem_addr_o,
    .imem_rdata_i,
    .imem_rvalid_i,

    // Instruction to fetch
    .insn_fetch_req_addr_i     (insn_fetch_req_addr),
    .insn_fetch_req_valid_i    (insn_fetch_req_valid),
    .insn_fetch_req_valid_raw_i(insn_fetch_req_valid_raw),

    // Fetched instruction
    .insn_fetch_resp_addr_o (insn_fetch_resp_addr),
    .insn_fetch_resp_valid_o(insn_fetch_resp_valid),
    .insn_fetch_resp_data_o (insn_fetch_resp_data),
    .insn_fetch_resp_clear_i(insn_fetch_resp_clear),
    .insn_fetch_err_o       (insn_fetch_err),
    .insn_addr_err_o        (insn_addr_err),

    .rf_predec_bignum_o       (rf_predec_bignum),
    .alu_predec_bignum_o      (alu_predec_bignum),
    .ctrl_flow_predec_o       (ctrl_flow_predec),
    .ctrl_flow_target_predec_o(ctrl_flow_target_predec),
    .ispr_predec_bignum_o     (ispr_predec_bignum),
    .mac_predec_bignum_o      (mac_predec_bignum),
    .lsu_addr_en_predec_o     (lsu_addr_en_predec),

    .rf_bignum_rd_a_indirect_onehot_i(rf_bignum_rd_a_indirect_onehot),
    .rf_bignum_rd_b_indirect_onehot_i(rf_bignum_rd_b_indirect_onehot),
    .rf_bignum_wr_indirect_onehot_i  (rf_bignum_wr_indirect_onehot),
    .rf_bignum_indirect_en_i         (rf_bignum_indirect_en),

    .prefetch_en_i             (prefetch_en),
    .prefetch_loop_active_i    (prefetch_loop_active),
    .prefetch_loop_iterations_i(prefetch_loop_iterations),
    .prefetch_loop_end_addr_i  (prefetch_loop_end_addr),
    .prefetch_loop_jump_addr_i (prefetch_loop_jump_addr),
    .prefetch_ignore_errs_i    (prefetch_ignore_errs),

    .sec_wipe_wdr_en_i  (sec_wipe_wdr_d),
    .sec_wipe_wdr_addr_i(sec_wipe_addr),

    .zero_flags_i(zero_flags)
  );

  // Instruction decoder
  otbn_decoder u_otbn_decoder (
    // The decoder is combinatorial; clk and rst are only used for assertions.
    .clk_i,
    .rst_ni,

    // Instruction to decode
    .insn_fetch_resp_data_i (insn_fetch_resp_data),
    .insn_fetch_resp_valid_i(insn_fetch_resp_valid),

    // Decoded instruction
    .insn_valid_o     (insn_valid),
    .insn_illegal_o   (insn_illegal),
    .insn_dec_base_o  (insn_dec_base),
    .insn_dec_bignum_o(insn_dec_bignum),
    .insn_dec_shared_o(insn_dec_shared)
  );

  // SEC_CM: CTRL.REDUN
  // ALU and MAC predecode is only relevant when there is a valid instruction, as without one it is
  // guaranteed there are no register reads (hence no sensitive data bits being fed into the blanked
  // data paths). RF and ISPR predecode must always be checked to ensure read and write data paths
  // are always correctly blanked.
  assign rd_predec_error = |{rf_predec_bignum.rf_ren_a,
                             rf_predec_bignum.rf_ren_b,
                             ispr_predec_bignum.ispr_rd_en} & ~insn_valid;

  assign predec_error =
    ((alu_bignum_predec_error | mac_bignum_predec_error | controller_predec_error) & insn_valid) |
     rf_bignum_predec_error                                                                      |
     ispr_predec_error                                                                           |
     rd_predec_error;

  // Controller: coordinate between functional units, prepare their inputs (e.g. by muxing between
  // operand sources), and post-process their outputs as needed.
  otbn_controller #(
    .ImemSizeByte(ImemSizeByte),
    .DmemSizeByte(DmemSizeByte)
  ) u_otbn_controller (
    .clk_i,
    .rst_ni,

    .start_i         (controller_start),
    .locking_o,
    .err_bit_clear_i (start_i),

    .fatal_escalate_en_i(controller_fatal_escalate_en),
    .recov_escalate_en_i(controller_recov_escalate_en),
    .rma_req_i,
    .err_bits_o         (controller_err_bits),
    .recoverable_err_o,

    // Next instruction selection (to instruction fetch)
    .insn_fetch_req_addr_o     (insn_fetch_req_addr),
    .insn_fetch_req_valid_o    (insn_fetch_req_valid),
    .insn_fetch_req_valid_raw_o(insn_fetch_req_valid_raw),
    .insn_fetch_resp_clear_o   (insn_fetch_resp_clear),

    // The current instruction
    .insn_valid_i  (insn_valid),
    .insn_illegal_i(insn_illegal),
    .insn_addr_i   (insn_addr),

    // Decoded instruction from decoder
    .insn_dec_base_i  (insn_dec_base),
    .insn_dec_bignum_i(insn_dec_bignum),
    .insn_dec_shared_i(insn_dec_shared),

    // To/from base register file
    .rf_base_wr_addr_o          (rf_base_wr_addr_ctrl),
    .rf_base_wr_en_o            (rf_base_wr_en_ctrl),
    .rf_base_wr_commit_o        (rf_base_wr_commit_ctrl),
    .rf_base_wr_data_no_intg_o  (rf_base_wr_data_no_intg_ctrl),
    .rf_base_wr_data_intg_o     (rf_base_wr_data_intg),
    .rf_base_wr_data_intg_sel_o (rf_base_wr_data_intg_sel_ctrl),
    .rf_base_rd_addr_a_o        (rf_base_rd_addr_a),
    .rf_base_rd_en_a_o          (rf_base_rd_en_a),
    .rf_base_rd_data_a_intg_i   (rf_base_rd_data_a_intg),
    .rf_base_rd_addr_b_o        (rf_base_rd_addr_b),
    .rf_base_rd_en_b_o          (rf_base_rd_en_b),
    .rf_base_rd_data_b_intg_i   (rf_base_rd_data_b_intg),
    .rf_base_rd_commit_o        (rf_base_rd_commit),
    .rf_base_call_stack_sw_err_i(rf_base_call_stack_sw_err),
    .rf_base_call_stack_hw_err_i(rf_base_call_stack_hw_err),

    // To/from bignum register file
    .rf_bignum_wr_addr_o         (rf_bignum_wr_addr_ctrl),
    .rf_bignum_wr_en_o           (rf_bignum_wr_en_ctrl),
    .rf_bignum_wr_commit_o       (rf_bignum_wr_commit_ctrl),
    .rf_bignum_wr_data_no_intg_o (rf_bignum_wr_data_no_intg_ctrl),
    .rf_bignum_wr_data_intg_o    (rf_bignum_wr_data_intg),
    .rf_bignum_wr_data_intg_sel_o(rf_bignum_wr_data_intg_sel_ctrl),
    .rf_bignum_rd_addr_a_o       (rf_bignum_rd_addr_a),
    .rf_bignum_rd_en_a_o         (rf_bignum_rd_en_a),
    .rf_bignum_rd_data_a_intg_i  (rf_bignum_rd_data_a_intg),
    .rf_bignum_rd_addr_b_o       (rf_bignum_rd_addr_b),
    .rf_bignum_rd_en_b_o         (rf_bignum_rd_en_b),
    .rf_bignum_rd_data_b_intg_i  (rf_bignum_rd_data_b_intg),
    .rf_bignum_intg_err_i        (rf_bignum_intg_err),
    .rf_bignum_spurious_we_err_i (rf_bignum_spurious_we_err),

    .rf_bignum_rd_a_indirect_onehot_o(rf_bignum_rd_a_indirect_onehot),
    .rf_bignum_rd_b_indirect_onehot_o(rf_bignum_rd_b_indirect_onehot),
    .rf_bignum_wr_indirect_onehot_o  (rf_bignum_wr_indirect_onehot),
    .rf_bignum_indirect_en_o         (rf_bignum_indirect_en),

    // To/from base ALU
    .alu_base_operation_o        (alu_base_operation),
    .alu_base_comparison_o       (alu_base_comparison),
    .alu_base_operation_result_i (alu_base_operation_result),
    .alu_base_comparison_result_i(alu_base_comparison_result),

    // To/from bignum ALU
    .alu_bignum_operation_o       (alu_bignum_operation),
    .alu_bignum_operation_valid_o (alu_bignum_operation_valid),
    .alu_bignum_operation_commit_o(alu_bignum_operation_commit),
    .alu_bignum_operation_result_i(alu_bignum_operation_result),
    .alu_bignum_selection_flag_i  (alu_bignum_selection_flag),

    // To/from bignum MAC
    .mac_bignum_operation_o       (mac_bignum_operation),
    .mac_bignum_operation_result_i(mac_bignum_operation_result),
    .mac_bignum_en_o              (mac_bignum_en),
    .mac_bignum_commit_o          (mac_bignum_commit),

    // To/from LSU (base and bignum)
    .lsu_load_req_o          (lsu_load_req),
    .lsu_store_req_o         (lsu_store_req),
    .lsu_req_subset_o        (lsu_req_subset),
    .lsu_addr_o              (lsu_addr),
    .lsu_addr_en_predec_i    (lsu_addr_en_predec),

    .lsu_base_wdata_o  (lsu_base_wdata),
    .lsu_bignum_wdata_o(lsu_bignum_wdata),

    .lsu_base_rdata_i  (lsu_base_rdata),
    .lsu_bignum_rdata_i(lsu_bignum_rdata),

    // Isprs read/write (base and bignum)
    .ispr_addr_o             (ispr_addr),
    .ispr_base_wdata_o       (ispr_base_wdata),
    .ispr_base_wr_en_o       (ispr_base_wr_en),
    .ispr_bignum_wdata_intg_o(ispr_bignum_wdata_intg),
    .ispr_bignum_wr_en_o     (ispr_bignum_wr_en),
    .ispr_flags_wr_o         (ispr_flags_wr),
    .ispr_wr_commit_o        (ispr_wr_commit),
    .ispr_rdata_intg_i       (ispr_rdata_intg),
    .ispr_rd_en_o            (ispr_rd_en),

    // RND interface
    .rnd_req_o         (rnd_req),
    .rnd_prefetch_req_o(rnd_prefetch_req),
    .rnd_valid_i       (rnd_valid),

    .urnd_reseed_err_i(urnd_reseed_err),

    // Secure wipe
    .secure_wipe_req_o     (secure_wipe_req),
    .secure_wipe_ack_i     (secure_wipe_ack),
    .sec_wipe_zero_i       (sec_wipe_zero),
    .secure_wipe_running_i (secure_wipe_running_o),

    .state_reset_i(state_reset),
    .insn_cnt_o   (insn_cnt),
    .insn_cnt_clear_i,
    .mems_sec_wipe_o,

    .software_errs_fatal_i,

    .sideload_key_shares_valid_i,

    .prefetch_en_o             (prefetch_en),
    .prefetch_loop_active_o    (prefetch_loop_active),
    .prefetch_loop_iterations_o(prefetch_loop_iterations),
    .prefetch_loop_end_addr_o  (prefetch_loop_end_addr),
    .prefetch_loop_jump_addr_o (prefetch_loop_jump_addr),
    .prefetch_ignore_errs_o    (prefetch_ignore_errs),

    .ctrl_flow_predec_i       (ctrl_flow_predec),
    .ctrl_flow_target_predec_i(ctrl_flow_target_predec),
    .predec_error_o           (controller_predec_error)
  );

  `ASSERT(InsnDataStableInStall, u_otbn_controller.state_q == OtbnStateStall |->
                                 insn_fetch_resp_data == $past(insn_fetch_resp_data))

  // Spot the fatal error bits from the controller
  logic controller_fatal_err;
  assign controller_fatal_err = |{controller_err_bits.fatal_software,
                                  controller_err_bits.bad_internal_state,
                                  controller_err_bits.reg_intg_violation};

  logic non_controller_reg_intg_violation;
  assign non_controller_reg_intg_violation =
      |{alu_bignum_reg_intg_violation_err, mac_bignum_reg_intg_violation_err, rf_base_intg_err};


  // Generate an err_bits output by combining errors from all the blocks in otbn_core
  assign err_bits_d = '{
    fatal_software:      controller_err_bits.fatal_software,
    bad_internal_state:  |{controller_err_bits.bad_internal_state,
                           start_stop_fatal_error,
                           urnd_all_zero,
                           predec_error,
                           insn_addr_err,
                           rf_base_spurious_we_err,
                           mubi_err},
    reg_intg_violation:  |{controller_err_bits.reg_intg_violation,
                           non_controller_reg_intg_violation},
    dmem_intg_violation: lsu_rdata_err,
    imem_intg_violation: insn_fetch_err,
    rnd_fips_chk_fail:   rnd_fips_err,
    rnd_rep_chk_fail:    rnd_rep_err,
    key_invalid:         controller_err_bits.key_invalid,
    loop:                controller_err_bits.loop,
    illegal_insn:        controller_err_bits.illegal_insn,
    call_stack:          controller_err_bits.call_stack,
    bad_insn_addr:       controller_err_bits.bad_insn_addr,
    bad_data_addr:       controller_err_bits.bad_data_addr
  };

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_bits_q <= '0;
    end else begin
      if (start_i && !locking_o) begin
        err_bits_q <= '0;
      end else begin
        err_bits_q <= err_bits_q | err_bits_d;
      end
    end
  end
  assign err_bits_o = err_bits_q | err_bits_d;

  // Pass an "escalation" signal down to the controller by ORing in error signals from the other
  // modules in otbn_core. Note that each error signal except escalate_en_i that appears here also
  // appears somewhere in err_bits_o above (checked in ErrBitsIfControllerEscalate_A)
  assign controller_fatal_escalate_en =
      mubi4_or_hi(escalate_en_i,
                  mubi4_bool_to_mubi(|{start_stop_fatal_error, urnd_all_zero, predec_error,
                                       rf_base_intg_err, rf_base_spurious_we_err, lsu_rdata_err,
                                       insn_fetch_err, non_controller_reg_intg_violation,
                                       insn_addr_err}));

  assign controller_recov_escalate_en =
      mubi4_bool_to_mubi(|{rnd_rep_err, rnd_fips_err});

  // Similarly for the start/stop controller
  assign start_stop_escalate_en =
      mubi4_or_hi(escalate_en_i,
                  mubi4_bool_to_mubi(|{urnd_all_zero, rf_base_intg_err, rf_base_spurious_we_err,
                                       predec_error, lsu_rdata_err, insn_fetch_err,
                                       controller_fatal_err, insn_addr_err}));

  // Signal error if MuBi input signals take on invalid values as this means something bad is
  // happening. The explicit error detection is required as the mubi4_or_hi operations above
  // might mask invalid values depending on other input operands.
  assign mubi_err = mubi4_test_invalid(escalate_en_i);

  assign insn_cnt_o = insn_cnt;

  // Load store unit: read and write data from data memory
  otbn_lsu u_otbn_lsu (
    .clk_i,
    .rst_ni,

    // Data memory interface
    .dmem_req_o,
    .dmem_write_o,
    .dmem_addr_o,
    .dmem_wdata_o,
    .dmem_wmask_o,
    .dmem_rmask_o,
    .dmem_rdata_i,
    .dmem_rvalid_i,
    .dmem_rerror_i,

    .lsu_load_req_i  (lsu_load_req),
    .lsu_store_req_i (lsu_store_req),
    .lsu_req_subset_i(lsu_req_subset),
    .lsu_addr_i      (lsu_addr),

    .lsu_base_wdata_i  (lsu_base_wdata),
    .lsu_bignum_wdata_i(lsu_bignum_wdata),

    .lsu_base_rdata_o  (lsu_base_rdata),
    .lsu_bignum_rdata_o(lsu_bignum_rdata),
    .lsu_rdata_err_o   (lsu_rdata_err)
  );

  // Base Instruction Subset =======================================================================

  otbn_rf_base #(
    .RegFile(RegFile)
  ) u_otbn_rf_base (
    .clk_i,
    .rst_ni,

    .state_reset_i         (state_reset),
    .sec_wipe_stack_reset_i(sec_wipe_zero),

    .wr_addr_i         (rf_base_wr_addr),
    .wr_en_i           (rf_base_wr_en),
    .wr_data_no_intg_i (rf_base_wr_data_no_intg),
    .wr_data_intg_i    (rf_base_wr_data_intg),
    .wr_data_intg_sel_i(rf_base_wr_data_intg_sel),
    .wr_commit_i       (rf_base_wr_commit),

    .rd_addr_a_i     (rf_base_rd_addr_a),
    .rd_en_a_i       (rf_base_rd_en_a),
    .rd_data_a_intg_o(rf_base_rd_data_a_intg),
    .rd_addr_b_i     (rf_base_rd_addr_b),
    .rd_en_b_i       (rf_base_rd_en_b),
    .rd_data_b_intg_o(rf_base_rd_data_b_intg),
    .rd_commit_i     (rf_base_rd_commit),

    .call_stack_sw_err_o(rf_base_call_stack_sw_err),
    .call_stack_hw_err_o(rf_base_call_stack_hw_err),
    .intg_err_o         (rf_base_intg_err),
    .spurious_we_err_o  (rf_base_spurious_we_err)
  );

  assign rf_base_wr_addr         = sec_wipe_base ? sec_wipe_addr : rf_base_wr_addr_ctrl;
  assign rf_base_wr_en           = sec_wipe_base ? 1'b1          : rf_base_wr_en_ctrl;
  assign rf_base_wr_commit       = sec_wipe_base ? 1'b1          : rf_base_wr_commit_ctrl;

  // Write data to Base RF
  always_comb begin
    if (sec_wipe_base) begin
      // Wipe the Base RF with either random numbers or zeroes.
      if (sec_wipe_base_urnd) begin
        rf_base_wr_data_no_intg = urnd_data[31:0];
      end else begin
        rf_base_wr_data_no_intg = 32'b0;
      end
      rf_base_wr_data_intg_sel = 0;
    end else begin
      rf_base_wr_data_no_intg = rf_base_wr_data_no_intg_ctrl;
      rf_base_wr_data_intg_sel = rf_base_wr_data_intg_sel_ctrl;
    end
  end

  otbn_alu_base u_otbn_alu_base (
    .clk_i,
    .rst_ni,

    .operation_i        (alu_base_operation),
    .comparison_i       (alu_base_comparison),
    .operation_result_o (alu_base_operation_result),
    .comparison_result_o(alu_base_comparison_result)
  );

  otbn_rf_bignum #(
    .RegFile(RegFile)
  ) u_otbn_rf_bignum (
    .clk_i,
    .rst_ni,

    .wr_addr_i         (rf_bignum_wr_addr),
    .wr_en_i           (rf_bignum_wr_en),
    .wr_commit_i       (rf_bignum_wr_commit),
    .wr_data_no_intg_i (rf_bignum_wr_data_no_intg),
    .wr_data_intg_i    (rf_bignum_wr_data_intg),
    .wr_data_intg_sel_i(rf_bignum_wr_data_intg_sel),

    .rd_addr_a_i     (rf_bignum_rd_addr_a),
    .rd_en_a_i       (rf_bignum_rd_en_a),
    .rd_data_a_intg_o(rf_bignum_rd_data_a_intg),
    .rd_addr_b_i     (rf_bignum_rd_addr_b),
    .rd_en_b_i       (rf_bignum_rd_en_b),
    .rd_data_b_intg_o(rf_bignum_rd_data_b_intg),

    .intg_err_o(rf_bignum_intg_err),

    .rf_predec_bignum_i(rf_predec_bignum),
    .predec_error_o    (rf_bignum_predec_error),

    .spurious_we_err_o(rf_bignum_spurious_we_err)
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if(!rst_ni) begin
      sec_wipe_wdr_q <= 1'b0;
    end else begin
      sec_wipe_wdr_q <= sec_wipe_wdr_d;
    end
  end

  always_ff @(posedge clk_i) begin
    if (sec_wipe_wdr_d) begin
      sec_wipe_wdr_addr_q <= sec_wipe_addr;
      sec_wipe_wdr_urnd_q <= sec_wipe_wdr_urnd_d;
    end
  end

  assign rf_bignum_wr_addr   = sec_wipe_wdr_q ? sec_wipe_wdr_addr_q : rf_bignum_wr_addr_ctrl;
  assign rf_bignum_wr_en     = sec_wipe_wdr_q ? 2'b11               : rf_bignum_wr_en_ctrl;
  assign rf_bignum_wr_commit = sec_wipe_wdr_q ? 1'b1                : rf_bignum_wr_commit_ctrl;

  // Write data to WDR
  always_comb begin
    if (sec_wipe_wdr_q) begin
      // Wipe the WDR with either random numbers or zeroes.
      if (sec_wipe_wdr_urnd_q) begin
        rf_bignum_wr_data_no_intg = urnd_data;
      end else begin
        rf_bignum_wr_data_no_intg = 256'b0;
      end
      rf_bignum_wr_data_intg_sel = 0;
    end else begin
      rf_bignum_wr_data_no_intg = rf_bignum_wr_data_no_intg_ctrl;
      rf_bignum_wr_data_intg_sel = rf_bignum_wr_data_intg_sel_ctrl;
    end
  end

  otbn_alu_bignum u_otbn_alu_bignum (
    .clk_i,
    .rst_ni,

    .operation_i       (alu_bignum_operation),
    .operation_valid_i (alu_bignum_operation_valid),
    .operation_commit_i(alu_bignum_operation_commit),
    .operation_result_o(alu_bignum_operation_result),
    .selection_flag_o  (alu_bignum_selection_flag),

    .alu_predec_bignum_i (alu_predec_bignum),
    .ispr_predec_bignum_i(ispr_predec_bignum),

    .ispr_addr_i             (ispr_addr),
    .ispr_base_wdata_i       (ispr_base_wdata),
    .ispr_base_wr_en_i       (ispr_base_wr_en),
    .ispr_bignum_wdata_intg_i(ispr_bignum_wdata_intg),
    .ispr_bignum_wr_en_i     (ispr_bignum_wr_en),
    .ispr_flags_wr_i         (ispr_flags_wr),
    .ispr_wr_commit_i        (ispr_wr_commit),
    .ispr_init_i             (ispr_init),
    .ispr_rdata_intg_o       (ispr_rdata_intg),
    .ispr_rd_en_i            (ispr_rd_en),

    .ispr_acc_intg_i        (ispr_acc_intg),
    .ispr_acc_wr_data_intg_o(ispr_acc_wr_data_intg),
    .ispr_acc_wr_en_o       (ispr_acc_wr_en),

    .reg_intg_violation_err_o(alu_bignum_reg_intg_violation_err),

    .sec_wipe_mod_urnd_i(sec_wipe_mod_urnd),

    .mac_operation_flags_i   (mac_bignum_operation_flags),
    .mac_operation_flags_en_i(mac_bignum_operation_flags_en),

    .rnd_data_i (rnd_data),
    .urnd_data_i(urnd_data),

    .sideload_key_shares_i,

    .alu_predec_error_o(alu_bignum_predec_error),
    .ispr_predec_error_o(ispr_predec_error)
  );

  otbn_mac_bignum u_otbn_mac_bignum (
    .clk_i,
    .rst_ni,

    .operation_i                    (mac_bignum_operation),
    .operation_result_o             (mac_bignum_operation_result),
    .operation_flags_o              (mac_bignum_operation_flags),
    .operation_flags_en_o           (mac_bignum_operation_flags_en),
    .operation_intg_violation_err_o (mac_bignum_reg_intg_violation_err),

    .mac_predec_bignum_i(mac_predec_bignum),
    .predec_error_o     (mac_bignum_predec_error),

    .urnd_data_i        (urnd_data),
    .sec_wipe_acc_urnd_i(sec_wipe_acc_urnd),

    .mac_en_i    (mac_bignum_en),
    .mac_commit_i(mac_bignum_commit),

    .ispr_acc_intg_o        (ispr_acc_intg),
    .ispr_acc_wr_data_intg_i(ispr_acc_wr_data_intg),
    .ispr_acc_wr_en_i       (ispr_acc_wr_en)
  );

  otbn_rnd #(
    .RndCnstUrndPrngSeed(RndCnstUrndPrngSeed)
  ) u_otbn_rnd (
    .clk_i,
    .rst_ni,

    .opn_start_i (controller_start),
    .opn_end_i   (secure_wipe_req),

    .rnd_req_i         (rnd_req),
    .rnd_prefetch_req_i(rnd_prefetch_req),
    .rnd_valid_o       (rnd_valid),
    .rnd_data_o        (rnd_data),
    .rnd_rep_err_o     (rnd_rep_err),
    .rnd_fips_err_o    (rnd_fips_err),

    .urnd_reseed_req_i (urnd_reseed_req),
    .urnd_reseed_ack_o (urnd_reseed_ack),
    .urnd_advance_i    (urnd_advance),
    .urnd_data_o       (urnd_data),
    .urnd_all_zero_o   (urnd_all_zero),

    .edn_rnd_req_o,
    .edn_rnd_ack_i,
    .edn_rnd_data_i,
    .edn_rnd_fips_i,
    .edn_rnd_err_i,

    .edn_urnd_req_o,
    .edn_urnd_ack_i,
    .edn_urnd_data_i
  );

  // Advance URND either when the start_stop_control commands it or when temporary secure wipe keys
  // are requested.
  // When SecMuteUrnd is enabled, signal urnd_advance_start_stop_control is muted. Therefore, it is
  // necessary to enable urnd_advance using ispr_predec_bignum.ispr_rd_en[IsprUrnd] whenever URND
  // data are consumed by the ALU.
  assign urnd_advance = urnd_advance_start_stop_control | req_sec_wipe_urnd_keys_q |
                        (SecMuteUrnd & ispr_predec_bignum.ispr_rd_en[IsprUrnd]);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      req_sec_wipe_urnd_keys_q <= 1'b0;
    end else begin
      req_sec_wipe_urnd_keys_q <= req_sec_wipe_urnd_keys_i;
    end
  end

  assign dmem_sec_wipe_urnd_key_o = urnd_data[127:0];
  assign imem_sec_wipe_urnd_key_o = urnd_data[255:128];

  // Asserts =======================================================================================

  // All outputs should be known.
  `ASSERT_KNOWN(DoneOKnown_A, done_o)
  `ASSERT_KNOWN(ImemReqOKnown_A, imem_req_o)
  `ASSERT_KNOWN_IF(ImemAddrOKnown_A, imem_addr_o, imem_req_o)
  `ASSERT_KNOWN(DmemReqOKnown_A, dmem_req_o)
  `ASSERT_KNOWN_IF(DmemWriteOKnown_A, dmem_write_o, dmem_req_o)
  `ASSERT_KNOWN_IF(DmemAddrOKnown_A, dmem_addr_o, dmem_req_o)
  `ASSERT_KNOWN_IF(DmemWdataOKnown_A, dmem_wdata_o, dmem_req_o & dmem_write_o)
  `ASSERT_KNOWN_IF(DmemWmaskOKnown_A, dmem_wmask_o, dmem_req_o & dmem_write_o)
  `ASSERT_KNOWN_IF(DmemRmaskOKnown_A, dmem_rmask_o, dmem_req_o)
  `ASSERT_KNOWN(EdnRndReqOKnown_A, edn_rnd_req_o)
  `ASSERT_KNOWN(EdnUrndReqOKnown_A, edn_urnd_req_o)
  `ASSERT_KNOWN(InsnCntOKnown_A, insn_cnt_o)
  `ASSERT_KNOWN(ErrBitsKnown_A, err_bits_o)

  // Keep the EDN requests active until they are acknowledged.
  `ASSERT(EdnRndReqStable_A, edn_rnd_req_o & ~edn_rnd_ack_i |=> edn_rnd_req_o)
  `ASSERT(EdnUrndReqStable_A, edn_urnd_req_o & ~edn_urnd_ack_i |=> edn_urnd_req_o)

  `ASSERT(OnlyWriteLoadDataBaseWhenDMemValid_A,
          rf_bignum_wr_en_ctrl & insn_dec_bignum.rf_wdata_sel == RfWdSelLsu |-> dmem_rvalid_i)
  `ASSERT(OnlyWriteLoadDataBignumWhenDMemValid_A,
          rf_base_wr_en_ctrl & insn_dec_base.rf_wdata_sel == RfWdSelLsu |-> dmem_rvalid_i)

  // Error handling: if we pass an error signal down to the controller then we should also be
  // setting an error flag, unless the signal came from above.
  `ASSERT(ErrBitsIfControllerEscalate_A,
          (mubi4_test_true_loose(controller_fatal_escalate_en) ||
           mubi4_test_true_loose(controller_recov_escalate_en)) &&
          mubi4_test_false_strict(escalate_en_i)
          |=> err_bits_q)

  // Similarly, if we pass an escalation signal down to the start/stop controller then we should
  // also be setting an error flag, unless the signal came from above.
  `ASSERT(ErrBitsIfStartStopEscalate_A,
          mubi4_test_true_loose(start_stop_escalate_en) && mubi4_test_false_strict(escalate_en_i)
          |=> err_bits_q)

  // The following assertions allow up to 400 cycles from escalation until the start/stop FSM locks.
  // This is a long time, but it's necessary because following an escalation the start/stop FSM goes
  // through two rounds of secure wiping with random data with an URND reseed in between.  Depending
  // on the delay configured in the EDN model, the reseed alone can take 200 cycles.

  `ASSERT(OtbnStartStopGlobalEscCntrMeasure_A, err_bits_q && mubi4_test_true_loose(escalate_en_i)
          && mubi4_test_true_loose(start_stop_escalate_en)|=> ##[1:400]
          u_otbn_start_stop_control.state_q == otbn_pkg::OtbnStartStopStateLocked)

  `ASSERT(OtbnStartStopLocalEscCntrMeasure_A, err_bits_q && mubi4_test_false_strict(escalate_en_i)
          && mubi4_test_true_loose(start_stop_escalate_en) |=>  ##[1:400]
          u_otbn_start_stop_control.state_q == otbn_pkg::OtbnStartStopStateLocked)

  // In contrast to the start/stop FSM, the controller FSM should lock quickly after an escalation,
  // independent of the secure wipe.

  `ASSERT(OtbnControllerGlobalEscCntrMeasure_A, err_bits_q && mubi4_test_true_loose(escalate_en_i)
          && mubi4_test_true_loose(controller_fatal_escalate_en)|=> ##[1:100]
          u_otbn_controller.state_q == otbn_pkg::OtbnStateLocked)

  `ASSERT(OtbnControllerLocalEscCntrMeasure_A, err_bits_q && mubi4_test_false_strict(escalate_en_i)
          && mubi4_test_true_loose(controller_fatal_escalate_en) |=>  ##[1:100]
          u_otbn_controller.state_q == otbn_pkg::OtbnStateLocked)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package otbn_reg_pkg;

  // Param list
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 16;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    logic        q;
  } otbn_reg2hw_intr_state_reg_t;

  typedef struct packed {
    logic        q;
  } otbn_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    logic        q;
    logic        qe;
  } otbn_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } fatal;
    struct packed {
      logic        q;
      logic        qe;
    } recov;
  } otbn_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic [7:0]  q;
    logic        qe;
  } otbn_reg2hw_cmd_reg_t;

  typedef struct packed {
    logic        q;
    logic        qe;
  } otbn_reg2hw_ctrl_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } bad_data_addr;
    struct packed {
      logic        q;
      logic        qe;
    } bad_insn_addr;
    struct packed {
      logic        q;
      logic        qe;
    } call_stack;
    struct packed {
      logic        q;
      logic        qe;
    } illegal_insn;
    struct packed {
      logic        q;
      logic        qe;
    } loop;
    struct packed {
      logic        q;
      logic        qe;
    } key_invalid;
    struct packed {
      logic        q;
      logic        qe;
    } rnd_rep_chk_fail;
    struct packed {
      logic        q;
      logic        qe;
    } rnd_fips_chk_fail;
    struct packed {
      logic        q;
      logic        qe;
    } imem_intg_violation;
    struct packed {
      logic        q;
      logic        qe;
    } dmem_intg_violation;
    struct packed {
      logic        q;
      logic        qe;
    } reg_intg_violation;
    struct packed {
      logic        q;
      logic        qe;
    } bus_intg_violation;
    struct packed {
      logic        q;
      logic        qe;
    } bad_internal_state;
    struct packed {
      logic        q;
      logic        qe;
    } illegal_bus_access;
    struct packed {
      logic        q;
      logic        qe;
    } lifecycle_escalation;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_software;
  } otbn_reg2hw_err_bits_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } otbn_reg2hw_insn_cnt_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } otbn_reg2hw_load_checksum_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } otbn_hw2reg_intr_state_reg_t;

  typedef struct packed {
    logic        d;
  } otbn_hw2reg_ctrl_reg_t;

  typedef struct packed {
    logic [7:0]  d;
    logic        de;
  } otbn_hw2reg_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } bad_data_addr;
    struct packed {
      logic        d;
    } bad_insn_addr;
    struct packed {
      logic        d;
    } call_stack;
    struct packed {
      logic        d;
    } illegal_insn;
    struct packed {
      logic        d;
    } loop;
    struct packed {
      logic        d;
    } key_invalid;
    struct packed {
      logic        d;
    } rnd_rep_chk_fail;
    struct packed {
      logic        d;
    } rnd_fips_chk_fail;
    struct packed {
      logic        d;
    } imem_intg_violation;
    struct packed {
      logic        d;
    } dmem_intg_violation;
    struct packed {
      logic        d;
    } reg_intg_violation;
    struct packed {
      logic        d;
    } bus_intg_violation;
    struct packed {
      logic        d;
    } bad_internal_state;
    struct packed {
      logic        d;
    } illegal_bus_access;
    struct packed {
      logic        d;
    } lifecycle_escalation;
    struct packed {
      logic        d;
    } fatal_software;
  } otbn_hw2reg_err_bits_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } imem_intg_violation;
    struct packed {
      logic        d;
      logic        de;
    } dmem_intg_violation;
    struct packed {
      logic        d;
      logic        de;
    } reg_intg_violation;
    struct packed {
      logic        d;
      logic        de;
    } bus_intg_violation;
    struct packed {
      logic        d;
      logic        de;
    } bad_internal_state;
    struct packed {
      logic        d;
      logic        de;
    } illegal_bus_access;
    struct packed {
      logic        d;
      logic        de;
    } lifecycle_escalation;
    struct packed {
      logic        d;
      logic        de;
    } fatal_software;
  } otbn_hw2reg_fatal_alert_cause_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } otbn_hw2reg_insn_cnt_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } otbn_hw2reg_load_checksum_reg_t;

  // Register -> HW type
  typedef struct packed {
    otbn_reg2hw_intr_state_reg_t intr_state; // [116:116]
    otbn_reg2hw_intr_enable_reg_t intr_enable; // [115:115]
    otbn_reg2hw_intr_test_reg_t intr_test; // [114:113]
    otbn_reg2hw_alert_test_reg_t alert_test; // [112:109]
    otbn_reg2hw_cmd_reg_t cmd; // [108:100]
    otbn_reg2hw_ctrl_reg_t ctrl; // [99:98]
    otbn_reg2hw_err_bits_reg_t err_bits; // [97:66]
    otbn_reg2hw_insn_cnt_reg_t insn_cnt; // [65:33]
    otbn_reg2hw_load_checksum_reg_t load_checksum; // [32:0]
  } otbn_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    otbn_hw2reg_intr_state_reg_t intr_state; // [107:106]
    otbn_hw2reg_ctrl_reg_t ctrl; // [105:105]
    otbn_hw2reg_status_reg_t status; // [104:96]
    otbn_hw2reg_err_bits_reg_t err_bits; // [95:80]
    otbn_hw2reg_fatal_alert_cause_reg_t fatal_alert_cause; // [79:64]
    otbn_hw2reg_insn_cnt_reg_t insn_cnt; // [63:32]
    otbn_hw2reg_load_checksum_reg_t load_checksum; // [31:0]
  } otbn_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] OTBN_INTR_STATE_OFFSET = 16'h 0;
  parameter logic [BlockAw-1:0] OTBN_INTR_ENABLE_OFFSET = 16'h 4;
  parameter logic [BlockAw-1:0] OTBN_INTR_TEST_OFFSET = 16'h 8;
  parameter logic [BlockAw-1:0] OTBN_ALERT_TEST_OFFSET = 16'h c;
  parameter logic [BlockAw-1:0] OTBN_CMD_OFFSET = 16'h 10;
  parameter logic [BlockAw-1:0] OTBN_CTRL_OFFSET = 16'h 14;
  parameter logic [BlockAw-1:0] OTBN_STATUS_OFFSET = 16'h 18;
  parameter logic [BlockAw-1:0] OTBN_ERR_BITS_OFFSET = 16'h 1c;
  parameter logic [BlockAw-1:0] OTBN_FATAL_ALERT_CAUSE_OFFSET = 16'h 20;
  parameter logic [BlockAw-1:0] OTBN_INSN_CNT_OFFSET = 16'h 24;
  parameter logic [BlockAw-1:0] OTBN_LOAD_CHECKSUM_OFFSET = 16'h 28;

  // Reset values for hwext registers and their fields
  parameter logic [0:0] OTBN_INTR_TEST_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_INTR_TEST_DONE_RESVAL = 1'h 0;
  parameter logic [1:0] OTBN_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] OTBN_ALERT_TEST_FATAL_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ALERT_TEST_RECOV_RESVAL = 1'h 0;
  parameter logic [7:0] OTBN_CMD_RESVAL = 8'h 0;
  parameter logic [7:0] OTBN_CMD_CMD_RESVAL = 8'h 0;
  parameter logic [0:0] OTBN_CTRL_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_CTRL_SOFTWARE_ERRS_FATAL_RESVAL = 1'h 0;
  parameter logic [23:0] OTBN_ERR_BITS_RESVAL = 24'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_BAD_DATA_ADDR_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_BAD_INSN_ADDR_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_CALL_STACK_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_ILLEGAL_INSN_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_LOOP_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_KEY_INVALID_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_RND_REP_CHK_FAIL_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_RND_FIPS_CHK_FAIL_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_IMEM_INTG_VIOLATION_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_DMEM_INTG_VIOLATION_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_REG_INTG_VIOLATION_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_BUS_INTG_VIOLATION_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_BAD_INTERNAL_STATE_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_ILLEGAL_BUS_ACCESS_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_LIFECYCLE_ESCALATION_RESVAL = 1'h 0;
  parameter logic [0:0] OTBN_ERR_BITS_FATAL_SOFTWARE_RESVAL = 1'h 0;
  parameter logic [31:0] OTBN_INSN_CNT_RESVAL = 32'h 0;
  parameter logic [31:0] OTBN_INSN_CNT_INSN_CNT_RESVAL = 32'h 0;
  parameter logic [31:0] OTBN_LOAD_CHECKSUM_RESVAL = 32'h 0;
  parameter logic [31:0] OTBN_LOAD_CHECKSUM_CHECKSUM_RESVAL = 32'h 0;

  // Window parameters
  parameter logic [BlockAw-1:0] OTBN_IMEM_OFFSET = 16'h 4000;
  parameter int unsigned        OTBN_IMEM_SIZE   = 'h 1000;
  parameter logic [BlockAw-1:0] OTBN_DMEM_OFFSET = 16'h 8000;
  parameter int unsigned        OTBN_DMEM_SIZE   = 'h c00;

  // Register index
  typedef enum int {
    OTBN_INTR_STATE,
    OTBN_INTR_ENABLE,
    OTBN_INTR_TEST,
    OTBN_ALERT_TEST,
    OTBN_CMD,
    OTBN_CTRL,
    OTBN_STATUS,
    OTBN_ERR_BITS,
    OTBN_FATAL_ALERT_CAUSE,
    OTBN_INSN_CNT,
    OTBN_LOAD_CHECKSUM
  } otbn_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] OTBN_PERMIT [11] = '{
    4'b 0001, // index[ 0] OTBN_INTR_STATE
    4'b 0001, // index[ 1] OTBN_INTR_ENABLE
    4'b 0001, // index[ 2] OTBN_INTR_TEST
    4'b 0001, // index[ 3] OTBN_ALERT_TEST
    4'b 0001, // index[ 4] OTBN_CMD
    4'b 0001, // index[ 5] OTBN_CTRL
    4'b 0001, // index[ 6] OTBN_STATUS
    4'b 0111, // index[ 7] OTBN_ERR_BITS
    4'b 0001, // index[ 8] OTBN_FATAL_ALERT_CAUSE
    4'b 1111, // index[ 9] OTBN_INSN_CNT
    4'b 1111  // index[10] OTBN_LOAD_CHECKSUM
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module otbn_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // Output port for window
  output tlul_pkg::tl_h2d_t tl_win_o  [2],
  input  tlul_pkg::tl_d2h_t tl_win_i  [2],

  // To HW
  output otbn_reg_pkg::otbn_reg2hw_t reg2hw, // Write
  input  otbn_reg_pkg::otbn_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import otbn_reg_pkg::* ;

  localparam int AW = 16;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [10:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(11)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(0)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  tlul_pkg::tl_h2d_t tl_socket_h2d [3];
  tlul_pkg::tl_d2h_t tl_socket_d2h [3];

  logic [1:0] reg_steer;

  // socket_1n connection
  assign tl_reg_h2d = tl_socket_h2d[2];
  assign tl_socket_d2h[2] = tl_reg_d2h;

  assign tl_win_o[0] = tl_socket_h2d[0];
  assign tl_socket_d2h[0] = tl_win_i[0];
  assign tl_win_o[1] = tl_socket_h2d[1];
  assign tl_socket_d2h[1] = tl_win_i[1];

  // Create Socket_1n
  tlul_socket_1n #(
    .N            (3),
    .HReqPass     (1'b1),
    .HRspPass     (1'b1),
    .DReqPass     ({3{1'b1}}),
    .DRspPass     ({3{1'b1}}),
    .HReqDepth    (4'h0),
    .HRspDepth    (4'h0),
    .DReqDepth    ({3{4'h0}}),
    .DRspDepth    ({3{4'h0}}),
    .ExplicitErrs (1'b0)
  ) u_socket (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),
    .tl_h_i (tl_i),
    .tl_h_o (tl_o_pre),
    .tl_d_o (tl_socket_h2d),
    .tl_d_i (tl_socket_d2h),
    .dev_select_i (reg_steer)
  );

  // Create steering logic
  always_comb begin
    reg_steer =
        tl_i.a_address[AW-1:0] inside {[16384:20479]} ? 2'd0 :
        tl_i.a_address[AW-1:0] inside {[32768:35839]} ? 2'd1 :
        // Default set to register
        2'd2;

    // Override this in case of an integrity error
    if (intg_err) begin
      reg_steer = 2'd2;
    end
  end

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(1)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_qs;
  logic intr_state_wd;
  logic intr_enable_we;
  logic intr_enable_qs;
  logic intr_enable_wd;
  logic intr_test_we;
  logic intr_test_wd;
  logic alert_test_we;
  logic alert_test_fatal_wd;
  logic alert_test_recov_wd;
  logic cmd_we;
  logic [7:0] cmd_wd;
  logic ctrl_re;
  logic ctrl_we;
  logic ctrl_qs;
  logic ctrl_wd;
  logic [7:0] status_qs;
  logic err_bits_re;
  logic err_bits_we;
  logic err_bits_bad_data_addr_qs;
  logic err_bits_bad_data_addr_wd;
  logic err_bits_bad_insn_addr_qs;
  logic err_bits_bad_insn_addr_wd;
  logic err_bits_call_stack_qs;
  logic err_bits_call_stack_wd;
  logic err_bits_illegal_insn_qs;
  logic err_bits_illegal_insn_wd;
  logic err_bits_loop_qs;
  logic err_bits_loop_wd;
  logic err_bits_key_invalid_qs;
  logic err_bits_key_invalid_wd;
  logic err_bits_rnd_rep_chk_fail_qs;
  logic err_bits_rnd_rep_chk_fail_wd;
  logic err_bits_rnd_fips_chk_fail_qs;
  logic err_bits_rnd_fips_chk_fail_wd;
  logic err_bits_imem_intg_violation_qs;
  logic err_bits_imem_intg_violation_wd;
  logic err_bits_dmem_intg_violation_qs;
  logic err_bits_dmem_intg_violation_wd;
  logic err_bits_reg_intg_violation_qs;
  logic err_bits_reg_intg_violation_wd;
  logic err_bits_bus_intg_violation_qs;
  logic err_bits_bus_intg_violation_wd;
  logic err_bits_bad_internal_state_qs;
  logic err_bits_bad_internal_state_wd;
  logic err_bits_illegal_bus_access_qs;
  logic err_bits_illegal_bus_access_wd;
  logic err_bits_lifecycle_escalation_qs;
  logic err_bits_lifecycle_escalation_wd;
  logic err_bits_fatal_software_qs;
  logic err_bits_fatal_software_wd;
  logic fatal_alert_cause_imem_intg_violation_qs;
  logic fatal_alert_cause_dmem_intg_violation_qs;
  logic fatal_alert_cause_reg_intg_violation_qs;
  logic fatal_alert_cause_bus_intg_violation_qs;
  logic fatal_alert_cause_bad_internal_state_qs;
  logic fatal_alert_cause_illegal_bus_access_qs;
  logic fatal_alert_cause_lifecycle_escalation_qs;
  logic fatal_alert_cause_fatal_software_qs;
  logic insn_cnt_re;
  logic insn_cnt_we;
  logic [31:0] insn_cnt_qs;
  logic [31:0] insn_cnt_wd;
  logic load_checksum_re;
  logic load_checksum_we;
  logic [31:0] load_checksum_qs;
  logic [31:0] load_checksum_wd;

  // Register instances
  // R[intr_state]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.de),
    .d      (hw2reg.intr_state.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_qs)
  );


  // R[intr_enable]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [0:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[fatal]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.fatal.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal.qe = alert_test_qe;

  //   F[recov]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.recov.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov.qe = alert_test_qe;


  // R[cmd]: V(True)
  logic cmd_qe;
  logic [0:0] cmd_flds_we;
  assign cmd_qe = &cmd_flds_we;
  prim_subreg_ext #(
    .DW    (8)
  ) u_cmd (
    .re     (1'b0),
    .we     (cmd_we),
    .wd     (cmd_wd),
    .d      ('0),
    .qre    (),
    .qe     (cmd_flds_we[0]),
    .q      (reg2hw.cmd.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.cmd.qe = cmd_qe;


  // R[ctrl]: V(True)
  logic ctrl_qe;
  logic [0:0] ctrl_flds_we;
  assign ctrl_qe = &ctrl_flds_we;
  prim_subreg_ext #(
    .DW    (1)
  ) u_ctrl (
    .re     (ctrl_re),
    .we     (ctrl_we),
    .wd     (ctrl_wd),
    .d      (hw2reg.ctrl.d),
    .qre    (),
    .qe     (ctrl_flds_we[0]),
    .q      (reg2hw.ctrl.q),
    .ds     (),
    .qs     (ctrl_qs)
  );
  assign reg2hw.ctrl.qe = ctrl_qe;


  // R[status]: V(False)
  prim_subreg #(
    .DW      (8),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (8'h4)
  ) u_status (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.status.de),
    .d      (hw2reg.status.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (status_qs)
  );


  // R[err_bits]: V(True)
  logic err_bits_qe;
  logic [15:0] err_bits_flds_we;
  assign err_bits_qe = &err_bits_flds_we;
  //   F[bad_data_addr]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_bad_data_addr (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_bad_data_addr_wd),
    .d      (hw2reg.err_bits.bad_data_addr.d),
    .qre    (),
    .qe     (err_bits_flds_we[0]),
    .q      (reg2hw.err_bits.bad_data_addr.q),
    .ds     (),
    .qs     (err_bits_bad_data_addr_qs)
  );
  assign reg2hw.err_bits.bad_data_addr.qe = err_bits_qe;

  //   F[bad_insn_addr]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_bad_insn_addr (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_bad_insn_addr_wd),
    .d      (hw2reg.err_bits.bad_insn_addr.d),
    .qre    (),
    .qe     (err_bits_flds_we[1]),
    .q      (reg2hw.err_bits.bad_insn_addr.q),
    .ds     (),
    .qs     (err_bits_bad_insn_addr_qs)
  );
  assign reg2hw.err_bits.bad_insn_addr.qe = err_bits_qe;

  //   F[call_stack]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_call_stack (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_call_stack_wd),
    .d      (hw2reg.err_bits.call_stack.d),
    .qre    (),
    .qe     (err_bits_flds_we[2]),
    .q      (reg2hw.err_bits.call_stack.q),
    .ds     (),
    .qs     (err_bits_call_stack_qs)
  );
  assign reg2hw.err_bits.call_stack.qe = err_bits_qe;

  //   F[illegal_insn]: 3:3
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_illegal_insn (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_illegal_insn_wd),
    .d      (hw2reg.err_bits.illegal_insn.d),
    .qre    (),
    .qe     (err_bits_flds_we[3]),
    .q      (reg2hw.err_bits.illegal_insn.q),
    .ds     (),
    .qs     (err_bits_illegal_insn_qs)
  );
  assign reg2hw.err_bits.illegal_insn.qe = err_bits_qe;

  //   F[loop]: 4:4
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_loop (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_loop_wd),
    .d      (hw2reg.err_bits.loop.d),
    .qre    (),
    .qe     (err_bits_flds_we[4]),
    .q      (reg2hw.err_bits.loop.q),
    .ds     (),
    .qs     (err_bits_loop_qs)
  );
  assign reg2hw.err_bits.loop.qe = err_bits_qe;

  //   F[key_invalid]: 5:5
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_key_invalid (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_key_invalid_wd),
    .d      (hw2reg.err_bits.key_invalid.d),
    .qre    (),
    .qe     (err_bits_flds_we[5]),
    .q      (reg2hw.err_bits.key_invalid.q),
    .ds     (),
    .qs     (err_bits_key_invalid_qs)
  );
  assign reg2hw.err_bits.key_invalid.qe = err_bits_qe;

  //   F[rnd_rep_chk_fail]: 6:6
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_rnd_rep_chk_fail (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_rnd_rep_chk_fail_wd),
    .d      (hw2reg.err_bits.rnd_rep_chk_fail.d),
    .qre    (),
    .qe     (err_bits_flds_we[6]),
    .q      (reg2hw.err_bits.rnd_rep_chk_fail.q),
    .ds     (),
    .qs     (err_bits_rnd_rep_chk_fail_qs)
  );
  assign reg2hw.err_bits.rnd_rep_chk_fail.qe = err_bits_qe;

  //   F[rnd_fips_chk_fail]: 7:7
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_rnd_fips_chk_fail (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_rnd_fips_chk_fail_wd),
    .d      (hw2reg.err_bits.rnd_fips_chk_fail.d),
    .qre    (),
    .qe     (err_bits_flds_we[7]),
    .q      (reg2hw.err_bits.rnd_fips_chk_fail.q),
    .ds     (),
    .qs     (err_bits_rnd_fips_chk_fail_qs)
  );
  assign reg2hw.err_bits.rnd_fips_chk_fail.qe = err_bits_qe;

  //   F[imem_intg_violation]: 16:16
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_imem_intg_violation (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_imem_intg_violation_wd),
    .d      (hw2reg.err_bits.imem_intg_violation.d),
    .qre    (),
    .qe     (err_bits_flds_we[8]),
    .q      (reg2hw.err_bits.imem_intg_violation.q),
    .ds     (),
    .qs     (err_bits_imem_intg_violation_qs)
  );
  assign reg2hw.err_bits.imem_intg_violation.qe = err_bits_qe;

  //   F[dmem_intg_violation]: 17:17
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_dmem_intg_violation (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_dmem_intg_violation_wd),
    .d      (hw2reg.err_bits.dmem_intg_violation.d),
    .qre    (),
    .qe     (err_bits_flds_we[9]),
    .q      (reg2hw.err_bits.dmem_intg_violation.q),
    .ds     (),
    .qs     (err_bits_dmem_intg_violation_qs)
  );
  assign reg2hw.err_bits.dmem_intg_violation.qe = err_bits_qe;

  //   F[reg_intg_violation]: 18:18
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_reg_intg_violation (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_reg_intg_violation_wd),
    .d      (hw2reg.err_bits.reg_intg_violation.d),
    .qre    (),
    .qe     (err_bits_flds_we[10]),
    .q      (reg2hw.err_bits.reg_intg_violation.q),
    .ds     (),
    .qs     (err_bits_reg_intg_violation_qs)
  );
  assign reg2hw.err_bits.reg_intg_violation.qe = err_bits_qe;

  //   F[bus_intg_violation]: 19:19
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_bus_intg_violation (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_bus_intg_violation_wd),
    .d      (hw2reg.err_bits.bus_intg_violation.d),
    .qre    (),
    .qe     (err_bits_flds_we[11]),
    .q      (reg2hw.err_bits.bus_intg_violation.q),
    .ds     (),
    .qs     (err_bits_bus_intg_violation_qs)
  );
  assign reg2hw.err_bits.bus_intg_violation.qe = err_bits_qe;

  //   F[bad_internal_state]: 20:20
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_bad_internal_state (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_bad_internal_state_wd),
    .d      (hw2reg.err_bits.bad_internal_state.d),
    .qre    (),
    .qe     (err_bits_flds_we[12]),
    .q      (reg2hw.err_bits.bad_internal_state.q),
    .ds     (),
    .qs     (err_bits_bad_internal_state_qs)
  );
  assign reg2hw.err_bits.bad_internal_state.qe = err_bits_qe;

  //   F[illegal_bus_access]: 21:21
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_illegal_bus_access (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_illegal_bus_access_wd),
    .d      (hw2reg.err_bits.illegal_bus_access.d),
    .qre    (),
    .qe     (err_bits_flds_we[13]),
    .q      (reg2hw.err_bits.illegal_bus_access.q),
    .ds     (),
    .qs     (err_bits_illegal_bus_access_qs)
  );
  assign reg2hw.err_bits.illegal_bus_access.qe = err_bits_qe;

  //   F[lifecycle_escalation]: 22:22
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_lifecycle_escalation (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_lifecycle_escalation_wd),
    .d      (hw2reg.err_bits.lifecycle_escalation.d),
    .qre    (),
    .qe     (err_bits_flds_we[14]),
    .q      (reg2hw.err_bits.lifecycle_escalation.q),
    .ds     (),
    .qs     (err_bits_lifecycle_escalation_qs)
  );
  assign reg2hw.err_bits.lifecycle_escalation.qe = err_bits_qe;

  //   F[fatal_software]: 23:23
  prim_subreg_ext #(
    .DW    (1)
  ) u_err_bits_fatal_software (
    .re     (err_bits_re),
    .we     (err_bits_we),
    .wd     (err_bits_fatal_software_wd),
    .d      (hw2reg.err_bits.fatal_software.d),
    .qre    (),
    .qe     (err_bits_flds_we[15]),
    .q      (reg2hw.err_bits.fatal_software.q),
    .ds     (),
    .qs     (err_bits_fatal_software_qs)
  );
  assign reg2hw.err_bits.fatal_software.qe = err_bits_qe;


  // R[fatal_alert_cause]: V(False)
  //   F[imem_intg_violation]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_imem_intg_violation (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.imem_intg_violation.de),
    .d      (hw2reg.fatal_alert_cause.imem_intg_violation.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_imem_intg_violation_qs)
  );

  //   F[dmem_intg_violation]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_dmem_intg_violation (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.dmem_intg_violation.de),
    .d      (hw2reg.fatal_alert_cause.dmem_intg_violation.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_dmem_intg_violation_qs)
  );

  //   F[reg_intg_violation]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_reg_intg_violation (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.reg_intg_violation.de),
    .d      (hw2reg.fatal_alert_cause.reg_intg_violation.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_reg_intg_violation_qs)
  );

  //   F[bus_intg_violation]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_bus_intg_violation (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.bus_intg_violation.de),
    .d      (hw2reg.fatal_alert_cause.bus_intg_violation.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_bus_intg_violation_qs)
  );

  //   F[bad_internal_state]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_bad_internal_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.bad_internal_state.de),
    .d      (hw2reg.fatal_alert_cause.bad_internal_state.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_bad_internal_state_qs)
  );

  //   F[illegal_bus_access]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_illegal_bus_access (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.illegal_bus_access.de),
    .d      (hw2reg.fatal_alert_cause.illegal_bus_access.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_illegal_bus_access_qs)
  );

  //   F[lifecycle_escalation]: 6:6
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_lifecycle_escalation (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.lifecycle_escalation.de),
    .d      (hw2reg.fatal_alert_cause.lifecycle_escalation.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_lifecycle_escalation_qs)
  );

  //   F[fatal_software]: 7:7
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_fatal_software (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.fatal_software.de),
    .d      (hw2reg.fatal_alert_cause.fatal_software.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_fatal_software_qs)
  );


  // R[insn_cnt]: V(True)
  logic insn_cnt_qe;
  logic [0:0] insn_cnt_flds_we;
  assign insn_cnt_qe = &insn_cnt_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_insn_cnt (
    .re     (insn_cnt_re),
    .we     (insn_cnt_we),
    .wd     (insn_cnt_wd),
    .d      (hw2reg.insn_cnt.d),
    .qre    (),
    .qe     (insn_cnt_flds_we[0]),
    .q      (reg2hw.insn_cnt.q),
    .ds     (),
    .qs     (insn_cnt_qs)
  );
  assign reg2hw.insn_cnt.qe = insn_cnt_qe;


  // R[load_checksum]: V(True)
  logic load_checksum_qe;
  logic [0:0] load_checksum_flds_we;
  assign load_checksum_qe = &load_checksum_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_load_checksum (
    .re     (load_checksum_re),
    .we     (load_checksum_we),
    .wd     (load_checksum_wd),
    .d      (hw2reg.load_checksum.d),
    .qre    (),
    .qe     (load_checksum_flds_we[0]),
    .q      (reg2hw.load_checksum.q),
    .ds     (),
    .qs     (load_checksum_qs)
  );
  assign reg2hw.load_checksum.qe = load_checksum_qe;



  logic [10:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == OTBN_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == OTBN_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == OTBN_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == OTBN_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == OTBN_CMD_OFFSET);
    addr_hit[ 5] = (reg_addr == OTBN_CTRL_OFFSET);
    addr_hit[ 6] = (reg_addr == OTBN_STATUS_OFFSET);
    addr_hit[ 7] = (reg_addr == OTBN_ERR_BITS_OFFSET);
    addr_hit[ 8] = (reg_addr == OTBN_FATAL_ALERT_CAUSE_OFFSET);
    addr_hit[ 9] = (reg_addr == OTBN_INSN_CNT_OFFSET);
    addr_hit[10] = (reg_addr == OTBN_LOAD_CHECKSUM_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(OTBN_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(OTBN_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(OTBN_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(OTBN_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(OTBN_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(OTBN_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(OTBN_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(OTBN_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(OTBN_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(OTBN_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(OTBN_PERMIT[10] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_wd = reg_wdata[0];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_wd = reg_wdata[0];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_wd = reg_wdata[0];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_fatal_wd = reg_wdata[0];

  assign alert_test_recov_wd = reg_wdata[1];
  assign cmd_we = addr_hit[4] & reg_we & !reg_error;

  assign cmd_wd = reg_wdata[7:0];
  assign ctrl_re = addr_hit[5] & reg_re & !reg_error;
  assign ctrl_we = addr_hit[5] & reg_we & !reg_error;

  assign ctrl_wd = reg_wdata[0];
  assign err_bits_re = addr_hit[7] & reg_re & !reg_error;
  assign err_bits_we = addr_hit[7] & reg_we & !reg_error;

  assign err_bits_bad_data_addr_wd = reg_wdata[0];

  assign err_bits_bad_insn_addr_wd = reg_wdata[1];

  assign err_bits_call_stack_wd = reg_wdata[2];

  assign err_bits_illegal_insn_wd = reg_wdata[3];

  assign err_bits_loop_wd = reg_wdata[4];

  assign err_bits_key_invalid_wd = reg_wdata[5];

  assign err_bits_rnd_rep_chk_fail_wd = reg_wdata[6];

  assign err_bits_rnd_fips_chk_fail_wd = reg_wdata[7];

  assign err_bits_imem_intg_violation_wd = reg_wdata[16];

  assign err_bits_dmem_intg_violation_wd = reg_wdata[17];

  assign err_bits_reg_intg_violation_wd = reg_wdata[18];

  assign err_bits_bus_intg_violation_wd = reg_wdata[19];

  assign err_bits_bad_internal_state_wd = reg_wdata[20];

  assign err_bits_illegal_bus_access_wd = reg_wdata[21];

  assign err_bits_lifecycle_escalation_wd = reg_wdata[22];

  assign err_bits_fatal_software_wd = reg_wdata[23];
  assign insn_cnt_re = addr_hit[9] & reg_re & !reg_error;
  assign insn_cnt_we = addr_hit[9] & reg_we & !reg_error;

  assign insn_cnt_wd = reg_wdata[31:0];
  assign load_checksum_re = addr_hit[10] & reg_re & !reg_error;
  assign load_checksum_we = addr_hit[10] & reg_we & !reg_error;

  assign load_checksum_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = cmd_we;
    reg_we_check[5] = ctrl_we;
    reg_we_check[6] = 1'b0;
    reg_we_check[7] = err_bits_we;
    reg_we_check[8] = 1'b0;
    reg_we_check[9] = insn_cnt_we;
    reg_we_check[10] = load_checksum_we;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[7:0] = '0;
      end

      addr_hit[5]: begin
        reg_rdata_next[0] = ctrl_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[7:0] = status_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[0] = err_bits_bad_data_addr_qs;
        reg_rdata_next[1] = err_bits_bad_insn_addr_qs;
        reg_rdata_next[2] = err_bits_call_stack_qs;
        reg_rdata_next[3] = err_bits_illegal_insn_qs;
        reg_rdata_next[4] = err_bits_loop_qs;
        reg_rdata_next[5] = err_bits_key_invalid_qs;
        reg_rdata_next[6] = err_bits_rnd_rep_chk_fail_qs;
        reg_rdata_next[7] = err_bits_rnd_fips_chk_fail_qs;
        reg_rdata_next[16] = err_bits_imem_intg_violation_qs;
        reg_rdata_next[17] = err_bits_dmem_intg_violation_qs;
        reg_rdata_next[18] = err_bits_reg_intg_violation_qs;
        reg_rdata_next[19] = err_bits_bus_intg_violation_qs;
        reg_rdata_next[20] = err_bits_bad_internal_state_qs;
        reg_rdata_next[21] = err_bits_illegal_bus_access_qs;
        reg_rdata_next[22] = err_bits_lifecycle_escalation_qs;
        reg_rdata_next[23] = err_bits_fatal_software_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[0] = fatal_alert_cause_imem_intg_violation_qs;
        reg_rdata_next[1] = fatal_alert_cause_dmem_intg_violation_qs;
        reg_rdata_next[2] = fatal_alert_cause_reg_intg_violation_qs;
        reg_rdata_next[3] = fatal_alert_cause_bus_intg_violation_qs;
        reg_rdata_next[4] = fatal_alert_cause_bad_internal_state_qs;
        reg_rdata_next[5] = fatal_alert_cause_illegal_bus_access_qs;
        reg_rdata_next[6] = fatal_alert_cause_lifecycle_escalation_qs;
        reg_rdata_next[7] = fatal_alert_cause_fatal_software_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = insn_cnt_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = load_checksum_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

/**
 * Scramble control for OTBN
 *
 * This provides a key and nonce for scrambling the OTBN IMem and DMem. The OTP
 * key interface is used to request a new key and nonce when they are requested.
 */
module otbn_scramble_ctrl
  import otbn_pkg::*;
#(
  // Default seed and nonce for scrambling
  parameter otp_ctrl_pkg::otbn_key_t   RndCnstOtbnKey   = otbn_pkg::RndCnstOtbnKeyDefault,
  parameter otp_ctrl_pkg::otbn_nonce_t RndCnstOtbnNonce = otbn_pkg::RndCnstOtbnNonceDefault
) (
  // OTBN clock
  input clk_i,
  input rst_ni,

  // OTP Clock (for key interface)
  input clk_otp_i,
  input rst_otp_ni,

  // OTP key interface
  output otp_ctrl_pkg::otbn_otp_key_req_t otbn_otp_key_o,
  input  otp_ctrl_pkg::otbn_otp_key_rsp_t otbn_otp_key_i,

  output otp_ctrl_pkg::otbn_key_t otbn_dmem_scramble_key_o,
  output otbn_dmem_nonce_t        otbn_dmem_scramble_nonce_o,
  output logic                    otbn_dmem_scramble_valid_o,
  output logic                    otbn_dmem_scramble_key_seed_valid_o,

  output otp_ctrl_pkg::otbn_key_t otbn_imem_scramble_key_o,
  output otbn_imem_nonce_t        otbn_imem_scramble_nonce_o,
  output logic                    otbn_imem_scramble_valid_o,
  output logic                    otbn_imem_scramble_key_seed_valid_o,

  input  logic                    otbn_dmem_scramble_sec_wipe_i,
  input  otp_ctrl_pkg::otbn_key_t otbn_dmem_scramble_sec_wipe_key_i,
  input  logic                    otbn_imem_scramble_sec_wipe_i,
  input  otp_ctrl_pkg::otbn_key_t otbn_imem_scramble_sec_wipe_key_i,

  output logic otbn_dmem_scramble_key_req_busy_o,
  output logic otbn_imem_scramble_key_req_busy_o,

  output logic state_error_o
);

  scramble_ctrl_state_e state_q, state_d;

  logic dmem_key_valid_q, dmem_key_valid_d;
  logic imem_key_valid_q, imem_key_valid_d;

  logic dmem_key_seed_valid_q, dmem_key_seed_valid_d;
  logic imem_key_seed_valid_q, imem_key_seed_valid_d;

  logic dmem_scramble_req_pending_q, dmem_scramble_req_pending_d;
  logic imem_scramble_req_pending_q, imem_scramble_req_pending_d;

  logic dmem_key_en, dmem_nonce_en;
  logic imem_key_en, imem_nonce_en;

  logic dmem_key_sel_otp;
  logic imem_key_sel_otp;

  otp_ctrl_pkg::otbn_key_t dmem_key_q, dmem_key_d;
  otp_ctrl_pkg::otbn_key_t imem_key_q, imem_key_d;

  otbn_dmem_nonce_t dmem_nonce_q;
  otbn_imem_nonce_t imem_nonce_q;

  logic                      otp_key_req, otp_key_ack;
  otp_ctrl_pkg::otbn_key_t   otp_key;
  otp_ctrl_pkg::otbn_nonce_t otp_nonce;
  logic                      otp_key_seed_valid;

  assign dmem_key_d = dmem_key_sel_otp ? otp_key : otbn_dmem_scramble_sec_wipe_key_i;
  assign imem_key_d = imem_key_sel_otp ? otp_key : otbn_imem_scramble_sec_wipe_key_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      dmem_key_q <= RndCnstOtbnKey;
    end else if (dmem_key_en) begin
      dmem_key_q <= dmem_key_d;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      dmem_nonce_q <= RndCnstOtbnNonce;
    end else if (dmem_nonce_en) begin
      dmem_nonce_q <= otp_nonce;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      imem_key_q <= RndCnstOtbnKey;
    end else if (imem_key_en) begin
      imem_key_q <= imem_key_d;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      imem_nonce_q <= RndCnstOtbnNonce;
    end else if (imem_nonce_en) begin
      imem_nonce_q <= otp_nonce;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      // Initial key and nonce are taken from defaults so on reset a valid key
      // is available.
      dmem_key_valid_q            <= 1'b1;
      imem_key_valid_q            <= 1'b1;
      dmem_key_seed_valid_q       <= 1'b0;
      imem_key_seed_valid_q       <= 1'b0;
      dmem_scramble_req_pending_q <= 1'b0;
      imem_scramble_req_pending_q <= 1'b0;
    end else begin
      dmem_key_valid_q            <= dmem_key_valid_d;
      imem_key_valid_q            <= imem_key_valid_d;
      dmem_key_seed_valid_q       <= dmem_key_seed_valid_d;
      imem_key_seed_valid_q       <= imem_key_seed_valid_d;
      dmem_scramble_req_pending_q <= dmem_scramble_req_pending_d;
      imem_scramble_req_pending_q <= imem_scramble_req_pending_d;
    end
  end

  // SEC_CM: SCRAMBLE_CTRL.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, scramble_ctrl_state_e, ScrambleCtrlIdle)

  always_comb begin
    dmem_key_valid_d            = dmem_key_valid_q;
    imem_key_valid_d            = imem_key_valid_q;
    dmem_key_seed_valid_d       = dmem_key_seed_valid_q;
    imem_key_seed_valid_d       = imem_key_seed_valid_q;
    dmem_key_en                 = 1'b0;
    dmem_nonce_en               = 1'b0;
    imem_key_en                 = 1'b0;
    imem_nonce_en               = 1'b0;
    dmem_scramble_req_pending_d = dmem_scramble_req_pending_q;
    imem_scramble_req_pending_d = imem_scramble_req_pending_q;
    dmem_key_sel_otp            = 1'b0;
    imem_key_sel_otp            = 1'b0;
    state_d                     = state_q;
    otp_key_req                 = 1'b0;
    state_error_o               = 1'b0;

    // Action dmem secure wipe request unless a new key request is already ongoing
    // SEC_CM: DATA.MEM.SEC_WIPE
    if (otbn_dmem_scramble_sec_wipe_i && state_q != ScrambleCtrlDmemReq) begin
      dmem_key_valid_d            = 1'b0;
      dmem_key_en                 = 1'b1;
      dmem_key_sel_otp            = 1'b0;
      dmem_scramble_req_pending_d = 1'b1;
    end

    // Action imem secure wipe request unless a new key request is already ongoing
    // SEC_CM: INSTRUCTION.MEM.SEC_WIPE
    if (otbn_imem_scramble_sec_wipe_i && state_q != ScrambleCtrlImemReq) begin
      imem_key_valid_d            = 1'b0;
      imem_key_en                 = 1'b1;
      imem_key_sel_otp            = 1'b0;
      imem_scramble_req_pending_d = 1'b1;
    end

    unique case (state_q)
      ScrambleCtrlIdle: begin
        if (dmem_scramble_req_pending_q) begin
          otp_key_req      = 1'b1;
          state_d          = ScrambleCtrlDmemReq;
        end else if (imem_scramble_req_pending_q) begin
          otp_key_req      = 1'b1;
          state_d          = ScrambleCtrlImemReq;
        end
      end
      ScrambleCtrlDmemReq: begin
        otp_key_req = 1'b1;

        if (otp_key_ack) begin
          state_d                     = ScrambleCtrlIdle;
          dmem_scramble_req_pending_d = 1'b0;
          dmem_key_en                 = 1'b1;
          dmem_nonce_en               = 1'b1;
          dmem_key_valid_d            = 1'b1;
          dmem_key_seed_valid_d       = otp_key_seed_valid;
          dmem_key_sel_otp            = 1'b1;
        end
      end ScrambleCtrlImemReq: begin
        otp_key_req = 1'b1;

        if (otp_key_ack) begin
          state_d                     = ScrambleCtrlIdle;
          imem_scramble_req_pending_d = 1'b0;
          imem_key_en                 = 1'b1;
          imem_nonce_en               = 1'b1;
          imem_key_valid_d            = 1'b1;
          imem_key_seed_valid_d       = otp_key_seed_valid;
          imem_key_sel_otp            = 1'b1;
        end
      end
      ScrambleCtrlError: begin
        // SEC_CM: SCRAMBLE_CTRL.FSM.LOCAL_ESC
        // Terminal error state
        state_error_o = 1'b1;
      end
      default: begin
        // We should never get here. If we do (e.g. via a malicious glitch), error out immediately.
        state_error_o = 1'b1;
        state_d = ScrambleCtrlError;
      end
    endcase
  end

  assign otbn_dmem_scramble_key_req_busy_o =
    (state_d == ScrambleCtrlDmemReq) | dmem_scramble_req_pending_d;

  assign otbn_imem_scramble_key_req_busy_o =
    (state_d == ScrambleCtrlImemReq) | imem_scramble_req_pending_d;

  prim_sync_reqack_data #(
    .Width($bits(otp_ctrl_pkg::otbn_otp_key_rsp_t)-1),
    .EnRstChks(1'b1),
    .DataSrc2Dst(1'b0)
  ) u_otp_key_req_sync (
    .clk_src_i (clk_i),
    .rst_src_ni(rst_ni),
    .clk_dst_i (clk_otp_i),
    .rst_dst_ni(rst_otp_ni),
    .req_chk_i (1'b1),
    .src_req_i (otp_key_req),
    .src_ack_o (otp_key_ack),
    .dst_req_o (otbn_otp_key_o.req),
    .dst_ack_i (otbn_otp_key_i.ack),
    .data_i    ({otbn_otp_key_i.key,
                 otbn_otp_key_i.nonce,
                 otbn_otp_key_i.seed_valid}),
    .data_o    ({otp_key,
                 otp_nonce,
                 otp_key_seed_valid})
  );

  assign otbn_dmem_scramble_key_o            = dmem_key_q;
  assign otbn_dmem_scramble_nonce_o          = dmem_nonce_q;
  assign otbn_dmem_scramble_valid_o          = dmem_key_valid_q;
  assign otbn_dmem_scramble_key_seed_valid_o = dmem_key_seed_valid_q;

  assign otbn_imem_scramble_key_o            = imem_key_q;
  assign otbn_imem_scramble_nonce_o          = imem_nonce_q;
  assign otbn_imem_scramble_valid_o          = imem_key_valid_q;
  assign otbn_imem_scramble_key_seed_valid_o = imem_key_seed_valid_q;

  `ASSERT(OtbnScrambleCtrlLocalEscCntrMeasure_A, state_error_o |=> state_q == ScrambleCtrlError)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

/**
 * OpenTitan Big Number Accelerator (OTBN)
 */
module otbn
  import prim_alert_pkg::*;
  import otbn_pkg::*;
  import otbn_reg_pkg::*;
#(
  parameter bit                   Stub         = 1'b0,
  parameter regfile_e             RegFile      = RegFileFF,
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},

  // Default seed for URND PRNG
  parameter urnd_prng_seed_t RndCnstUrndPrngSeed = RndCnstUrndPrngSeedDefault,

  // Disable URND advance when not in use. Useful for SCA only.
  parameter bit SecMuteUrnd = 1'b0,
  // Skip URND re-seed at the start of an operation. Useful for SCA only.
  parameter bit SecSkipUrndReseedAtStart = 1'b0,

  // Default seed and nonce for scrambling
  parameter otp_ctrl_pkg::otbn_key_t   RndCnstOtbnKey   = RndCnstOtbnKeyDefault,
  parameter otp_ctrl_pkg::otbn_nonce_t RndCnstOtbnNonce = RndCnstOtbnNonceDefault
) (
  input clk_i,
  input rst_ni,

  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // Inter-module signals
  output prim_mubi_pkg::mubi4_t idle_o,

  // Interrupts
  output logic intr_done_o,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // Lifecycle interfaces
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  input  lc_ctrl_pkg::lc_tx_t lc_rma_req_i,
  output lc_ctrl_pkg::lc_tx_t lc_rma_ack_o,

  // Memory configuration
  input prim_ram_1p_pkg::ram_1p_cfg_t ram_cfg_i,

  // EDN clock and interface
  input                     clk_edn_i,
  input                     rst_edn_ni,
  output edn_pkg::edn_req_t edn_rnd_o,
  input  edn_pkg::edn_rsp_t edn_rnd_i,

  output edn_pkg::edn_req_t edn_urnd_o,
  input  edn_pkg::edn_rsp_t edn_urnd_i,

  // Key request to OTP (running on clk_fixed)
  input                                   clk_otp_i,
  input                                   rst_otp_ni,
  output otp_ctrl_pkg::otbn_otp_key_req_t otbn_otp_key_o,
  input  otp_ctrl_pkg::otbn_otp_key_rsp_t otbn_otp_key_i,

  input keymgr_pkg::otbn_key_req_t keymgr_key_i
);

  import prim_mubi_pkg::*;
  import prim_util_pkg::vbits;

  logic rst_n;

  // hold module in reset permanently when stubbing
  if (Stub) begin : gen_stub_otbn
    assign rst_n = 1'b0;
  end else begin : gen_real_otbn
    assign rst_n = rst_ni;
  end

  // The OTBN_*_SIZE parameters are auto-generated by regtool and come from the bus window sizes;
  // they are given in bytes and must be powers of two.
  //
  // DMEM is actually a bit bigger than OTBN_DMEM_SIZE: there are an extra DmemScratchSizeByte bytes
  // that aren't accessible over the bus.
  localparam int ImemSizeByte = int'(otbn_reg_pkg::OTBN_IMEM_SIZE);
  localparam int DmemSizeByte = int'(otbn_reg_pkg::OTBN_DMEM_SIZE + DmemScratchSizeByte);

  localparam int ImemAddrWidth = vbits(ImemSizeByte);
  localparam int DmemAddrWidth = vbits(DmemSizeByte);

  `ASSERT_INIT(ImemSizePowerOfTwo, 2 ** ImemAddrWidth == ImemSizeByte)
  `ASSERT_INIT(DmemSizePowerOfTwo, 2 ** DmemAddrWidth == DmemSizeByte)

  logic start_d, start_q;
  logic busy_execute_d, busy_execute_q;
  logic done, done_core, locking, locking_q;
  logic busy_secure_wipe;
  logic init_sec_wipe_done_d, init_sec_wipe_done_q;
  logic illegal_bus_access_d, illegal_bus_access_q;
  logic missed_gnt_error_d, missed_gnt_error_q;
  logic dmem_sec_wipe;
  logic imem_sec_wipe;
  logic mems_sec_wipe;
  logic req_sec_wipe_urnd_keys;
  logic [127:0] dmem_sec_wipe_urnd_key, imem_sec_wipe_urnd_key;

  logic core_recoverable_err, recoverable_err_d, recoverable_err_q;
  mubi4_t core_escalate_en;

  core_err_bits_t     core_err_bits;
  non_core_err_bits_t non_core_err_bits, non_core_err_bits_d, non_core_err_bits_q;
  err_bits_t          err_bits, err_bits_d, err_bits_q;
  logic               err_bits_en;

  // ERR_BITS register should be cleared due to a write request from the host processor
  // when OTBN is not running.
  logic err_bits_clear;

  logic software_errs_fatal_q, software_errs_fatal_d;

  otbn_reg2hw_t reg2hw;
  otbn_hw2reg_t hw2reg;
  status_e      status_d, status_q;

  // Bus device windows, as specified in otbn.hjson
  typedef enum logic {
    TlWinImem = 1'b0,
    TlWinDmem = 1'b1
  } tl_win_e;

  tlul_pkg::tl_h2d_t tl_win_h2d[2];
  tlul_pkg::tl_d2h_t tl_win_d2h[2];

  // The clock can be gated and some registers can be updated as long as OTBN isn't currently
  // running. Other registers can only be updated when OTBN is in the Idle state (which also implies
  // we are not locked).
  logic is_not_running_d, is_not_running_q;
  logic otbn_dmem_scramble_key_req_busy, otbn_imem_scramble_key_req_busy;

  assign is_not_running_d = ~|{busy_execute_d,
                               otbn_dmem_scramble_key_req_busy,
                               otbn_imem_scramble_key_req_busy,
                               busy_secure_wipe};

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if(!rst_ni) begin
      // OTBN starts busy, performing the initial secure wipe.
      is_not_running_q  <= 1'b0;
    end else begin
      is_not_running_q  <= is_not_running_d;
    end
  end

  // Inter-module signals ======================================================

  // Note: This is not the same thing as STATUS == IDLE. For example, we want to allow clock gating
  // when locked.
  prim_mubi4_sender #(
    .ResetValue(prim_mubi_pkg::MuBi4True)
  ) u_prim_mubi4_sender (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi4_bool_to_mubi(is_not_running_q)),
    .mubi_o(idle_o)
  );

  // Lifecycle ==================================================================

  localparam int unsigned LcEscalateCopies = 2;
  lc_ctrl_pkg::lc_tx_t [LcEscalateCopies-1:0] lc_escalate_en;
  prim_lc_sync #(
    .NumCopies(LcEscalateCopies)
  ) u_lc_escalate_en_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i(lc_escalate_en_i),
    .lc_en_o(lc_escalate_en)
  );

  lc_ctrl_pkg::lc_tx_t lc_rma_req;
  prim_lc_sync #(
    .NumCopies(1)
  ) u_lc_rma_req_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i(lc_rma_req_i),
    .lc_en_o({lc_rma_req})
  );

  // Internally, OTBN uses MUBI types.
  mubi4_t mubi_rma_req, mubi_rma_ack;
  assign mubi_rma_req = lc_ctrl_pkg::lc_to_mubi4(lc_rma_req);

  // When stubbing, forward req to ack.
  if (Stub) begin : gen_stub_rma_ack
    assign lc_rma_ack_o = lc_rma_req;
  end else begin : gen_real_rma_ack
    assign lc_rma_ack_o = lc_ctrl_pkg::mubi4_to_lc(mubi_rma_ack);
  end

  // Interrupts ================================================================

  assign done = is_busy_status(status_q) & ~is_busy_status(status_d) & init_sec_wipe_done_q;

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_done (
    .clk_i,
    .rst_ni                (rst_n),
    .event_intr_i          (done),
    .reg2hw_intr_enable_q_i(reg2hw.intr_enable.q),
    .reg2hw_intr_test_q_i  (reg2hw.intr_test.q),
    .reg2hw_intr_test_qe_i (reg2hw.intr_test.qe),
    .reg2hw_intr_state_q_i (reg2hw.intr_state.q),
    .hw2reg_intr_state_de_o(hw2reg.intr_state.de),
    .hw2reg_intr_state_d_o (hw2reg.intr_state.d),
    .intr_o                (intr_done_o)
  );

  // Instruction Memory (IMEM) =================================================

  localparam int ImemSizeWords = ImemSizeByte / 4;
  localparam int ImemIndexWidth = vbits(ImemSizeWords);

  // Access select to IMEM: core (1), or bus (0)
  logic imem_access_core;

  logic imem_req;
  logic imem_gnt;
  logic imem_write;
  logic [ImemIndexWidth-1:0] imem_index;
  logic [38:0] imem_wdata;
  logic [38:0] imem_wmask;
  logic [38:0] imem_rdata;
  logic imem_rvalid;
  logic imem_illegal_bus_access;
  logic imem_missed_gnt;

  logic imem_req_core;
  logic imem_write_core;
  logic [ImemIndexWidth-1:0] imem_index_core;
  logic [38:0] imem_rdata_core;
  logic imem_rvalid_core;

  logic imem_req_bus;
  logic imem_dummy_response_q, imem_dummy_response_d;
  logic imem_write_bus;
  logic [ImemIndexWidth-1:0] imem_index_bus;
  logic [38:0] imem_wdata_bus;
  logic [38:0] imem_wmask_bus;
  logic [38:0] imem_rdata_bus, imem_rdata_bus_raw;
  logic imem_rdata_bus_en_q, imem_rdata_bus_en_d;
  logic [top_pkg::TL_DBW-1:0] imem_byte_mask_bus;
  logic imem_rvalid_bus;
  logic [1:0] imem_rerror_bus;

  logic imem_bus_intg_violation;

  typedef struct packed {
    logic        imem;
    logic [14:0] index;
    logic [31:0] wr_data;
  } mem_crc_data_in_t;

  logic             mem_crc_data_in_valid;
  mem_crc_data_in_t mem_crc_data_in;
  logic             set_crc;
  logic [31:0]      crc_in, crc_out;

  logic [ImemAddrWidth-1:0] imem_addr_core;
  assign imem_index_core = imem_addr_core[ImemAddrWidth-1:2];

  logic [1:0] unused_imem_addr_core_wordbits;
  assign unused_imem_addr_core_wordbits = imem_addr_core[1:0];

  otp_ctrl_pkg::otbn_key_t otbn_imem_scramble_key;
  otbn_imem_nonce_t        otbn_imem_scramble_nonce;
  logic                    otbn_imem_scramble_valid;
  logic                    unused_otbn_imem_scramble_key_seed_valid;

  otp_ctrl_pkg::otbn_key_t otbn_dmem_scramble_key;
  otbn_dmem_nonce_t        otbn_dmem_scramble_nonce;
  logic                    otbn_dmem_scramble_valid;
  logic                    unused_otbn_dmem_scramble_key_seed_valid;


  logic otbn_scramble_state_error;

  // SEC_CM: SCRAMBLE.KEY.SIDELOAD
  otbn_scramble_ctrl #(
    .RndCnstOtbnKey  (RndCnstOtbnKey),
    .RndCnstOtbnNonce(RndCnstOtbnNonce)
  ) u_otbn_scramble_ctrl (
    .clk_i,
    .rst_ni,

    .clk_otp_i,
    .rst_otp_ni,

    .otbn_otp_key_o,
    .otbn_otp_key_i,

    .otbn_dmem_scramble_key_o           (otbn_dmem_scramble_key),
    .otbn_dmem_scramble_nonce_o         (otbn_dmem_scramble_nonce),
    .otbn_dmem_scramble_valid_o         (otbn_dmem_scramble_valid),
    .otbn_dmem_scramble_key_seed_valid_o(unused_otbn_dmem_scramble_key_seed_valid),

    .otbn_imem_scramble_key_o           (otbn_imem_scramble_key),
    .otbn_imem_scramble_nonce_o         (otbn_imem_scramble_nonce),
    .otbn_imem_scramble_valid_o         (otbn_imem_scramble_valid),
    .otbn_imem_scramble_key_seed_valid_o(unused_otbn_imem_scramble_key_seed_valid),

    .otbn_dmem_scramble_sec_wipe_i    (dmem_sec_wipe),
    .otbn_dmem_scramble_sec_wipe_key_i(dmem_sec_wipe_urnd_key),
    .otbn_imem_scramble_sec_wipe_i    (imem_sec_wipe),
    .otbn_imem_scramble_sec_wipe_key_i(imem_sec_wipe_urnd_key),

    .otbn_dmem_scramble_key_req_busy_o(otbn_dmem_scramble_key_req_busy),
    .otbn_imem_scramble_key_req_busy_o(otbn_imem_scramble_key_req_busy),

    .state_error_o(otbn_scramble_state_error)
  );

  // SEC_CM: MEM.SCRAMBLE
  prim_ram_1p_scr #(
    .Width          (39),
    .Depth          (ImemSizeWords),
    .DataBitsPerMask(39),
    .EnableParity   (0),
    .DiffWidth      (39)
  ) u_imem (
    .clk_i,
    .rst_ni(rst_n),

    .key_valid_i(otbn_imem_scramble_valid),
    .key_i      (otbn_imem_scramble_key),
    .nonce_i    (otbn_imem_scramble_nonce),

    .req_i       (imem_req),
    .gnt_o       (imem_gnt),
    .write_i     (imem_write),
    .addr_i      (imem_index),
    .wdata_i     (imem_wdata),
    .wmask_i     (imem_wmask),
    .intg_error_i(locking),

    .rdata_o (imem_rdata),
    .rvalid_o(imem_rvalid),
    .raddr_o (),
    .rerror_o(),
    .cfg_i   (ram_cfg_i)
  );

  // We should never see a request that doesn't get granted. A fatal error is raised if this occurs.
  assign imem_missed_gnt = imem_req & ~imem_gnt;

  // IMEM access from main TL-UL bus
  logic imem_gnt_bus;
  // Always grant to bus accesses, when OTBN is running a dummy response is returned
  assign imem_gnt_bus = imem_req_bus;

  tlul_adapter_sram #(
    .SramAw          (ImemIndexWidth),
    .SramDw          (32),
    .Outstanding     (1),
    .ByteAccess      (0),
    .ErrOnRead       (0),
    .EnableDataIntgPt(1),
    .SecFifoPtr      (1)  // SEC_CM: TLUL_FIFO.CTR.REDUN
  ) u_tlul_adapter_sram_imem (
    .clk_i,
    .rst_ni      (rst_n),
    .tl_i        (tl_win_h2d[TlWinImem]),
    .tl_o        (tl_win_d2h[TlWinImem]),
    .en_ifetch_i (MuBi4False),
    .req_o       (imem_req_bus),
    .req_type_o  (),
    .gnt_i       (imem_gnt_bus),
    .we_o        (imem_write_bus),
    .addr_o      (imem_index_bus),
    .wdata_o     (imem_wdata_bus),
    .wmask_o     (imem_wmask_bus),
    .intg_error_o(imem_bus_intg_violation),
    .rdata_i     (imem_rdata_bus),
    .rvalid_i    (imem_rvalid_bus),
    .rerror_i    (imem_rerror_bus)
  );


  // Mux core and bus access into IMEM
  assign imem_access_core = busy_execute_q | start_q;

  assign imem_req   = imem_access_core ? imem_req_core        : imem_req_bus;
  assign imem_write = imem_access_core ? imem_write_core      : imem_write_bus;
  assign imem_index = imem_access_core ? imem_index_core      : imem_index_bus;
  assign imem_wdata = imem_access_core ? '0                   : imem_wdata_bus;

  assign imem_illegal_bus_access = imem_req_bus & imem_access_core;

  assign imem_dummy_response_d = imem_illegal_bus_access;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      imem_dummy_response_q <= 1'b0;
    end else begin
      imem_dummy_response_q <= imem_dummy_response_d;
    end
  end

  // The instruction memory only supports 32b word writes, so we hardcode its
  // wmask here.
  //
  // Since this could cause confusion if the bus tried to do a partial write
  // (which wasn't caught in the TLUL adapter for some reason), we assert that
  // the wmask signal from the bus is indeed '1 when it requests a write. We
  // don't have the corresponding check for writes from the core because the
  // core cannot perform writes (and has no imem_wmask_o port).
  assign imem_wmask = imem_access_core ? '1 : imem_wmask_bus;
  `ASSERT(ImemWmaskBusIsFullWord_A, imem_req_bus && imem_write_bus |-> imem_wmask_bus == '1)

  // SEC_CM: DATA_REG_SW.SCA
  // Blank bus read data interface during core operation to avoid leaking the currently executed
  // instruction from IMEM through the bus unintentionally. Also blank when OTBN is returning
  // a dummy response (responding to an illegal bus access) and when OTBN is locked.
  assign imem_rdata_bus_en_d = ~(busy_execute_d | start_d) & ~imem_dummy_response_d & ~locking;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
        imem_rdata_bus_en_q <= 1'b1;
    end else begin
        imem_rdata_bus_en_q <= imem_rdata_bus_en_d;
    end
  end

  prim_blanker #(.Width(39)) u_imem_rdata_bus_blanker (
    .in_i (imem_rdata),
    .en_i (imem_rdata_bus_en_q),
    .out_o(imem_rdata_bus_raw)
  );

  // When OTBN is locked all imem bus reads should return 0. The blanker produces the 0s, this adds
  // the appropriate ECC. When OTBN is not locked the output of the blanker is passed straight
  // through. Data bits are always left un-modified. A registered version of `locking` is used for
  // timing reasons. When a read comes in when `locking` has just been asserted, `locking_q` will be
  // set the following cycle and the rdata will be forced to 0 with appropriate ECC. When `locking`
  // is asserted the cycle the rdata is being returned no locking was ocurring when the request came
  // in so it is reasonable to proceed with returning the supplied integrity.
  assign imem_rdata_bus =
    {locking_q ? prim_secded_pkg::SecdedInv3932ZeroEcc : imem_rdata_bus_raw[38:32],
     imem_rdata_bus_raw[31:0]};

  `ASSERT(ImemRDataBusDisabledWhenCoreAccess_A, imem_access_core |-> !imem_rdata_bus_en_q)
  `ASSERT(ImemRDataBusEnabledWhenIdle_A, status_q == StatusIdle |-> imem_rdata_bus_en_q)
  `ASSERT(ImemRDataBusDisabledWhenLocked_A, locking |=> !imem_rdata_bus_en_q)
  `ASSERT(ImemRDataBusReadAsZeroWhenLocked_A,
    imem_rvalid_bus & locking |-> imem_rdata_bus_raw == '0)

  assign imem_rdata_core = imem_rdata;

  // When an illegal bus access is seen, always return a dummy response the follow cycle.
  assign imem_rvalid_bus = (~imem_access_core & imem_rvalid) | imem_dummy_response_q;
  assign imem_rvalid_core = imem_access_core ? imem_rvalid : 1'b0;

  assign imem_byte_mask_bus = tl_win_h2d[TlWinImem].a_mask;

  // No imem errors reported for bus reads. Integrity is carried through on the bus so integrity
  // checking on TL responses will pick up any errors.
  assign imem_rerror_bus = 2'b00;

  // Data Memory (DMEM) ========================================================

  localparam int DmemSizeWords = DmemSizeByte / (WLEN / 8);
  localparam int DmemIndexWidth = vbits(DmemSizeWords);

  localparam int DmemBusSizeWords = int'(otbn_reg_pkg::OTBN_DMEM_SIZE) / (WLEN / 8);
  localparam int DmemBusIndexWidth = vbits(DmemBusSizeWords);

  // Access select to DMEM: core (1), or bus (0)
  logic dmem_access_core;

  logic dmem_req;
  logic dmem_gnt;
  logic dmem_write;
  logic [DmemIndexWidth-1:0] dmem_index;
  logic [ExtWLEN-1:0] dmem_wdata;
  logic [ExtWLEN-1:0] dmem_wmask;
  logic [ExtWLEN-1:0] dmem_rdata;
  logic dmem_rvalid;
  logic [BaseWordsPerWLEN*2-1:0] dmem_rerror_vec;
  logic dmem_rerror;
  logic dmem_illegal_bus_access;
  logic dmem_missed_gnt;

  logic dmem_req_core;
  logic dmem_write_core;
  logic [DmemIndexWidth-1:0] dmem_index_core;
  logic [ExtWLEN-1:0] dmem_wdata_core;
  logic [ExtWLEN-1:0] dmem_wmask_core;
  logic [BaseWordsPerWLEN-1:0] dmem_rmask_core_q, dmem_rmask_core_d;
  logic [ExtWLEN-1:0] dmem_rdata_core;
  logic dmem_rvalid_core;
  logic dmem_rerror_core;

  logic dmem_req_bus;
  logic dmem_dummy_response_q, dmem_dummy_response_d;
  logic dmem_write_bus;
  logic [DmemBusIndexWidth-1:0] dmem_index_bus;
  logic [ExtWLEN-1:0] dmem_wdata_bus;
  logic [ExtWLEN-1:0] dmem_wmask_bus;
  logic [ExtWLEN-1:0] dmem_rdata_bus, dmem_rdata_bus_raw;
  logic dmem_rdata_bus_en_q, dmem_rdata_bus_en_d;
  logic [DmemAddrWidth-1:0] dmem_addr_bus;
  logic unused_dmem_addr_bus;
  logic [31:0] dmem_wdata_narrow_bus;
  logic [top_pkg::TL_DBW-1:0] dmem_byte_mask_bus;
  logic dmem_rvalid_bus;
  logic [1:0] dmem_rerror_bus;

  logic dmem_bus_intg_violation;

  logic [DmemAddrWidth-1:0] dmem_addr_core;
  assign dmem_index_core = dmem_addr_core[DmemAddrWidth-1:DmemAddrWidth-DmemIndexWidth];

  logic unused_dmem_addr_core_wordbits;
  assign unused_dmem_addr_core_wordbits = ^dmem_addr_core[DmemAddrWidth-DmemIndexWidth-1:0];

  logic mubi_err;

  // SEC_CM: MEM.SCRAMBLE
  prim_ram_1p_scr #(
    .Width             (ExtWLEN),
    .Depth             (DmemSizeWords),
    .DataBitsPerMask   (39),
    .EnableParity      (0),
    .DiffWidth         (39),
    .ReplicateKeyStream(1)
  ) u_dmem (
    .clk_i,
    .rst_ni(rst_n),

    .key_valid_i(otbn_dmem_scramble_valid),
    .key_i      (otbn_dmem_scramble_key),
    .nonce_i    (otbn_dmem_scramble_nonce),

    .req_i       (dmem_req),
    .gnt_o       (dmem_gnt),
    .write_i     (dmem_write),
    .addr_i      (dmem_index),
    .wdata_i     (dmem_wdata),
    .wmask_i     (dmem_wmask),
    .intg_error_i(locking),

    .rdata_o (dmem_rdata),
    .rvalid_o(dmem_rvalid),
    .raddr_o (),
    .rerror_o(),
    .cfg_i   (ram_cfg_i)
  );

  // We should never see a request that doesn't get granted. A fatal error is raised if this occurs.
  assign dmem_missed_gnt = dmem_req & !dmem_gnt;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      dmem_rmask_core_q <= '0;
    end else begin
      if (dmem_req_core) begin
        dmem_rmask_core_q <= dmem_rmask_core_d;
      end
    end
  end

  // SEC_CM: DATA.MEM.INTEGRITY
  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; ++i_word) begin : g_dmem_intg_check
    logic [1:0] dmem_rerror_raw;

    // Separate check for dmem read data integrity outside of `u_dmem` as `prim_ram_1p_adv` doesn't
    // have functionality for only integrity checking, just fully integrated ECC. Integrity bits are
    // implemented on a 32-bit granule so separate checks are required for each.
    prim_secded_inv_39_32_dec u_dmem_intg_check (
      .data_i    (dmem_rdata[i_word*39+:39]),
      .data_o    (),
      .syndrome_o(),
      .err_o     (dmem_rerror_raw)
    );

    // Only report an error where the word was actually accessed. Otherwise uninitialised memory
    // that OTBN isn't using will cause false errors. dmem_rerror is only reported for reads from
    // OTBN. For Ibex reads integrity checking on TL responses will serve the same purpose.
    assign dmem_rerror_vec[i_word*2 +: 2] = dmem_rerror_raw &
        {2{dmem_rmask_core_q[i_word] & dmem_rvalid & dmem_access_core}};
  end

  // dmem_rerror_vec is 2 bits wide and is used to report ECC errors. Bit 1 is set if there's an
  // uncorrectable error and bit 0 is set if there's a correctable error. However, we're treating
  // all errors as fatal, so OR the two signals together.
  //zdr: dmem ecc disable
  assign dmem_rerror = (|dmem_rerror_vec)  & 1'b0;
  // assign dmem_rerror = |dmem_rerror_vec;

  // DMEM access from main TL-UL bus
  logic dmem_gnt_bus;
  // Always grant to bus accesses, when OTBN is running a dummy response is returned
  assign dmem_gnt_bus = dmem_req_bus;

  tlul_adapter_sram #(
    .SramAw          (DmemBusIndexWidth),
    .SramDw          (WLEN),
    .Outstanding     (1),
    .ByteAccess      (0),
    .ErrOnRead       (0),
    .EnableDataIntgPt(1),
    .SecFifoPtr      (1)  // SEC_CM: TLUL_FIFO.CTR.REDUN
  ) u_tlul_adapter_sram_dmem (
    .clk_i,
    .rst_ni      (rst_n),
    .tl_i        (tl_win_h2d[TlWinDmem]),
    .tl_o        (tl_win_d2h[TlWinDmem]),
    .en_ifetch_i (MuBi4False),
    .req_o       (dmem_req_bus),
    .req_type_o  (),
    .gnt_i       (dmem_gnt_bus),
    .we_o        (dmem_write_bus),
    .addr_o      (dmem_index_bus),
    .wdata_o     (dmem_wdata_bus),
    .wmask_o     (dmem_wmask_bus),
    .intg_error_o(dmem_bus_intg_violation),
    .rdata_i     (dmem_rdata_bus),
    .rvalid_i    (dmem_rvalid_bus),
    .rerror_i    (dmem_rerror_bus)
  );

  // Mux core and bus access into dmem
  assign dmem_access_core = busy_execute_q;

  assign dmem_req = dmem_access_core ? dmem_req_core : dmem_req_bus;
  assign dmem_write = dmem_access_core ? dmem_write_core : dmem_write_bus;
  assign dmem_wmask = dmem_access_core ? dmem_wmask_core : dmem_wmask_bus;
  // SEC_CM: DATA.MEM.SW_NOACCESS
  assign dmem_index = dmem_access_core ? dmem_index_core : dmem_index_bus;
  assign dmem_wdata = dmem_access_core ? dmem_wdata_core : dmem_wdata_bus;

  assign dmem_illegal_bus_access = dmem_req_bus & dmem_access_core;

  assign dmem_dummy_response_d = dmem_illegal_bus_access;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      dmem_dummy_response_q <= 1'b0;
    end else begin
      dmem_dummy_response_q <= dmem_dummy_response_d;
    end
  end

  // SEC_CM: DATA_REG_SW.SCA
  // Blank bus read data interface during core operation to avoid leaking DMEM data through the bus
  // unintentionally. Also blank when OTBN is returning a dummy response (responding to an illegal
  // bus access) and when OTBN is locked.
  assign dmem_rdata_bus_en_d = ~(busy_execute_d | start_d) & ~dmem_dummy_response_d & ~locking;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
        dmem_rdata_bus_en_q <= 1'b1;
    end else begin
        dmem_rdata_bus_en_q <= dmem_rdata_bus_en_d;
    end
  end

  prim_blanker #(.Width(ExtWLEN)) u_dmem_rdata_bus_blanker (
    .in_i (dmem_rdata),
    .en_i (dmem_rdata_bus_en_q),
    .out_o(dmem_rdata_bus_raw)
  );

  // When OTBN is locked all dmem bus reads should return 0. The blanker produces the 0s, this adds
  // the appropriate ECC. When OTBN is not locked the output of the blanker is passed straight
  // through. Data bits are always left un-modified. A registered version of `locking` is used for
  // timing reasons. When a read comes in when `locking` has just been asserted, `locking_q` will be
  // timing reasons. When a read comes in when `locking` has just been asserted, `locking_q` will be
  // set the following cycle and the rdata will be forced to 0 with appropriate ECC. When `locking`
  // is asserted the cycle the rdata is being returned no locking was ocurring when the request came
  // in so it is reasonable to proceed with returning the supplied integrity.
  for (genvar i_word = 0; i_word < BaseWordsPerWLEN; ++i_word) begin : g_dmem_rdata_bus
    assign dmem_rdata_bus[i_word*39+:39] =
      {locking_q ? prim_secded_pkg::SecdedInv3932ZeroEcc : dmem_rdata_bus_raw[i_word*39+32+:7],
       dmem_rdata_bus_raw[i_word*39+:32]};
  end

  `ASSERT(DmemRDataBusDisabledWhenCoreAccess_A, dmem_access_core |-> !dmem_rdata_bus_en_q)
  `ASSERT(DmemRDataBusEnabledWhenIdle_A, status_q == StatusIdle |-> dmem_rdata_bus_en_q)
  `ASSERT(DmemRDataBusDisabledWhenLocked_A, locking |=> !dmem_rdata_bus_en_q)
  `ASSERT(DmemRDataBusReadAsZeroWhenLocked_A,
    dmem_rvalid_bus & locking |-> dmem_rdata_bus_raw == '0)

  assign dmem_rdata_core = dmem_rdata;

  // When an illegal bus access is seen, always return a dummy response the follow cycle.
  assign dmem_rvalid_bus  = (~dmem_access_core & dmem_rvalid) | dmem_dummy_response_q;
  assign dmem_rvalid_core = dmem_access_core ? dmem_rvalid : 1'b0;

  // No dmem errors reported for bus reads. Integrity is carried through on the bus so integrity
  // checking on TL responses will pick up any errors.
  assign dmem_rerror_bus  = 2'b00;
  assign dmem_rerror_core = dmem_rerror;

  assign dmem_addr_bus = tl_win_h2d[TlWinDmem].a_address[DmemAddrWidth-1:0];
  assign dmem_wdata_narrow_bus = tl_win_h2d[TlWinDmem].a_data[31:0];
  assign dmem_byte_mask_bus = tl_win_h2d[TlWinDmem].a_mask;

  // Memory Load Integrity =====================================================
  // CRC logic below assumes a incoming data bus width of 32 bits
  `ASSERT_INIT(TLDWIs32Bit_A, top_pkg::TL_DW == 32)

  // Only advance CRC calculation on full 32-bit writes;
  assign mem_crc_data_in_valid   = ~(dmem_access_core | imem_access_core) &
      ((imem_req_bus & (imem_byte_mask_bus == 4'hf)) |
       (dmem_req_bus & (dmem_byte_mask_bus == 4'hf)));

  assign mem_crc_data_in.wr_data = imem_req_bus ? imem_wdata_bus[31:0] :
                                                  dmem_wdata_narrow_bus[31:0];
  assign mem_crc_data_in.index   = imem_req_bus ? {{15 - ImemIndexWidth{1'b0}}, imem_index_bus} :
                                                   {{15 - (DmemAddrWidth - 2){1'b0}},
                                                    dmem_addr_bus[DmemAddrWidth-1:2]};
  assign mem_crc_data_in.imem    = imem_req_bus;

  // Only the bits that factor into the dmem index and dmem word enables are required
  assign unused_dmem_addr_bus = ^{dmem_addr_bus[DmemAddrWidth-1:DmemIndexWidth],
                                  dmem_addr_bus[1:0]};

  // SEC_CM: WRITE.MEM.INTEGRITY
  prim_crc32 #(
    .BytesPerWord(6)
  ) u_mem_load_crc32 (
    .clk_i (clk_i),
    .rst_ni(rst_ni),

    .set_crc_i(set_crc),
    .crc_in_i (crc_in),

    .data_valid_i(mem_crc_data_in_valid),
    .data_i      (mem_crc_data_in),
    .crc_out_o   (crc_out)
  );

  assign set_crc = reg2hw.load_checksum.qe;
  assign crc_in = reg2hw.load_checksum.q;
  assign hw2reg.load_checksum.d = crc_out;

  // Registers =================================================================

  logic reg_bus_intg_violation;

  otbn_reg_top u_reg (
    .clk_i,
    .rst_ni  (rst_n),
    .tl_i,
    .tl_o,
    .tl_win_o(tl_win_h2d),
    .tl_win_i(tl_win_d2h),

    .reg2hw,
    .hw2reg,

    .intg_err_o(reg_bus_intg_violation),
    .devmode_i (1'b1)
  );

  // SEC_CM: BUS.INTEGRITY
  // SEC_CM: TLUL_FIFO.CTR.REDUN
  logic bus_intg_violation;
  assign bus_intg_violation = (imem_bus_intg_violation | dmem_bus_intg_violation |
                               reg_bus_intg_violation);

  // CMD register
  always_comb begin
    // start is flopped to avoid long timing paths from the TL fabric into OTBN internals.
    start_d       = 1'b0;
    dmem_sec_wipe = 1'b0;
    imem_sec_wipe = 1'b0;

    // Can only start a new command when idle.
    if (status_q == StatusIdle) begin
      if (reg2hw.cmd.qe) begin
        unique case (reg2hw.cmd.q)
          CmdExecute:     start_d       = 1'b1;
          CmdSecWipeDmem: dmem_sec_wipe = 1'b1;
          CmdSecWipeImem: imem_sec_wipe = 1'b1;
          default: ;
        endcase
      end
    end else if (busy_execute_q) begin
      // OTBN can command a secure wipe of IMEM and DMEM. This occurs when OTBN encounters a fatal
      // error.
      if (mems_sec_wipe) begin
        dmem_sec_wipe = 1'b1;
        imem_sec_wipe = 1'b1;
      end
    end
  end

  assign req_sec_wipe_urnd_keys = dmem_sec_wipe | imem_sec_wipe;

  assign illegal_bus_access_d = dmem_illegal_bus_access | imem_illegal_bus_access;

  // It should not be possible to request an imem or dmem access without it being granted. Either
  // a scramble key is present so the request will be granted or the core is busy obtaining a new
  // key, so no request can occur (the core won't generate one whilst awaiting a scrambling key and
  // the bus requests get an immediate dummy response bypassing the dmem or imem). A fatal error is
  // raised if request is seen without a grant.
  assign missed_gnt_error_d = dmem_missed_gnt | imem_missed_gnt;

  // Flop `illegal_bus_access_q` and `missed_gnt_error_q` to break timing paths from the TL
  // interface into the OTBN core.
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      start_q              <= 1'b0;
      illegal_bus_access_q <= 1'b0;
      missed_gnt_error_q   <= 1'b0;
    end else begin
      start_q              <= start_d;
      illegal_bus_access_q <= illegal_bus_access_d;
      missed_gnt_error_q   <= missed_gnt_error_d;
    end
  end

  // STATUS register
  // imem/dmem scramble req can be busy when locked, so use a priority selection so locked status
  // always takes priority.
  //
  // Note that these signals are all "a cycle early". For example, the locking signal gets asserted
  // combinatorially on the cycle that an error is injected. The STATUS register change, done
  // interrupt and any change to the idle signal will be delayed by 2 cycles.
  assign status_d = locking                         ? StatusLocked          :
                    busy_secure_wipe                ? StatusBusySecWipeInt  :
                    busy_execute_d                  ? StatusBusyExecute     :
                    otbn_dmem_scramble_key_req_busy ? StatusBusySecWipeDmem :
                    otbn_imem_scramble_key_req_busy ? StatusBusySecWipeImem :
                                                      StatusIdle;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      status_q <= StatusBusySecWipeInt;
    end else begin
      status_q <= status_d;
    end
  end

  assign hw2reg.status.d = status_q;
  assign hw2reg.status.de = 1'b1;

  // Only certain combinations of the state variable {locking, busy_execute_d,
  // otbn_dmem_scramble_key_req_busy, otbn_imem_scramble_key_req_busy} are possible.
  //
  // (1) When we finish (with a pulse on "done_core", which might stay high in the "locking"
  //     signal), busy_execute_d is guaranteed to be low. (Assertion: NotBusyAndDone_A)
  //
  // (2) There aren't really any other restrictions when locking is low: if there is an error during
  //     an operation, we'll start rotating memory keys while doing the internal secure wipe, so
  //     may see all of the signals high except locking.
  //
  // (3) Once locking is high, we guarantee never to see a new execution or the start of a key
  //     rotation. (Assertion: NoStartWhenLocked_A)

  `ASSERT(NotBusyAndDone_A, !((done_core | locking) && busy_execute_d))
  `ASSERT(NoStartWhenLocked_A,
          locking |=> !($rose(busy_execute_d) ||
                        $rose(otbn_dmem_scramble_key_req_busy) ||
                        $rose(otbn_imem_scramble_key_req_busy)))

  // CTRL register
  assign software_errs_fatal_d =
    reg2hw.ctrl.qe && (status_q == StatusIdle) ? reg2hw.ctrl.q :
                                                 software_errs_fatal_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      software_errs_fatal_q <= 1'b0;
    end else begin
      software_errs_fatal_q <= software_errs_fatal_d;
    end
  end

  assign hw2reg.ctrl.d = software_errs_fatal_q;

  // ERR_BITS register
  // The error bits for an OTBN operation get stored on the cycle that done is
  // asserted. Software is expected to read them out before starting the next operation.

  assign hw2reg.err_bits.bad_data_addr.d = err_bits_q.bad_data_addr;
  assign hw2reg.err_bits.bad_insn_addr.d = err_bits_q.bad_insn_addr;
  assign hw2reg.err_bits.call_stack.d = err_bits_q.call_stack;
  assign hw2reg.err_bits.illegal_insn.d = err_bits_q.illegal_insn;
  assign hw2reg.err_bits.loop.d = err_bits_q.loop;
  assign hw2reg.err_bits.key_invalid.d = err_bits_q.key_invalid;
  assign hw2reg.err_bits.rnd_rep_chk_fail.d = err_bits_q.rnd_rep_chk_fail;
  assign hw2reg.err_bits.rnd_fips_chk_fail.d = err_bits_q.rnd_fips_chk_fail;
  assign hw2reg.err_bits.imem_intg_violation.d = err_bits_q.imem_intg_violation;
  assign hw2reg.err_bits.dmem_intg_violation.d = err_bits_q.dmem_intg_violation;
  assign hw2reg.err_bits.reg_intg_violation.d = err_bits_q.reg_intg_violation;
  assign hw2reg.err_bits.bus_intg_violation.d = err_bits_q.bus_intg_violation;
  assign hw2reg.err_bits.bad_internal_state.d = err_bits_q.bad_internal_state;
  assign hw2reg.err_bits.illegal_bus_access.d = err_bits_q.illegal_bus_access;
  assign hw2reg.err_bits.lifecycle_escalation.d = err_bits_q.lifecycle_escalation;
  assign hw2reg.err_bits.fatal_software.d = err_bits_q.fatal_software;

  assign err_bits_clear = reg2hw.err_bits.bad_data_addr.qe & is_not_running_q;
  assign err_bits_d = err_bits_clear ? '0 : err_bits;
  assign err_bits_en = err_bits_clear | done_core;

  logic unused_reg2hw_err_bits;

  // Majority of reg2hw.err_bits is unused as write values are ignored, all writes clear the
  // register to 0.
  assign unused_reg2hw_err_bits = ^{reg2hw.err_bits.bad_data_addr.q,
                                    reg2hw.err_bits.bad_insn_addr,
                                    reg2hw.err_bits.call_stack,
                                    reg2hw.err_bits.illegal_insn,
                                    reg2hw.err_bits.loop,
                                    reg2hw.err_bits.key_invalid,
                                    reg2hw.err_bits.rnd_rep_chk_fail,
                                    reg2hw.err_bits.rnd_fips_chk_fail,
                                    reg2hw.err_bits.imem_intg_violation,
                                    reg2hw.err_bits.dmem_intg_violation,
                                    reg2hw.err_bits.reg_intg_violation,
                                    reg2hw.err_bits.bus_intg_violation,
                                    reg2hw.err_bits.bad_internal_state,
                                    reg2hw.err_bits.illegal_bus_access,
                                    reg2hw.err_bits.lifecycle_escalation,
                                    reg2hw.err_bits.fatal_software};

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_bits_q <= '0;
    end else if (err_bits_en) begin
      err_bits_q <= err_bits_d;
    end
  end

  // Latch the recoverable error signal from the core. This will be generated as a pulse some time
  // during the run (and before secure wipe finishes). Collect up this bit, clearing on the start or
  // end of an operation (start_q / done_core, respectively)
  assign recoverable_err_d = (recoverable_err_q | core_recoverable_err) & ~(start_q | done_core);
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      recoverable_err_q <= '0;
    end else begin
      recoverable_err_q <= recoverable_err_d;
    end
  end

  // FATAL_ALERT_CAUSE register. The .de and .d values are equal for each bit, so that it can only
  // be set, not cleared.
`define DEF_FAC_BIT(NAME)                                         \
  assign hw2reg.fatal_alert_cause.``NAME``.d = 1'b1;              \
  assign hw2reg.fatal_alert_cause.``NAME``.de = err_bits.``NAME;

  `DEF_FAC_BIT(fatal_software)
  `DEF_FAC_BIT(lifecycle_escalation)
  `DEF_FAC_BIT(illegal_bus_access)
  `DEF_FAC_BIT(bad_internal_state)
  `DEF_FAC_BIT(bus_intg_violation)
  `DEF_FAC_BIT(reg_intg_violation)
  `DEF_FAC_BIT(dmem_intg_violation)
  `DEF_FAC_BIT(imem_intg_violation)

`undef DEF_FAC_BIT

  // INSN_CNT register
  logic [31:0] insn_cnt;
  logic        insn_cnt_clear;
  logic        unused_insn_cnt_q;
  assign hw2reg.insn_cnt.d = insn_cnt;
  assign insn_cnt_clear = reg2hw.insn_cnt.qe & is_not_running_q;
  // Ignore all write data to insn_cnt. All writes zero the register.
  assign unused_insn_cnt_q = ^reg2hw.insn_cnt.q;

  // Alerts ====================================================================

  logic [NumAlerts-1:0] alert_test;
  assign alert_test[AlertFatal] = reg2hw.alert_test.fatal.q & reg2hw.alert_test.fatal.qe;
  assign alert_test[AlertRecov] = reg2hw.alert_test.recov.q & reg2hw.alert_test.recov.qe;

  logic [NumAlerts-1:0] alerts;
  assign alerts[AlertFatal] = |{err_bits.fatal_software,
                                err_bits.lifecycle_escalation,
                                err_bits.illegal_bus_access,
                                err_bits.bad_internal_state,
                                err_bits.bus_intg_violation,
                                err_bits.reg_intg_violation,
                                err_bits.dmem_intg_violation,
                                err_bits.imem_intg_violation};

  assign alerts[AlertRecov] = (core_recoverable_err | recoverable_err_q) & done_core;

  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i == AlertFatal)
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni       (rst_n),
      .alert_test_i (alert_test[i]),
      .alert_req_i  (alerts[i]),
      .alert_ack_o  (),
      .alert_state_o(),
      .alert_rx_i   (alert_rx_i[i]),
      .alert_tx_o   (alert_tx_o[i])
    );
  end


  // EDN Connections ============================================================
  logic edn_rnd_req, edn_rnd_ack;
  logic [EdnDataWidth-1:0] edn_rnd_data;
  logic edn_rnd_fips, edn_rnd_err;

  logic edn_urnd_req, edn_urnd_ack;
  logic [EdnDataWidth-1:0] edn_urnd_data;

  // These synchronize the data coming from EDN and stack the 32 bit EDN words to achieve an
  // internal entropy width of 256 bit.

  prim_edn_req #(
    .EnRstChks(1'b1),
    .OutWidth(EdnDataWidth),
    // SEC_CM: RND.BUS.CONSISTENCY
    .RepCheck(1'b1)
  ) u_prim_edn_rnd_req (
    .clk_i,
    .rst_ni     ( rst_n        ),
    .req_chk_i  ( 1'b1         ),
    .req_i      ( edn_rnd_req  ),
    .ack_o      ( edn_rnd_ack  ),
    .data_o     ( edn_rnd_data ),
    .fips_o     ( edn_rnd_fips ),
    .err_o      ( edn_rnd_err  ),
    .clk_edn_i,
    .rst_edn_ni,
    .edn_o      ( edn_rnd_o ),
    .edn_i      ( edn_rnd_i )
  );

  prim_edn_req #(
    .EnRstChks(1'b1),
    .OutWidth(EdnDataWidth)
  ) u_prim_edn_urnd_req (
    .clk_i,
    .rst_ni     ( rst_n         ),
    .req_chk_i  ( 1'b1          ),
    .req_i      ( edn_urnd_req  ),
    .ack_o      ( edn_urnd_ack  ),
    .data_o     ( edn_urnd_data ),
    .fips_o     (               ), // unused
    .err_o      (               ), // unused
    .clk_edn_i,
    .rst_edn_ni,
    .edn_o      ( edn_urnd_o    ),
    .edn_i      ( edn_urnd_i    )
  );


  // OTBN Core =================================================================

  always_ff @(posedge clk_i or negedge rst_n) begin
    if (!rst_n) begin
      busy_execute_q       <= 1'b0;
      init_sec_wipe_done_q <= 1'b0;
    end else begin
      busy_execute_q       <= busy_execute_d;
      init_sec_wipe_done_q <= init_sec_wipe_done_d;
    end
  end
  assign busy_execute_d = (busy_execute_q | start_d) & ~done_core;
  assign init_sec_wipe_done_d = init_sec_wipe_done_q | ~busy_secure_wipe;

  otbn_core #(
    .RegFile(RegFile),
    .DmemSizeByte(DmemSizeByte),
    .ImemSizeByte(ImemSizeByte),
    .RndCnstUrndPrngSeed(RndCnstUrndPrngSeed),
    .SecMuteUrnd(SecMuteUrnd),
    .SecSkipUrndReseedAtStart(SecSkipUrndReseedAtStart)
  ) u_otbn_core (
    .clk_i,
    .rst_ni                      (rst_n),

    .start_i                     (start_q),
    .done_o                      (done_core),
    .locking_o                   (locking),
    .secure_wipe_running_o       (busy_secure_wipe),

    .err_bits_o                  (core_err_bits),
    .recoverable_err_o           (core_recoverable_err),

    .imem_req_o                  (imem_req_core),
    .imem_addr_o                 (imem_addr_core),
    .imem_rdata_i                (imem_rdata_core),
    .imem_rvalid_i               (imem_rvalid_core),

    .dmem_req_o                  (dmem_req_core),
    .dmem_write_o                (dmem_write_core),
    .dmem_addr_o                 (dmem_addr_core),
    .dmem_wdata_o                (dmem_wdata_core),
    .dmem_wmask_o                (dmem_wmask_core),
    .dmem_rmask_o                (dmem_rmask_core_d),
    .dmem_rdata_i                (dmem_rdata_core),
    .dmem_rvalid_i               (dmem_rvalid_core),
    .dmem_rerror_i               (dmem_rerror_core),

    .edn_rnd_req_o               (edn_rnd_req),
    .edn_rnd_ack_i               (edn_rnd_ack),
    .edn_rnd_data_i              (edn_rnd_data),
    .edn_rnd_fips_i              (edn_rnd_fips),
    .edn_rnd_err_i               (edn_rnd_err),

    .edn_urnd_req_o              (edn_urnd_req),
    .edn_urnd_ack_i              (edn_urnd_ack),
    .edn_urnd_data_i             (edn_urnd_data),

    .insn_cnt_o                  (insn_cnt),
    .insn_cnt_clear_i            (insn_cnt_clear),

    .mems_sec_wipe_o             (mems_sec_wipe),
    .dmem_sec_wipe_urnd_key_o    (dmem_sec_wipe_urnd_key),
    .imem_sec_wipe_urnd_key_o    (imem_sec_wipe_urnd_key),
    .req_sec_wipe_urnd_keys_i    (req_sec_wipe_urnd_keys),

    .escalate_en_i               (core_escalate_en),
    .rma_req_i                   (mubi_rma_req),
    .rma_ack_o                   (mubi_rma_ack),

    .software_errs_fatal_i       (software_errs_fatal_q),

    .sideload_key_shares_i       (keymgr_key_i.key),
    .sideload_key_shares_valid_i ({2{keymgr_key_i.valid}})
  );

  always_ff @(posedge clk_i or negedge rst_n) begin
    if (!rst_n) begin
      locking_q <= 1'b0;
    end else begin
      locking_q <= locking;
    end
  end

  // Collect up the error bits that don't come from the core itself and latch them so that they'll
  // be available when an operation finishes.
  assign non_core_err_bits = '{
    lifecycle_escalation: lc_escalate_en[0] != lc_ctrl_pkg::Off,
    illegal_bus_access:   illegal_bus_access_q,
    bad_internal_state:   otbn_scramble_state_error | missed_gnt_error_q | mubi_err,
    bus_intg_violation:   bus_intg_violation
  };

  assign non_core_err_bits_d = non_core_err_bits_q | non_core_err_bits;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      non_core_err_bits_q <= '0;
    end else begin
      non_core_err_bits_q <= non_core_err_bits_d;
    end
  end

  // Construct a full set of error bits from the core output
  assign err_bits = '{
    fatal_software:       core_err_bits.fatal_software,
    lifecycle_escalation: non_core_err_bits_d.lifecycle_escalation,
    illegal_bus_access:   non_core_err_bits_d.illegal_bus_access,
    bad_internal_state:   |{core_err_bits.bad_internal_state,
                            non_core_err_bits_d.bad_internal_state},
    bus_intg_violation:   non_core_err_bits_d.bus_intg_violation,
    reg_intg_violation:   core_err_bits.reg_intg_violation,
    dmem_intg_violation:  core_err_bits.dmem_intg_violation,
    imem_intg_violation:  core_err_bits.imem_intg_violation,
    rnd_fips_chk_fail:    core_err_bits.rnd_fips_chk_fail,
    rnd_rep_chk_fail:     core_err_bits.rnd_rep_chk_fail,
    key_invalid:          core_err_bits.key_invalid,
    loop:                 core_err_bits.loop,
    illegal_insn:         core_err_bits.illegal_insn,
    call_stack:           core_err_bits.call_stack,
    bad_insn_addr:        core_err_bits.bad_insn_addr,
    bad_data_addr:        core_err_bits.bad_data_addr
  };

  // Internally, OTBN uses MUBI types.
  mubi4_t mubi_escalate_en;
  assign mubi_escalate_en = lc_ctrl_pkg::lc_to_mubi4(lc_escalate_en[1]);

  // An error signal going down into the core to show that it should locally escalate
  assign core_escalate_en = mubi4_or_hi(
      mubi4_bool_to_mubi(|{non_core_err_bits.illegal_bus_access,
                           non_core_err_bits.bad_internal_state,
                           non_core_err_bits.bus_intg_violation}),
      mubi_escalate_en
  );

  // Signal error if MuBi input signals take on invalid values as this means something bad is
  // happening. The explicit error detection is required as the mubi4_or_hi operations above
  // might mask invalid values depending on other input operands.
  assign mubi_err = mubi4_test_invalid(mubi_escalate_en);

  // The core can never signal a write to IMEM
  assign imem_write_core = 1'b0;


  // Asserts ===================================================================
  for (genvar i = 0; i < LoopStackDepth; ++i) begin : gen_loop_stack_cntr_asserts
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(
      LoopStackCntAlertCheck_A,
      u_otbn_core.u_otbn_controller.u_otbn_loop_controller.g_loop_counters[i].u_loop_count,
      alert_tx_o[AlertFatal]
    )
  end

  // GPR assertions for secure wipe
  // 1. urnd_reseed_err disables the assertion because secure wipe finishes with failure and OTBN
  // goes to LOCKED state immediately after this error which means that it's not guaranteed to have
  // secure wiping complete.
  // 2. mubi_err_d of start_stop_control disables the internal secure wipe related assertion
  // because a fatal error affecting internal secure wiping could cause an immediate locking
  // behaviour in which it's not guaranteed to see a succesful secure wipe.
  for (genvar i = 2; i < NGpr; ++i) begin : gen_sec_wipe_gpr_asserts
    // Initial secure wipe needs to initialise all registers to nonzero
    `ASSERT(InitSecWipeNonZeroBaseRegs_A,
      $fell(busy_secure_wipe) |->
      u_otbn_core.u_otbn_rf_base.gen_rf_base_ff.u_otbn_rf_base_inner.g_rf_flops[i].rf_reg_q !=
        EccZeroWord,
      clk_i,
      !rst_ni || u_otbn_core.urnd_reseed_err || u_otbn_core.u_otbn_start_stop_control.mubi_err_d)
    // After execution, it's expected to see a change resulting with a nonzero register value
    `ASSERT(SecWipeChangedBaseRegs_A,
      $rose(busy_secure_wipe) |-> ((##[0:$]
        u_otbn_core.u_otbn_rf_base.gen_rf_base_ff.u_otbn_rf_base_inner.g_rf_flops[i].rf_reg_q !=
          EccZeroWord &&
        $changed(
          u_otbn_core.u_otbn_rf_base.gen_rf_base_ff.u_otbn_rf_base_inner.g_rf_flops[i].rf_reg_q))
        within ($rose(busy_secure_wipe) ##[0:$] $fell(busy_secure_wipe))),
      clk_i,
      !rst_ni || u_otbn_core.urnd_reseed_err || u_otbn_core.u_otbn_start_stop_control.mubi_err_d)
  end

  // WDR assertions for secure wipe
  // 1. urnd_reseed_err disables the assertion because secure wipe finishes with failure and OTBN
  // goes to LOCKED state immediately after this error which means that it's not guaranteed to have
  // secure wiping complete.
  // 2. mubi_err_d of start_stop_control disables the internal secure wipe related assertion
  // because a fatal error affecting internal secure wiping could cause an immediate locking
  // behaviour in which it's not guaranteed to see a succesful secure wipe.
  for (genvar i = 0; i < NWdr; ++i) begin : gen_sec_wipe_wdr_asserts
    // Initial secure wipe needs to initialise all registers to nonzero
    `ASSERT(InitSecWipeNonZeroWideRegs_A,
            $fell(busy_secure_wipe) |->
              u_otbn_core.u_otbn_rf_bignum.gen_rf_bignum_ff.u_otbn_rf_bignum_inner.rf[i] !=
                EccWideZeroWord,
            clk_i,
            !rst_ni || u_otbn_core.urnd_reseed_err ||
              u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

    // After execution, it's expected to see a change resulting with a nonzero register value
    `ASSERT(SecWipeChangedWideRegs_A,
            $rose(busy_secure_wipe) |-> ((##[0:$]
              u_otbn_core.u_otbn_rf_bignum.gen_rf_bignum_ff.u_otbn_rf_bignum_inner.rf[i] !=
                EccWideZeroWord &&
              $changed(
                u_otbn_core.u_otbn_rf_bignum.gen_rf_bignum_ff.u_otbn_rf_bignum_inner.rf[i]))
              within ($rose(busy_secure_wipe) ##[0:$] $fell(busy_secure_wipe))),
          clk_i, !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)
  end

  // Secure wipe needs to invalidate call and loop stack, initialize MOD, ACC to nonzero and set
  // FLAGS CSR to zero
  // 1. urnd_reseed_err disables the assertion because secure wipe finishes with failure and OTBN
  // goes to LOCKED state immediately after this error which means that it's not guaranteed to have
  // secure wiping complete.
  // 2. mubi_err_d of start_stop_control disables the secure wipe related assertions because a
  // fatal error affecting internal secure wiping could cause an immediate locking behaviour
  // in which it's not guaranteed to see a succesful secure wipe.
  `ASSERT(SecWipeInvalidCallStack_A,
          $fell(busy_secure_wipe) |-> (!u_otbn_core.u_otbn_rf_base.u_call_stack.top_valid_o),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)
  `ASSERT(SecWipeInvalidLoopStack_A,
          $fell(busy_secure_wipe) |->
            (!u_otbn_core.u_otbn_controller.u_otbn_loop_controller.loop_info_stack.top_valid_o),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

  `ASSERT(SecWipeNonZeroMod_A,
          $fell(busy_secure_wipe) |-> u_otbn_core.u_otbn_alu_bignum.mod_intg_q != EccWideZeroWord,
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

  `ASSERT(SecWipeNonZeroACC_A,
          $fell(busy_secure_wipe) |->
            u_otbn_core.u_otbn_alu_bignum.ispr_acc_intg_i != EccWideZeroWord,
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

  `ASSERT(SecWipeNonZeroFlags_A,
          $fell(busy_secure_wipe) |-> (!u_otbn_core.u_otbn_alu_bignum.flags_flattened),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

  // Secure wipe of IMEM and DMEM first happens with a key change from URND (while valid is zero)
  `ASSERT(ImemSecWipeRequiresUrndKey_A,
          $rose(imem_sec_wipe) |=> (otbn_imem_scramble_key == $past(imem_sec_wipe_urnd_key)),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)
  `ASSERT(DmemSecWipeRequiresUrndKey_A,
          $rose(dmem_sec_wipe) |=> (otbn_dmem_scramble_key == $past(dmem_sec_wipe_urnd_key)),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

  // Then it is guaranteed to have a valid key from OTP interface which is different from URND key
  `ASSERT(ImemSecWipeRequiresOtpKey_A,
          $rose(imem_sec_wipe) ##1 (otbn_imem_scramble_key == $past(imem_sec_wipe_urnd_key)) |=>
            ##[0:$] otbn_imem_scramble_valid && $changed(otbn_imem_scramble_key),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)
  `ASSERT(DmemSecWipeRequiresOtpKey_A,
          $rose(dmem_sec_wipe) ##1 (otbn_dmem_scramble_key == $past(dmem_sec_wipe_urnd_key)) |=>
            ##[0:$] otbn_dmem_scramble_valid && $changed(otbn_dmem_scramble_key),
          clk_i,
          !rst_ni || u_otbn_core.urnd_reseed_err ||
            u_otbn_core.u_otbn_start_stop_control.mubi_err_d)

  // All outputs should be known value after reset
  `ASSERT_KNOWN(TlODValidKnown_A, tl_o.d_valid)
  `ASSERT_KNOWN(TlOAReadyKnown_A, tl_o.a_ready)
  `ASSERT_KNOWN(IdleOKnown_A, idle_o)
  `ASSERT_KNOWN(IntrDoneOKnown_A, intr_done_o)
  `ASSERT_KNOWN(AlertTxOKnown_A, alert_tx_o)
  `ASSERT_KNOWN(EdnRndOKnown_A, edn_rnd_o, clk_edn_i, !rst_edn_ni)
  `ASSERT_KNOWN(EdnUrndOKnown_A, edn_urnd_o, clk_edn_i, !rst_edn_ni)
  `ASSERT_KNOWN(OtbnOtpKeyO_A, otbn_otp_key_o, clk_otp_i, !rst_otp_ni)
  `ASSERT_KNOWN(ErrBitsKnown_A, err_bits)

  // Incoming key must be valid (other inputs go via prim modules that handle the X checks).
  `ASSERT_KNOWN(KeyMgrKeyValid_A, keymgr_key_i.valid)

  // In locked state, the readable registers INSN_CNT, IMEM, and DMEM are expected to always read 0
  // when accessed from the bus. For INSN_CNT, we use "|=>" so that the assertion lines up with
  // "status.q" (a signal that isn't directly accessible here).
  `ASSERT(LockedInsnCntReadsZero_A, (hw2reg.status.d == StatusLocked) |=> insn_cnt == 'd0)
  `ASSERT(ExecuteOrLockedImemReadsZero_A,
          (hw2reg.status.d inside {StatusBusyExecute, StatusLocked}) & imem_rvalid_bus
          |-> imem_rdata_bus == 'd0)
  `ASSERT(ExecuteOrLockedDmemReadsZero_A,
          (hw2reg.status.d inside {StatusBusyExecute, StatusLocked}) & dmem_rvalid_bus
          |-> dmem_rdata_bus == 'd0)

  // From the cycle the core is told to start to when it is done, it must always be busy executing,
  // locking, or both -- even if the core is never done.  We use this property to enable blanking
  // while the core is executing or locking, and this assertion ensures that there is no gap
  // between execution and locking.
  `ASSERT(BusyOrLockingFromStartToDone_A,
          $rose(start_q) |-> (busy_execute_d | locking) |-> ##[0:$] $rose(done_core))

  // Error handling: if we pass an error signal down to the core then we should also be setting an
  // error flag. Note that this uses err_bits, not err_bits_q, because the latter signal only gets
  // asserted when an operation finishes.
  `ASSERT(ErrBitIfEscalate_A, mubi4_test_true_loose(core_escalate_en) |=> |err_bits)

  // Constraint from package, check here as we cannot have `ASSERT_INIT in package
  `ASSERT_INIT(WsrESizeMatchesParameter_A, $bits(wsr_e) == WsrNumWidth)

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(OtbnStartStopFsmCheck_A,
    u_otbn_core.u_otbn_start_stop_control.u_state_regs, alert_tx_o[AlertFatal])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(OtbnControllerFsmCheck_A,
    u_otbn_core.u_otbn_controller.u_state_regs, alert_tx_o[AlertFatal])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(OtbnScrambleCtrlFsmCheck_A,
    u_otbn_scramble_ctrl.u_state_regs, alert_tx_o[AlertFatal])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(OtbnCallStackWrPtrAlertCheck_A,
    u_otbn_core.u_otbn_rf_base.u_call_stack.u_stack_wr_ptr, alert_tx_o[AlertFatal])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(OtbnLoopInfoStackWrPtrAlertCheck_A,
    u_otbn_core.u_otbn_controller.u_otbn_loop_controller.loop_info_stack.u_stack_wr_ptr,
    alert_tx_o[AlertFatal])

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A,
      u_reg, alert_tx_o[AlertFatal])
  // other onehot checks
  `ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ALERT(RfBaseOnehotCheck_A,
      u_otbn_core.u_otbn_rf_base.gen_rf_base_ff.u_otbn_rf_base_inner.u_prim_onehot_check,
      alert_tx_o[AlertFatal])
  `ASSERT_PRIM_ONEHOT_ERROR_TRIGGER_ALERT(RfBignumOnehotCheck_A,
      u_otbn_core.u_otbn_rf_bignum.gen_rf_bignum_ff.u_otbn_rf_bignum_inner.u_prim_onehot_check,
      alert_tx_o[AlertFatal])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(DmemFifoWptrCheck_A,
      u_tlul_adapter_sram_dmem.u_rspfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_wptr,
      alert_tx_o[AlertFatal])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(DmemFifoRptrCheck_A,
      u_tlul_adapter_sram_dmem.u_rspfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_rptr,
      alert_tx_o[AlertFatal])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(ImemFifoWptrCheck_A,
      u_tlul_adapter_sram_imem.u_rspfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_wptr,
      alert_tx_o[AlertFatal])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(ImemFifoRptrCheck_A,
      u_tlul_adapter_sram_imem.u_rspfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_rptr,
      alert_tx_o[AlertFatal])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// sha3_pkg

package sha3_pkg;

  // StateW represents the width of Keccak state variable.
  // As Sha3 assume the state value as 1600, this shouldn't be modified.
  // Note that keccak_round is flexible. It can have any values defined in SHA3
  // specification. But sha3pad logic assumes the value as 1600.
  parameter int StateW = 1600;

  // Function Name (N) and Customzation String (S) shall be
  // smaller than 2**256 bits and integer divisiable by 8.
  parameter int FnWidth = 32;  // up to 32bit Function Name
  parameter int CsWidth = 256; // up to 256bit Customization Input

  // Calculate left_encode(len( X )) bit size.
  // Assume the enc_8(n) is always 1 (up to 255 byte of len(S) size)
  // e.g) 248bit --> two bytes , 256bit --> three bytes
  //  round8bit(clog2(X+1))/8

  parameter int MaxFnEncodeSize = ($clog2(FnWidth+1) + 8 - 1) / 8 + 1;
  parameter int MaxCsEncodeSize = ($clog2(CsWidth+1) + 8 - 1) / 8 + 1;

  parameter int NSRegisterSizePre = FnWidth/8       + CsWidth/8
                                  + MaxFnEncodeSize + MaxCsEncodeSize;
  // Round up to 32bit word base
  parameter int NSRegisterSize = ((NSRegisterSizePre + 4 - 1 ) / 4) * 4;

  // Prefix represents bytepad(encode_string(N) || encode_string(S), 168 or 136)
  // +2 represents left_encoding(168 or 136) which could be either:
  // 10000000 || 00010101 // 168
  // 10000000 || 00010001 // 136
  parameter int PrefixSize = NSRegisterSize + 2;

  // index width for `N` and `S`
  parameter int PrefixIndexW = $clog2(PrefixSize/64);

  // Datapath width in KMAC, this also affects the output of MSG_FIFO
  // This is assumed as 64 in KMAC design. If this value is changed, some parts
  // of the KMAC design need to be changed.
  //
  // 1. keccak_round logic datapath. Keccak round logic assumes MsgWidth
  //    divides 1600 keccak state `Width`. Choose the value accordingly.
  // 2. sha3pad module has fixed width mux for funcpad logic. If MsgWidth is
  //    changed, the logic also need to be revised.
  // 3. kmac core logic also has fixed size mux for appeding output length.
  //    Revise the case statement to fit into revised MsgWidth value.
  parameter int MsgWidth = 64;
  parameter int MsgStrbW = MsgWidth / 8;

  // Keccak module supports SHA3, SHAKE, cSHAKE function.
  // This mode determines if the module uses encoded N and S or not.
  // Also it chooses the padding value.
  //
  //    mode   |  little-endian
  //    -------|----------------
  //    Sha3   |  2'b   10
  //    Shake  |  4'b 1111
  //    CShake |  2'b   00
  //
  // Please remind that if input strings N and S are empty, SW shall
  // choose SHAKE even for cSHAKE operation.
  typedef enum logic[1:0] {
    Sha3   = 2'b 00,
    Shake  = 2'b 10,
    CShake = 2'b 11
  } sha3_mode_e;

  // keccak_strength_e determines the security strength against collision attack
  // This value decides the _rate_ and _capacity_ of the keccak states.
  // It affects the sha3pad module too. the padding module implements
  // `bytepad(X,168)` for L128, `bytepad(X,136)` for L256 in cSHAKE
  typedef enum logic [2:0] {
    L128 = 3'b 000, // rate: 1344 bit / capacity:  256 bit Keccak[ 256](, 128)
    L224 = 3'b 001, // rate: 1152 bit / capacity:  448 bit Keccak[ 448](, 224)
    L256 = 3'b 010, // rate: 1088 bit / capacity:  512 bit Keccak[ 512](, 256)
    L384 = 3'b 011, // rate:  832 bit / capacity:  768 bit Keccak[ 768](, 384)
    L512 = 3'b 100  // rate:  576 bit / capacity: 1024 bit Keccak[1024](, 512)
  } keccak_strength_e;

  parameter int unsigned KeccakRate [5] = '{
    1344/MsgWidth,  // 21 depth := (1600 - 128*2)
    1152/MsgWidth,  // 18 depth := (1600 - 224*2)
    1088/MsgWidth,  // 17 depth := (1600 - 256*2)
     832/MsgWidth,  // 13 depth := (1600 - 384*2)
     576/MsgWidth   //  9 depth := (1600 - 512*2)
  };

  parameter int unsigned KeccakBitCapacity [5] = '{
    2 * 128, // capacity for L128
    2 * 224, // capacity for L224
    2 * 256, // capacity for L256
    2 * 384, // capacity for L384
    2 * 512  // capacity for L512
  };

  parameter int unsigned MaxBlockSize = KeccakRate[0];

  parameter int unsigned KeccakEntries = 1600/MsgWidth;
  parameter int unsigned KeccakMsgAddrW = $clog2(KeccakEntries);

  parameter int unsigned KeccakCountW = $clog2(KeccakEntries+1);

  // SHA3 core state. This state value is used in sha3core module
  // and also in KMAC top module and the register interface for sw to track the
  // sha3 status.
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 7 -n 6 \
  //      -s 4082450958 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (57.14%)
  //  4: ||||||||||||||| (42.86%)
  //  5: --
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4
  //
  localparam int StateWidth = 6;
  typedef enum logic [StateWidth-1:0] {
    StIdle_sparse = 6'b101100,

    // Absorb stage receives the message bitstream and computes the keccak
    // rounds. This internal operation is mainly done inside sha3pad module
    // not sha3core. The core module and this state machine observe the status
    // of the process and mainly waits until all the sponge absorbing is
    // completed. The main indicator is `absorbed` signal.
    StAbsorb_sparse = 6'b100001,

    // Reserved state for context-switching. See #3479.
    // Abort stage can be moved from StAbsorb stage. It basically holds the
    // keccak round operation and opens up the internal state variable to the
    // software. This stage is for the software to pause current operation and
    // store the internal state elsewhere then initiates new KMAC/SHA3 process.
    // StAbort only can be moved to _StFlush_.
    //StAbort_sparse = 6'b011101,

    // Squeeze stage allows the software to read the internal state.
    // If `EnMasking`, it opens the read permission of two share of the state.
    // The squeezing in SHA3 specification describes the software to read up to
    // the rate of SHA3 algorithm but this logic opens up the entire 1600 bits
    // of the state (3200bits if `EnMasking`).
    StSqueeze_sparse = 6'b001011,

    // ManualRun stage initiaties the keccak round and waits the completion.
    // This state is moved from Squeeze state by writing 1 to manual_run CSR.
    // When keccak round is completed, it goes back to Squeeze state.
    StManualRun_sparse = 6'b010000,

    // Flush stage, the core clears out the internal variables and also
    // submodules' variables too. Then moves back to Idle state.
    StFlush_sparse =  6'b000110,

    StTerminalError_sparse = 6'b111010
  } sha3_st_sparse_e;

  localparam int StateWidthLogic = 3;
  typedef enum logic [StateWidthLogic-1:0] {
    StIdle,
    StAbsorb,
    //StAbort,
    StSqueeze,
    StManualRun,
    StFlush,
    StError
  } sha3_st_e;

  function automatic sha3_st_e sparse2logic(sha3_st_sparse_e st);
    unique case (st)
      StIdle_sparse      : return StIdle;
      StAbsorb_sparse    : return StAbsorb;
      //StAbort_sparse   : return StAbort;
      StSqueeze_sparse   : return StSqueeze;
      StManualRun_sparse : return StManualRun;
      StFlush_sparse     : return StFlush;
      default            : return StError;
    endcase
  endfunction : sparse2logic


  //////////////////////
  // Keccak Round FSM //
  //////////////////////

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 8 -n 6 \
  //      -s 1363425333 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (57.14%)
  //  4: ||||||||||||||| (42.86%)
  //  5: --
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 5
  //
  localparam int KeccakFsmWidth = 6;
  typedef enum logic [KeccakFsmWidth-1:0] {
    KeccakStIdle = 6'b011111,

    // Active state is used in Unmasked version only.
    // It handles keccak round in a cycle
    KeccakStActive = 6'b000100,

    // Phase1 --> Phase2Cycle1 --> Phase2Cycle2 --> Phase2Cycle3
    // Activated only in Masked version.
    // Phase1 processes Theta, Rho, Pi steps in a cycle and stores the states
    // into storage. It only moves to Phase2 once the randomness required for
    // Phase2 is available.
    KeccakStPhase1 = 6'b101101,

    // Chi Stage 1 for first lane halves. Unconditionally move to Phase2Cycle2.
    KeccakStPhase2Cycle1 = 6'b000011,

    // Chi Stage 2 and Iota for first lane halves. Chi Stage 1 for second
    // lane halves. We only move forward if the fresh randomness required for
    // remasking is available. Otherwise, keep computing Phase2Cycle1.
    KeccakStPhase2Cycle2 = 6'b011000,

    // Chi Stage 2 and Iota for second lane halves.
    // This state doesn't require random value as it is XORed into the states
    // in Phase1 and Phase2Cycle2. When doing the last round (MaxRound -1)
    // it completes the process and goes back to Idle. If not, it repeats
    // the phases again.
    KeccakStPhase2Cycle3 = 6'b101010,

    // Error state. Not clearly defined yet.
    // Intention is if any unexpected input in the process, state moves to
    // here and report through the error fifo with debugging information.
    KeccakStError = 6'b110001,

    KeccakStTerminalError = 6'b110110
  } keccak_st_e;


  //////////////////
  // Error Report //
  //////////////////
  typedef enum logic [7:0] {
    ErrNone = 8'h 00,

    // ErrSha3SwControl occurs when software sent wrong flow signal.
    // e.g) Sw set `process_i` without `start_i`. The state machine ignores
    //      the signal and report through the error FIFO.
    ErrSha3SwControl = 8'h 80
  } err_code_e;

  typedef struct packed {
    logic        valid;
    err_code_e   code; // Type of error
    logic [23:0] info; // Additional Debug info
  } err_t;


  ///////////////
  // Functions //
  ///////////////

  // Bytepading function
  // `encode_bytepad_len` represents the first two bytes of bytepad()
  // It depends on the block size. We can reuse KeccakRate
  // 10000000 || 00010101 // 168
  // 10000000 || 00010001 // 136
  function automatic logic [15:0] encode_bytepad_len(keccak_strength_e kstrength);
    logic [15:0] result;
    unique case (kstrength)
      L128: result = 16'h A801; // cSHAKE128
      L224: result = 16'h 9001; // not used
      L256: result = 16'h 8801; // cSHAKE256
      L384: result = 16'h 6801; // not used
      L512: result = 16'h 4801; // not used

      default: result = 16'h 0000;
    endcase
    return result;
  endfunction : encode_bytepad_len


endpackage : sha3_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Keccak full round logic based on given input `Width`
// e.g. Width 800 requires 22 rounds

`include "prim_assert.sv"

module keccak_round
  import prim_mubi_pkg::*;
#(
  parameter int Width = 1600, // b= {25, 50, 100, 200, 400, 800, 1600}

  // Derived
  localparam int W        = Width/25,
  localparam int L        = $clog2(W),
  localparam int MaxRound = 12 + 2*L,           // Keccak-f only
  localparam int RndW     = $clog2(MaxRound+1), // Representing up to MaxRound-1

  // Feed parameters
  parameter  int DInWidth = 64, // currently only 64bit supported
  localparam int DInEntry = Width / DInWidth,
  localparam int DInAddr  = $clog2(DInEntry),

  // Control parameters
  parameter  bit EnMasking = 1'b0,  // Enable SCA hardening, requires Width >= 50
  localparam int Share     = EnMasking ? 2 : 1
) (
  input clk_i,
  input rst_ni,

  // Message Feed
  input                valid_i,
  input [DInAddr-1:0]  addr_i,
  input [DInWidth-1:0] data_i [Share],
  output               ready_o,

  // In-process control
  input                    run_i,  // Pulse signal to initiates Keccak full round
  input                    rand_valid_i,
  input                    rand_early_i,
  input      [Width/2-1:0] rand_data_i,
  input                    rand_aux_i,
  output logic             rand_consumed_o,

  output logic             complete_o, // Indicates full round is done

  // State out. This can be used as Digest
  output logic [Width-1:0] state_o [Share],

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  // Errors:
  //  sparse_fsm_error: Checking if FSM state falls into unknown value
  output logic             sparse_fsm_error_o,
  //  round_count_error: prim_count checks round value consistency
  output logic             round_count_error_o,
  //  rst_storage_error: check if reset signal asserted out of the
  //                     permitted window
  output logic             rst_storage_error_o,

  input  prim_mubi_pkg::mubi4_t clear_i     // Clear internal state to '0
);

  import sha3_pkg::*;

  /////////////////////
  // Control signals //
  /////////////////////

  // Update storage register
  logic update_storage;

  // Reset the storage to 0 to initiate new Hash operation
  logic rst_storage;

  // XOR message into storage register
  // It only does based on the given DInWidth.
  // If DInWidth < Width, it takes multiple cycles to XOR all message
  logic xor_message;

  // Select Keccak_p datapath
  // 0: Select Phase1 (Theta -> Rho -> Pi)
  // 1: Select Phase2 (Chi -> Iota)
  // `phase_sel` needs to be asserted until the Chi stage is consumed,
  mubi4_t phase_sel;

  // Cycle index used for controlling input/output muxes and write enables inside
  // keccak_2share.
  logic [1:0] cycle;

  // Increase/ Reset Round number
  logic inc_rnd_num;
  logic rst_rnd_num;

  // Round reaches end
  // This signal indicates the round reaches desired number, which is MaxRound -1.
  // MaxRound is dependant on the Width. In case of SHA3/SHAKE, MaxRound is 24.
  logic rnd_eq_end;

  // Complete of Keccak_f
  // State machine asserts `complete_d` when it reaches at the end of round and
  // operation (Phase3 if Masked). The stage, the storage still doesn't have
  // the valid states. So precisely it is not completed yet.
  // State generated `complete_d` is latched with the clock and creates a pulse
  // signal one cycle later. The signal is the indication of completion.
  //
  // Intentionally removed any intermediate step (so called StComplete) in order
  // to save a clock to proceeds next round.
  logic complete_d;

  //////////////////////
  // Datapath Signals //
  //////////////////////

  // Single round keccak output data
  logic [Width-1:0] keccak_out [Share];

  // Keccak Round indicator: range from 0 .. MaxRound
  logic [RndW-1:0] round;

  // Random value and valid signal used in Keccak_p
  logic               keccak_rand_consumed;
  logic [Width/2-1:0] keccak_rand_data;
  logic               keccak_rand_aux;

  //////////////////////
  // Keccak Round FSM //
  //////////////////////

  // state inputs
  assign rnd_eq_end = (int'(round) == MaxRound - 1);

  keccak_st_e keccak_st, keccak_st_d;
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, keccak_st_d, keccak_st, keccak_st_e, KeccakStIdle)

  // Next state logic and output logic
  // SEC_CM: FSM.SPARSE
  always_comb begin
    // Default values
    keccak_st_d = keccak_st;

    xor_message    = 1'b 0;
    update_storage = 1'b 0;
    rst_storage    = 1'b 0;

    inc_rnd_num = 1'b 0;
    rst_rnd_num = 1'b 0;

    keccak_rand_consumed = 1'b 0;

    phase_sel = MuBi4False;
    cycle = 2'h 0;

    complete_d = 1'b 0;

    sparse_fsm_error_o = 1'b 0;

    unique case (keccak_st)
      KeccakStIdle: begin
        if (valid_i) begin
          // State machine allows Sponge Absorbing only in Idle state.
          keccak_st_d = KeccakStIdle;

          xor_message    = 1'b 1;
          update_storage = 1'b 1;
        end else if (prim_mubi_pkg::mubi4_test_true_strict(clear_i)) begin
          // Opt1. State machine allows resetting the storage only in Idle
          // Opt2. storage resets regardless of states but clear_i
          // Both are added in the design at this time. Will choose the
          // direction later.
          keccak_st_d = KeccakStIdle;

          rst_storage = 1'b 1;
        end else if (EnMasking && run_i) begin
          // Masked version of Keccak handling
          keccak_st_d = KeccakStPhase1;
        end else if (!EnMasking && run_i) begin
          // Unmasked version of Keccak handling
          keccak_st_d = KeccakStActive;
        end else begin
          keccak_st_d = KeccakStIdle;
        end
      end

      KeccakStActive: begin
        // Run Keccak single round logic until it reaches MaxRound - 1
        update_storage = 1'b 1;

        if (rnd_eq_end) begin
          keccak_st_d = KeccakStIdle;

          rst_rnd_num = 1'b 1;
          complete_d  = 1'b 1;
        end else begin
          keccak_st_d = KeccakStActive;

          inc_rnd_num = 1'b 1;
        end
      end

      KeccakStPhase1: begin
        // Theta, Rho and Pi
        phase_sel = MuBi4False;
        cycle =  2'h 0;

        // Only update state and move on once we know the randomness required
        // for Phase2 will be available in the next clock cycle. This way the
        // DOM multipliers inside keccak_2share will be presented the new
        // state (updated with update_storage) at the same time as the new
        // randomness (updated with rand_early_i). Otherwise, stale entropy is
        // paired with fresh data or vice versa. This could lead to undesired
        // SCA leakage.
        if (rand_early_i || rand_valid_i) begin
          keccak_st_d = KeccakStPhase2Cycle1;
          update_storage = 1'b 1;
        end else begin
          keccak_st_d = KeccakStPhase1;
        end
      end

      KeccakStPhase2Cycle1: begin
        // Chi Stage 1 for first lane halves.
        phase_sel = MuBi4True;
        cycle =  2'h 1;

        // Trigger randomness update for next cycle.
        keccak_rand_consumed = 1'b 1;

        // Unconditionally move to next phase/cycle.
        keccak_st_d = KeccakStPhase2Cycle2;
      end

      KeccakStPhase2Cycle2: begin
        // Chi Stage 1 for second lane halves.
        // Chi Stage 2 and Iota for first lane halves.
        phase_sel = MuBi4True;

        // Only update state and move on if the required randomness is
        // available. This way the DOM multipliers inside keccak_2share will be
        // presented the second lane halves at the same time as the new
        // randomness. Otherwise, stale entropy is paired with fresh data or
        // vice versa. This could lead to undesired SCA leakage.
        if (rand_valid_i) begin
          cycle =  2'h 2;

          // Trigger randomness update for next round.
          keccak_rand_consumed = 1'b 1;

          // Update first lane halves.
          update_storage = 1'b 1;

          keccak_st_d = KeccakStPhase2Cycle3;
        end else begin
          cycle =  2'h 1;
          keccak_st_d = KeccakStPhase2Cycle2;
        end
      end

      KeccakStPhase2Cycle3: begin
        // Chi Stage 2 and Iota for second lane halves.
        phase_sel = MuBi4True;
        cycle =  2'h 3;

        // Update second lane halves.
        update_storage = 1'b 1;

        if (rnd_eq_end) begin
          keccak_st_d = KeccakStIdle;

          rst_rnd_num    = 1'b 1;
          complete_d     = 1'b 1;
        end else begin
          keccak_st_d = KeccakStPhase1;

          inc_rnd_num = 1'b 1;
        end
      end

      KeccakStError: begin
        keccak_st_d = KeccakStError;
      end

      KeccakStTerminalError: begin
        //this state is terminal
        keccak_st_d = keccak_st;
        sparse_fsm_error_o = 1'b 1;
      end

      default: begin
        keccak_st_d = KeccakStTerminalError;
        sparse_fsm_error_o = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      keccak_st_d = KeccakStTerminalError;
    end
  end

  // Ready indicates the keccak_round is able to receive new message.
  // While keccak_round is processing the data, it blocks the new message to be
  // XORed into the current state.
  assign ready_o = (keccak_st == KeccakStIdle) ? 1'b 1 : 1'b 0;

  ////////////////////////////
  // Keccak state registers //
  ////////////////////////////

  // SEC_CM: LOGIC.INTEGRITY
  logic rst_n;
  prim_sec_anchor_buf #(
   .Width(1)
  ) u_prim_sec_anchor_buf (
    .in_i(rst_ni),
    .out_o(rst_n)
  );

  logic [Width-1:0] storage   [Share];
  logic [Width-1:0] storage_d [Share];
  always_ff @(posedge clk_i or negedge rst_n) begin
    if (!rst_n) begin
      storage <= '{default:'0};
    end else if (rst_storage) begin
      storage <= '{default:'0};
    end else if (update_storage) begin
      storage <= storage_d;
    end
  end

  assign state_o = storage;

  // Storage register input
  // The incoming message is XORed with the existing storage registers.
  // The logic can accept not a block size incoming message chunk but
  // the size defined in `DInWidth` parameter with its position.

  always_comb begin
    storage_d = keccak_out;
    if (xor_message) begin
      for (int j = 0 ; j < Share ; j++) begin
        for (int unsigned i = 0 ; i < DInEntry ; i++) begin
          // ICEBOX(#18029): handle If Width is not integer divisable by DInWidth
          // Currently it is not allowed to have partial write
          // Please see the Assertion `WidthDivisableByDInWidth_A`
          if (addr_i == i[DInAddr-1:0]) begin
            storage_d[j][i*DInWidth+:DInWidth] =
              storage[j][i*DInWidth+:DInWidth] ^ data_i[j];
          end else begin
            storage_d[j][i*DInWidth+:DInWidth] = storage[j][i*DInWidth+:DInWidth];
          end
        end // for i
      end // for j
    end // if xor_message
  end

  // Check the rst_storage integrity
  logic rst_storage_error;

  always_comb begin : chk_rst_storage
    rst_storage_error = 1'b 0;

    if (rst_storage) begin
      // FSM should be in KeccakStIdle and clear_i should be high
      if ((keccak_st != KeccakStIdle) ||
        prim_mubi_pkg::mubi4_test_false_loose(clear_i)) begin
        rst_storage_error = 1'b 1;
      end
    end
  end : chk_rst_storage

  assign rst_storage_error_o = rst_storage_error ;

  //////////////
  // Datapath //
  //////////////
  keccak_2share #(
    .Width     (Width),
    .EnMasking (EnMasking)
  ) u_keccak_p (
    .clk_i,
    .rst_ni,

    .lc_escalate_en_i,

    .rnd_i           (round),
    .phase_sel_i     (phase_sel),
    .cycle_i         (cycle),
    .rand_aux_i      (keccak_rand_aux),
    .rand_i          (keccak_rand_data),
    .s_i             (storage),
    .s_o             (keccak_out)
  );

  // keccak entropy handling
  assign rand_consumed_o = keccak_rand_consumed;

  assign keccak_rand_data = rand_data_i;
  assign keccak_rand_aux = rand_aux_i;

  // Round number
  // This primitive is used to place a hardened counter
  // SEC_CM: CTR.REDUN
  prim_count #(
    .Width(RndW)
  ) u_round_count (
    .clk_i,
    .rst_ni,
    .clr_i(rst_rnd_num),
    .set_i(1'b0),
    .set_cnt_i('0),
    .incr_en_i(inc_rnd_num),
    .decr_en_i(1'b0),
    .step_i(RndW'(1)),
    .cnt_o(round),
    .cnt_next_o(),
    .err_o(round_count_error_o)
  );

  // completion signal
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      complete_o <= 1'b 0;
    end else begin
      complete_o <= complete_d;
    end
  end

  ////////////////
  // Assertions //
  ////////////////

  // Only allow `DInWidth` that `Width` is integer divisable by `DInWidth`
  `ASSERT_INIT(WidthDivisableByDInWidth_A, (Width % DInWidth) == 0)

  // If `run_i` triggerred, it shall complete
  //`ASSERT(RunResultComplete_A, run_i ##[MaxRound:] complete_o, clk_i, !rst_ni)

  // valid_i and run_i cannot be asserted at the same time
  `ASSUME(OneHot0ValidAndRun_A, $onehot0({valid_i, run_i}), clk_i, !rst_ni)

  // valid_i, run_i only asserted in Idle state
  `ASSUME(ValidRunAssertStIdle_A, valid_i || run_i |-> keccak_st == KeccakStIdle, clk_i, !rst_ni)

  // clear_i is assumed to be asserted in Idle state
  `ASSUME(ClearAssertStIdle_A,
    prim_mubi_pkg::mubi4_test_true_strict(clear_i)
     |-> keccak_st == KeccakStIdle, clk_i, !rst_ni)

  // EnMasking controls the valid states
  if (EnMasking) begin : gen_mask_st_chk
    `ASSERT(EnMaskingValidStates_A, keccak_st != KeccakStActive, clk_i, !rst_ni)
  end else begin : gen_unmask_st_chk
    `ASSERT(UnmaskValidStates_A, !(keccak_st
        inside {KeccakStPhase1, KeccakStPhase2Cycle1, KeccakStPhase2Cycle2, KeccakStPhase2Cycle3}),
        clk_i, !rst_ni)
  end
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// This module is the single round keccak permutation module
// It supports Keccak with up to 1600b of state

`include "prim_assert.sv"

module keccak_2share
  import prim_mubi_pkg::*;
#(
  parameter int Width = 1600, // b= {25, 50, 100, 200, 400, 800, 1600}

  // Derived
  localparam int W        = Width/25,
  localparam int L        = $clog2(W),
  localparam int MaxRound = 12 + 2*L,           // Keccak-f only
  localparam int RndW     = $clog2(MaxRound+1), // Representing up to MaxRound

  // Control parameters
  parameter  bit EnMasking = 0,                // Enable secure hardening
  localparam int Share     = EnMasking ? 2 : 1
) (
  input clk_i,
  input rst_ni,

  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i, // Used to disable SVAs when escalating.

  input         [RndW-1:0] rnd_i, // Current round index
  input mubi4_t            phase_sel_i, // Output mux contol. Used when EnMasking := 1
  input              [1:0] cycle_i, // Current cycle index. Used when EnMasking := 1
  input                    rand_aux_i, // Auxiliary randomness input. Used when EnMasking := 1
  input      [Width/2-1:0] rand_i, // Randomness for remasking. Used when EnMasking := 1
  input        [Width-1:0] s_i      [Share],
  output logic [Width-1:0] s_o      [Share]
);
  ///////////
  // Types //
  ///////////
  //             x    y    z
  typedef logic [4:0][4:0][W-1:0] box_t;   // (x,y,z) state
  typedef logic           [W-1:0] lane_t;  // (z)
  typedef logic [4:0]     [W-1:0] plane_t; // (x,z)
  typedef logic [4:0][4:0]        slice_t; // (x,y)
  typedef logic      [4:0][W-1:0] sheet_t; // (y,z) identical to plane_t
  typedef logic [4:0]             row_t;   // (x)
  typedef logic      [4:0]        col_t;   // (y) identical to row_t

  //////////////
  // Keccak_f //
  //////////////
  box_t state_in   [Share];
  box_t state_out  [Share];
  box_t theta_data [Share];
  box_t rho_data   [Share];
  box_t pi_data    [Share];
  box_t chi_data   [Share];
  box_t iota_data  [Share];

  box_t phase1_in  [Share];
  box_t phase1_out [Share];
  box_t phase2_in  [Share];
  box_t phase2_out [Share];

  /////////////////
  // Unused nets //
  /////////////////
  // Tie off input signals that aren't used in the unmasked implementation.
  if (!EnMasking) begin : gen_tie_unused
    logic unused_clk;
    logic unused_rst_n;
    mubi4_t unused_phase_sel;
    logic [1:0] unused_cycle;
    logic unused_rand_aux;
    logic [Width/2-1:0] unused_rand;
    assign unused_clk = clk_i;
    assign unused_rst_n = rst_ni;
    assign unused_phase_sel = phase_sel_i;
    assign unused_cycle = cycle_i;
    assign unused_rand_aux = rand_aux_i;
    assign unused_rand = rand_i;
  end

  //////////////////////////////////////////////////
  // Input/output type conversion and interfacing //
  //////////////////////////////////////////////////
  for (genvar i = 0 ; i < Share ; i++) begin : g_state_inout
    assign state_in[i] = bitarray_to_box(s_i[i]);
    assign s_o[i]      = box_to_bitarray(state_out[i]);
  end : g_state_inout

  if (EnMasking) begin : g_2share_data
    assign phase1_in = state_in;
    assign phase2_in = state_in;

    always_comb begin
      unique case (phase_sel_i)
        MuBi4False: state_out = phase1_out;
        MuBi4True:  state_out = phase2_out;
        default:    state_out = phase1_out;
      endcase
    end
  end else begin : g_single_data
    assign phase1_in = state_in;
    assign phase2_in = phase1_out;
    assign state_out = phase2_out;
  end

  //////////////
  // Datapath //
  //////////////
  // This module has two phases. First phase, it calculates Theta, Rho, Pi steps
  // in SHA3. At the second phase, it computes Chi and Iota steps. If masking is
  // not enabled, the two phases are completed within a single clock cycle.
  //
  // If masking is enabled, the first phase (Phase1) completes in one cycle.
  // Then, the output should be stored in the state and given to the input of
  // this module again. The second phase in the masked version needs three
  // clock cycles to complete. In the first clock cycle, the first stage of Chi
  // is computed for the first lane halves. In the second clock cycle, the
  // module then outputs the updated first lane halves. In the third clock
  // cycle, the new second lane halves are output. To aggravate SCA, we
  // randomly decide which lane halves to process first on a per-round basis.
  // We use additional randomness generated by the PRNG to take this decision
  // (rand_aux_i). For more details, refer to the comments in the "MUX control"
  // section below.

  for (genvar i = 0 ; i < Share ; i++) begin : g_datapath

    // Phase 1:
    assign theta_data[i] = theta(phase1_in[i]);
    // Commented out rho function as vcs complains z-Offset%W isn't constant
    // assign rho_data[i]   = rho(theta_data[i]);

    assign pi_data[i]    = pi(rho_data[i]);

    // Phase 2 (Cycles 1, 2 and 3):
    // Chi : See below
    // Iota: See below
  end : g_datapath

  assign phase1_out = pi_data;

  // Iota adds Round Constants(RC), so only one share should be XORed
  if (EnMasking) begin : g_2share_iota
    assign iota_data[0]  = iota(chi_data[0], rnd_i);
    assign iota_data[1]  = chi_data[1];
  end else begin : g_single_iota
    assign iota_data[0]  = iota(chi_data[0], rnd_i);
  end

  if (EnMasking) begin : g_2share_chi
    // Domain-Oriented Masking
    // reference: https://eprint.iacr.org/2017/395.pdf

    localparam int unsigned WSheetHalf = $bits(sheet_t)/2;
    logic [4:0][WSheetHalf-1:0] in_prd, out_prd;

    logic low_then_high_d, low_then_high_q;
    logic in_data_low, out_data_low;
    logic in_rand_ext;
    logic update_dom;

    /////////////////
    // MUX control //
    /////////////////

    // Update lane-half processing order in Phase 1 and keep the value constant
    // for the entire round.
    assign low_then_high_d =
        mubi4_test_false_strict(phase_sel_i) ? rand_aux_i : low_then_high_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        low_then_high_q <= 1'b 0;
      end else begin
        low_then_high_q <= low_then_high_d;
      end
    end

    // This implementation uses both randomness provided from an external PRNG
    // as well as intermediate results for remasking the DOM multipliers below.
    // Per clock cycle, 800b of pseudo-random data (PRD) are required. The
    // following schedule is used to only ever update the input data when also
    // providing fresh randomness and vice versa.
    //
    // Cycle 0: Compute Theta, Rho, Pi - The DOM multipliers are not evaluated
    //          at all: the inputs are driven by the first lane halves (same
    //          values as in Cycle 3). Also the intermediate results we already
    //          had in Cycle 3 didn't change.
    // Cycle 1: Compute first stage of Chi for first lane halves using the DOM
    //          multipliers. We use the fresh randomness provided from the
    //          PRNG for remasking.
    // Cycle 2: Compute second stage of Chi and Iota for first lane halves.
    //          Compute first stage of Chi for second lane halves. We use the
    //          fresh randomness provided from the PRNG for remasking the
    //          DOM multipliers.
    // Cycle 3: Compute second stage of Chi and Iota for second lane halves.
    //          Feed again first lane halves to DOM multiplier inputs (now
    //          the updated values become visible) together with intermediate
    //          results of Cycle 2. Don't update the register stage inside
    //          the DOM multipliers.
    always_comb begin
      unique case (cycle_i)
        2'h0: begin
          in_data_low = low_then_high_q;
          in_rand_ext = 1'b0;
          update_dom  = 1'b0;
        end
        2'h1: begin
          in_data_low = low_then_high_q;
          in_rand_ext = 1'b1;
          update_dom  = 1'b1;
        end
        2'h2: begin
          in_data_low = ~low_then_high_q;
          in_rand_ext = 1'b1;
          update_dom  = 1'b1;
        end
        2'h3: begin
          in_data_low = low_then_high_q;
          in_rand_ext = 1'b0;
          update_dom  = 1'b0;
        end
        default: begin
          in_data_low = low_then_high_q;
          in_rand_ext = 1'b0;
          update_dom  = 1'b0;
        end
      endcase
    end

    // When taking the lower lane halves in, the upper lane halves are output
    // and vice versa.
    assign out_data_low = ~in_data_low;

    /////////////////////
    // DOM multipliers //
    /////////////////////

    for (genvar x = 0 ; x < 5 ; x++) begin : g_chi_w
      localparam int X1 = (x + 1) % 5;
      localparam int X2 = (x + 2) % 5;

      sheet_t sheet0[Share]; // Inverted input X1
      sheet_t sheet1[Share]; // X2
      sheet_t sheet2[Share]; // DOM output

      assign sheet0[0] = ~phase2_in[0][X1];
      assign sheet0[1] = phase2_in[1][X1];

      assign sheet1[0] = phase2_in[0][X2];
      assign sheet1[1] = phase2_in[1][X2];

      // Convert sheet_t to 1D arrays, one for the upper and lower half lane.
      logic [WSheetHalf-1:0] a0_l, a1_l, b0_l, b1_l;
      logic [WSheetHalf-1:0] a0_h, a1_h, b0_h, b1_h;
      logic [WSheetHalf-1:0] a0, a1, b0, b1, q0, q1;

      assign a0_l = {sheet0[0][0][W/2-1:0],
                     sheet0[0][1][W/2-1:0],
                     sheet0[0][2][W/2-1:0],
                     sheet0[0][3][W/2-1:0],
                     sheet0[0][4][W/2-1:0]};
      assign a1_l = {sheet0[1][0][W/2-1:0],
                     sheet0[1][1][W/2-1:0],
                     sheet0[1][2][W/2-1:0],
                     sheet0[1][3][W/2-1:0],
                     sheet0[1][4][W/2-1:0]};

      assign a0_h = {sheet0[0][0][W-1:W/2],
                     sheet0[0][1][W-1:W/2],
                     sheet0[0][2][W-1:W/2],
                     sheet0[0][3][W-1:W/2],
                     sheet0[0][4][W-1:W/2]};
      assign a1_h = {sheet0[1][0][W-1:W/2],
                     sheet0[1][1][W-1:W/2],
                     sheet0[1][2][W-1:W/2],
                     sheet0[1][3][W-1:W/2],
                     sheet0[1][4][W-1:W/2]};

      assign b0_l = {sheet1[0][0][W/2-1:0],
                     sheet1[0][1][W/2-1:0],
                     sheet1[0][2][W/2-1:0],
                     sheet1[0][3][W/2-1:0],
                     sheet1[0][4][W/2-1:0]};
      assign b1_l = {sheet1[1][0][W/2-1:0],
                     sheet1[1][1][W/2-1:0],
                     sheet1[1][2][W/2-1:0],
                     sheet1[1][3][W/2-1:0],
                     sheet1[1][4][W/2-1:0]};

      assign b0_h = {sheet1[0][0][W-1:W/2],
                     sheet1[0][1][W-1:W/2],
                     sheet1[0][2][W-1:W/2],
                     sheet1[0][3][W-1:W/2],
                     sheet1[0][4][W-1:W/2]};
      assign b1_h = {sheet1[1][0][W-1:W/2],
                     sheet1[1][1][W-1:W/2],
                     sheet1[1][2][W-1:W/2],
                     sheet1[1][3][W-1:W/2],
                     sheet1[1][4][W-1:W/2]};

      // Input muxing
      assign a0 = in_data_low ? a0_l : a0_h;
      assign a1 = in_data_low ? a1_l : a1_h;
      assign b0 = in_data_low ? b0_l : b0_h;
      assign b1 = in_data_low ? b1_l : b1_h;

      // Randomness muxing
      // Intermediate results are rotated across rows. The new Row x depends on
      // data from Rows x + 1 and x + 2. Hence we don't want to use intermediate
      // results from Rows x, x + 1, and x + 2 for remasking.
      assign in_prd[x] = in_rand_ext ? rand_i[x * WSheetHalf +: WSheetHalf] :
                                       out_prd[rot_int(x, 5)];

      prim_dom_and_2share #(
        .DW (WSheetHalf), // a half sheet
        .Pipeline(1) // Process the full sheet in 3 clock cycles. This reduces
                     // SCA leakage.
      ) u_dom (
        .clk_i,
        .rst_ni,

        .a0_i      (a0),
        .a1_i      (a1),
        .b0_i      (b0),
        .b1_i      (b1),
        .z_valid_i (update_dom),
        .z_i       (in_prd[x]),
        .q0_o      (q0),
        .q1_o      (q1),
        .prd_o     (out_prd[x])
      );

      // Output conversion from q0, q1 to sheet_t
      // For simplicity, we forward the generated lane half to both the upper
      // and lower lane halves at this point. The actual output muxing/selection
      // happens after the Iota step when generating phase2_out from iota_data
      // and state_in below.
      assign sheet2[0][4] = {2{q0[W/2*0+:W/2]}};
      assign sheet2[0][3] = {2{q0[W/2*1+:W/2]}};
      assign sheet2[0][2] = {2{q0[W/2*2+:W/2]}};
      assign sheet2[0][1] = {2{q0[W/2*3+:W/2]}};
      assign sheet2[0][0] = {2{q0[W/2*4+:W/2]}};

      assign sheet2[1][4] = {2{q1[W/2*0+:W/2]}};
      assign sheet2[1][3] = {2{q1[W/2*1+:W/2]}};
      assign sheet2[1][2] = {2{q1[W/2*2+:W/2]}};
      assign sheet2[1][1] = {2{q1[W/2*3+:W/2]}};
      assign sheet2[1][0] = {2{q1[W/2*4+:W/2]}};

      // Final XOR to generate the output
      assign chi_data[0][x] = sheet2[0] ^ phase2_in[0][x];
      assign chi_data[1][x] = sheet2[1] ^ phase2_in[1][x];
    end : g_chi_w

    // Since Chi and thus Iota are separately applied to the lower and upper half
    // lanes, we need to forward the input to the other half.
    for (genvar x = 0 ; x < 5 ; x++) begin : g_2share_phase2_out_row
      for (genvar y = 0 ; y < 5 ; y++) begin : g_2share_phase2_out_col
        assign phase2_out[0][x][y] = out_data_low ?
            { state_in[0][x][y][W-1:W/2], iota_data[0][x][y][W/2-1:0]} :
            {iota_data[0][x][y][W-1:W/2],  state_in[0][x][y][W/2-1:0]};
        assign phase2_out[1][x][y] = out_data_low ?
            { state_in[1][x][y][W-1:W/2], iota_data[1][x][y][W/2-1:0]} :
            {iota_data[1][x][y][W-1:W/2],  state_in[1][x][y][W/2-1:0]};
      end
    end

  end else begin : g_single_chi
    assign chi_data[0] = chi(phase2_in[0]);
    assign phase2_out = iota_data;
  end

  // Rho ======================================================================
  // As RhoOffset[x][y] is considered as variable int in VCS,
  // it is replaced with generate statement.
  // Revised to meet verilator lint. Now RhoOffset is 1-D array
  localparam int RhoOffset [25]  = '{
    //y  0    1    2    3    4     x
         0,  36,   3, 105, 210, // 0:  0  1  2  3  4
         1, 300,  10,  45,  66, // 1:  5  6  7  8  9
       190,   6, 171,  15, 253, // 2: 10 11 12 13 14
        28,  55, 153,  21, 120, // 3: 15 16 17 18 19
        91, 276, 231, 136,  78  // 4: 20 21 22 23 24
  };
  for (genvar i = 0 ; i < Share ; i++) begin : g_rho
    box_t rho_in, rho_out;
    assign rho_in = theta_data[i];
    assign rho_data[i] = rho_out;

    for (genvar x = 0 ; x < 5 ; x++) begin : gen_rho_x
      for (genvar y = 0 ; y < 5 ; y++) begin : gen_rho_y
        localparam int Offset = RhoOffset[5*x+y]%W;
        localparam int ShiftAmt = W- Offset;
        if (Offset == 0) begin : gen_offset0
          assign rho_out[x][y][W-1:0] = rho_in[x][y][W-1:0];
        end else begin : gen_others
          assign rho_out[x][y][W-1:0] = {rho_in[x][y][0+:ShiftAmt],
                                         rho_in[x][y][ShiftAmt+:Offset]};
        end
      end
    end
  end : g_rho

  ////////////////
  // Assertions //
  ////////////////

  `ASSERT_INIT(ValidWidth_A,
      EnMasking == 0 && Width inside {25, 50, 100, 200, 400, 800, 1600} ||
      EnMasking == 1 && Width inside {50, 100, 200, 400, 800, 1600})
  `ASSERT_INIT(ValidW_A, W inside {1, 2, 4, 8, 16, 32, 64})
  `ASSERT_INIT(ValidL_A, L inside {0, 1, 2, 3, 4, 5, 6})
  `ASSERT_INIT(ValidRound_A, MaxRound <= 24) // Keccak-f only

  // phase_sel_i shall stay for two cycle after change to 1.
  lc_ctrl_pkg::lc_tx_t unused_lc_sig;
  assign unused_lc_sig = lc_escalate_en_i;
  if (EnMasking) begin : gen_selperiod_chk
    `ASSUME(SelStayTwoCycleIfTrue_A,
        ($past(phase_sel_i) == MuBi4False) && (phase_sel_i == MuBi4True)
        |=> phase_sel_i == MuBi4True, clk_i, !rst_ni || lc_escalate_en_i != lc_ctrl_pkg::Off)
  end

  ///////////////
  // Functions //
  ///////////////

  // Convert bitarray to 3D box
  // Please take a look at FIPS PUB 202
  // https://nvlpubs.nist.gov/nistpubs/FIPS/NIST.FIPS.202.pdf
  // > For all triples (x,y,z) such that 0<=x<5, 0<=y<5, and 0<=z<w,
  // >    A[x,y,z]=S[w(5y+x)+z]
  function automatic box_t bitarray_to_box(logic [Width-1:0] s_in);
    automatic box_t box;
    for (int y = 0 ; y < 5 ; y++) begin
      for (int x = 0 ; x < 5 ; x++) begin
        for (int z = 0 ; z < W ; z++) begin
          box[x][y][z] = s_in[W*(5*y+x) + z];
        end
      end
    end
    return box;
  endfunction : bitarray_to_box

  // Convert 3D cube to bitarray
  function automatic logic [Width-1:0] box_to_bitarray(box_t state);
    automatic logic [Width-1:0] bitarray;
    for (int y = 0 ; y < 5 ; y++) begin
      for (int x = 0 ; x < 5 ; x++) begin
        for (int z = 0 ; z < W ; z++) begin
          bitarray[W*(5*y+x)+z] = state[x][y][z];
        end
      end
    end
    return bitarray;
  endfunction : box_to_bitarray

  // Rotate integer indices
  function automatic integer rot_int(integer in, integer num);
    integer out;
    if (in == 0) begin
      out = num - 1;
    end else begin
      out = in - 1;
    end
    return out;
  endfunction

  // Step Mapping =============================================================
  // theta
  // XOR each bit in the state with the parity of two columns
  // C[x,z] = A[x,0,z] ^ A[x,1,z] ^ A[x,2,z] ^ A[x,3,z] ^ A[x,4,z]
  // D[x,z] = C[x-1,z] ^ C[x+1,z-1]
  // theta = A[x,y,z] ^ D[x,z]
  parameter int ThetaIndexX1 [5] = '{4, 0, 1, 2, 3}; // (x-1)%5
  parameter int ThetaIndexX2 [5] = '{1, 2, 3, 4, 0}; // (x+1)%5
  function automatic box_t theta(box_t state);
    plane_t c;
    plane_t d;
    box_t result;
    for (int x = 0 ; x < 5 ; x++) begin
      c[x] = state[x][0] ^ state[x][1] ^ state[x][2] ^ state[x][3] ^ state[x][4];
    end
    for (int x = 0 ; x < 5 ; x++) begin
      for (int z = 0 ; z < W ; z++) begin
        int index_z;
        index_z = (z == 0) ? W-1 : z-1; // (z+1)%W
        d[x][z] = c[ThetaIndexX1[x]][z] ^ c[ThetaIndexX2[x]][index_z];
      end
    end
    for (int x = 0 ; x < 5 ; x++) begin
      for (int y = 0 ; y < 5 ; y++) begin
        result[x][y] = state[x][y] ^ d[x];
      end
    end
    return result;
  endfunction : theta

  // rho

  // Commented out entire rho function due to VCS elaboration error.
  // (z-RhoOffset[x][y]%W) isn't considered as a constant in VCS.
  // Even changing it to W-RhoOffset[x][y]%W and assign to ShiftAmt
  // creates same error.

  // Offset : Look at Table 2 in FIPS PUB 202
  //localparam int RhoOffset [5][5]  = '{
  //  //y  0    1    2    3    4     x
  //  '{   0,  36,   3, 105, 210},// 0
  //  '{   1, 300,  10,  45,  66},// 1
  //  '{ 190,   6, 171,  15, 253},// 2
  //  '{  28,  55, 153,  21, 120},// 3
  //  '{  91, 276, 231, 136,  78} // 4
  //};

  // rotate bits of each lane by offset
  // 1. rho[0,0,z] = A[0,0,z]
  // 2. Offset swap
  //    a. (x,y) := (1,0)
  //    b. for t [0..23]
  //       i. rho[x,y,z] = A[x,y,z-(t+1)(t+2)/2]
  //       ii. (x,y) = (y, (2x+3y))
  //function automatic box_t rho(box_t state);
  //  box_t result;
  //  for (int x = 0 ; x < 5 ; x++) begin
  //    for (int y = 0 ; y < 5 ; y++) begin
  //      for (int z = 0 ; z < W ; z++) begin
  //        automatic int index_z;
  //        index_z = (z-RhoOffset[x][y])%W;
  //        result[x][y][z] = state[x][y][(z-RhoOffset[x][y])%W];
  //      end
  //    end
  //  end
  //  return result;
  //endfunction : rho

  // pi
  // rearrange the position of lanes
  // pi[x,y,z] = state[(x+3y),x,z]
  localparam int PiRotate [5][5] = '{
    //y  0    1    2    3    4     x
    '{   0,   3,   1,   4,   2},// 0
    '{   1,   4,   2,   0,   3},// 1
    '{   2,   0,   3,   1,   4},// 2
    '{   3,   1,   4,   2,   0},// 3
    '{   4,   2,   0,   3,   1} // 4
  };
  function automatic box_t pi(box_t state);
    box_t result;
    for (int x = 0 ; x < 5 ; x++) begin
      for (int y = 0 ; y < 5 ; y++) begin
        result[x][y][W-1:0] = state[PiRotate[x][y]][x][W-1:0];
      end
    end
    return result;
  endfunction : pi

  // chi
  // chi[x,y,z] = state[x,y,z] ^ ((state[x+1,y,z] ^ 1) & state[x+2,y,z])
  parameter int ChiIndexX1 [5] = '{1, 2, 3, 4, 0}; // (x+1)%5
  parameter int ChiIndexX2 [5] = '{2, 3, 4, 0, 1}; // (x+2)%5
  function automatic box_t chi(box_t state);
    box_t result;
    for (int x = 0 ; x < 5 ; x++) begin
      result[x] = state[x] ^ ((~state[ChiIndexX1[x]]) & state[ChiIndexX2[x]]);
    end
    return result;
  endfunction : chi

  // iota
  // XOR (x,y) = (0,0) with Round Constant (RC)

  // RC parameter: Precomputed by util/keccak_rc.py. Only up-to 0..L-1 is used
  // RC = '0
  // RC[2**j-1] = rc(j+7*rnd)
  // rc(t) =
  //    1. t%255 == 0 -> 1
  //    2. R[0:7] = 'b10000000
  //    3. for i = [1..t%255]
  //      a. R = 0 || R
  //      b. R[0] = R[0] ^ R[8]
  //      c. R[4] = R[4] ^ R[8]
  //      d. R[5] = R[5] ^ R[8]
  //      e. R[6] = R[6] ^ R[8]
  //      f. R = R[0:7]
  //    4. return R[0]
  // RC has L = [0..6]
  // for lower L case, only chopping lower part of 64bit RC is sufficient.
  localparam logic [63:0] RC [24] = '{
     64'h 0000_0000_0000_0001, // Round 0
     64'h 0000_0000_0000_8082, // Round 1
     64'h 8000_0000_0000_808A, // Round 2
     64'h 8000_0000_8000_8000, // Round 3
     64'h 0000_0000_0000_808B, // Round 4
     64'h 0000_0000_8000_0001, // Round 5
     64'h 8000_0000_8000_8081, // Round 6
     64'h 8000_0000_0000_8009, // Round 7
     64'h 0000_0000_0000_008A, // Round 8
     64'h 0000_0000_0000_0088, // Round 9
     64'h 0000_0000_8000_8009, // Round 10
     64'h 0000_0000_8000_000A, // Round 11
     64'h 0000_0000_8000_808B, // Round 12
     64'h 8000_0000_0000_008B, // Round 13
     64'h 8000_0000_0000_8089, // Round 14
     64'h 8000_0000_0000_8003, // Round 15
     64'h 8000_0000_0000_8002, // Round 16
     64'h 8000_0000_0000_0080, // Round 17
     64'h 0000_0000_0000_800A, // Round 18
     64'h 8000_0000_8000_000A, // Round 19
     64'h 8000_0000_8000_8081, // Round 20
     64'h 8000_0000_0000_8080, // Round 21
     64'h 0000_0000_8000_0001, // Round 22
     64'h 8000_0000_8000_8008  // Round 23
  };

  // iota: XOR with RC for (x,y) = (0,0)
  function automatic box_t iota(box_t state, logic [RndW-1:0] rnd);
    box_t result;
    result = state;
    result[0][0][W-1:0] = state[0][0][W-1:0] ^ RC[rnd][W-1:0];

    return result;
  endfunction : iota

  // Round function : Rnd(A,i_r)
  // Not used due to rho function issue described above.

  //function automatic box_t keccak_rnd(box_t state, logic [RndW-1:0] rnd);
  //  box_t keccak_state;
  //  keccak_state = iota(chi(pi(rho(theta(state)))), rnd);
  //
  //  return keccak_state;
  //endfunction : keccak_rnd

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SHA3 padding logic

`include "prim_assert.sv"

module sha3pad
  import sha3_pkg::*;
#(
  parameter  bit EnMasking = 0,
  localparam int Share = (EnMasking) ? 2 : 1
) (
  input clk_i,
  input rst_ni,

  // Message interface (FIFO)
  input                       msg_valid_i,
  input        [MsgWidth-1:0] msg_data_i [Share],
  input        [MsgStrbW-1:0] msg_strb_i,         // one strobe for shares
  output logic                msg_ready_o,

  // N, S: Used in cSHAKE mode only
  input [NSRegisterSize*8-1:0] ns_data_i, // See sha3_pkg for details

  // output to keccak_round: message path
  output logic                       keccak_valid_o,
  output logic [KeccakMsgAddrW-1:0]  keccak_addr_o,
  output logic [MsgWidth-1:0]        keccak_data_o [Share],
  input  logic                       keccak_ready_i,

  // keccak_round control and status
  // `run` initiates the keccak_round to process full keccak_f (24rounds).
  // `complete` is an input from keccak round showing the current keccak_f is
  // completed.
  output logic keccak_run_o,
  input        keccak_complete_i,

  // configurations
  input sha3_mode_e       mode_i,
  // strength_i is used in bytepad operation. bytepad() is used in cSHAKE only.
  // SHA3, SHAKE doesn't have encode_N,S
  input keccak_strength_e strength_i,

  // control signal
  // start_i is a pulse signal triggers the padding logic (and the rest of SHA)
  // to accept the incoming messages. This signal is used in the pad module,
  // to initiate the prefix transmitting to keccak_round
  input start_i,
  // process_i is a pulse signal triggers the pad logic to stop receiving the
  // message from MSG_FIFO and pad the trailing bits specified in the SHA3
  // standard. Look at `funcpad` signal for the values.
  input process_i,
  // done_i is a pulse signal to make the pad logic to clear internal variables
  // and to move back to the Idle state for next hashing process.
  // done_i may not needed if sw controls the keccak_round directly.
  input prim_mubi_pkg::mubi4_t done_i,

  // Indication of the Keccak Sponge Absorbing is complete, it is time for SW to
  // control the Keccak-round if it needs more digest, or complete by asserting
  // `done_i`
  output prim_mubi_pkg::mubi4_t absorbed_o,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  // Indication that there was a fault in the sparse encoding
  output logic sparse_fsm_error_o,

  // Indication that there was a fault in the counter
  output logic msg_count_error_o
);

  /////////////////
  // Definitions //
  /////////////////

  // Padding States
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 10 -n 7 \
  //      -s 1116691466 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (42.22%)
  //  4: |||||||||||||||||| (40.00%)
  //  5: ||||| (11.11%)
  //  6: || (4.44%)
  //  7: | (2.22%)
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 7
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 5
  //
  localparam int StateWidthPad = 7;
  typedef enum logic [StateWidthPad-1:0] {
    StPadIdle = 7'b1000010,

    // Sending a block of prefix, if cSHAKE mode is turned on. For the rest
    // (SHA3, SHAKE), sending prefix is not needed. FSM moves from Idle to
    // Message directly in that case.
    //
    // As prim_slicer is instantiated, zerofill after the actual prefix is done
    // by the module.
    StPrefix = 7'b0111100,
    StPrefixWait =7'b1001100,

    // Sending Message. In this state, it directly forwards the incoming data
    // to Keccak round module. If `process_i` is asserted, then the rest of the
    // messages will be discarded until new `start_i` is asserted.
    //
    // The incoming data can be partial write. Padding logic counts the number
    // of bytes received and pause if a block size is transferred.
    StMessage = 7'b0100101,
    StMessageWait = 7'b0001111,

    // After sending the messages, then `process_i` is set, the FSM pads at the
    // end of the message based on `mode_i`. If this is the last byte of the
    // block, then it pads [7] to 1 to complete `pad10*1()` function.
    StPad = 7'b1111010,
    StPadRun = 7'b0011001,

    // If the padding isn't the end of the block byte (which will be rare case),
    // FSM moves to another zerofill state. In contrast to StZerofill, this state
    StPad01 = 7'b1101001,

    // Flushing the internal packers in front of the Keccak data output port.
    StPadFlush = 7'b1010111,

    StTerminalError = 7'b0110011
  } pad_st_e;

  typedef enum logic [2:0] {
    MuxNone    = 3'b 000,
    MuxFifo    = 3'b 001,
    MuxPrefix  = 3'b 010,
    MuxFuncPad = 3'b 011,
    MuxZeroEnd = 3'b 100
  } mux_sel_e;

  ////////////////////
  // Configurations //
  ////////////////////

  logic [KeccakCountW-1:0] block_addr_limit;

  // Block size based on the address.
  // This is used for bytepad() and also pad10*1()
  // assign block_addr_limit = KeccakRate[strength_i];
  // but below is easier to understand
  always_comb begin
    unique case (strength_i)
      L128: block_addr_limit = KeccakCountW'(KeccakRate[L128]);
      L224: block_addr_limit = KeccakCountW'(KeccakRate[L224]);
      L256: block_addr_limit = KeccakCountW'(KeccakRate[L256]);
      L384: block_addr_limit = KeccakCountW'(KeccakRate[L384]);
      L512: block_addr_limit = KeccakCountW'(KeccakRate[L512]);

      default: block_addr_limit = '0;
    endcase
  end

  /////////////////////
  // Control Signals //
  /////////////////////

  // `sel_mux` selects the output data among the incoming or internally generated data.
  // MuxFifo:    data from external (msg_data_i)
  // MuxPrefix:  bytepad(encode_string(N)||encode_string(S), )
  // MuxFuncPad: function_pad with end of message
  // MuxZeroEnd: all 0
  mux_sel_e sel_mux;

  // `sent_message` indicates the number of entries sent to keccak round per
  // block. The value shall be enough to cover Maximum entry of the Keccak
  // storage as defined in sha3_pkg, `$clog2(KeccakEntries+1)`. Logically,
  // it is not needed to have more than KeccakEntries but for safety in case of
  // SHA3 context switch resuming the SHA3 from the middle of sponge
  // construction. If needed, the software should be able to write whole 1600
  // bits. The `sent_message` is used to check sent_blocksize.
  logic [KeccakCountW-1:0] sent_message;
  logic inc_sentmsg, clr_sentmsg;

  // This primitive is used to place a hardened counter
  // SEC_CM: CTR.REDUN
  prim_count #(
    .Width(KeccakCountW)
  ) u_sentmsg_count (
    .clk_i,
    .rst_ni,
    .clr_i(clr_sentmsg),
    .set_i(1'b0),
    .set_cnt_i(KeccakCountW'(0)),
    .incr_en_i(inc_sentmsg),
    .decr_en_i(1'b0),
    .step_i(KeccakCountW'(1)),
    .cnt_o(sent_message),
    .cnt_next_o(),
    .err_o(msg_count_error_o)
  );


  assign inc_sentmsg = keccak_valid_o & keccak_ready_i ;

  // Prefix index to slice the `prefix` n-bits into multiple of 64bit.
  logic [KeccakMsgAddrW-1:0] prefix_index;
  assign prefix_index = (sent_message < block_addr_limit) ? sent_message : '0;

  // fsm_keccak_valid is an output signal from FSM which to send data generated
  // inside the pad logic to keccak_round
  logic fsm_keccak_valid;

  // hold_msg to prevent message from being forwarded into keccak_round and
  // acked. Mainly the usage is to hold the message and initiates the
  // keccak_round for current block.
  logic hold_msg;

  // latch the partial write. Latched data is used for funcpad_merged
  logic en_msgbuf;
  logic clr_msgbuf;

  ///////////////////
  // State Machine //
  ///////////////////

  // Inputs

  // FSM moves to StPrefix only when cSHAKE is enabled
  logic mode_eq_cshake;
  assign mode_eq_cshake = (mode_i == CShake) ? 1'b 1 : 1'b 0;

  // `sent_blocksize` indicates the pad logic pushed block size data into
  // keccak round logic.
  logic sent_blocksize;

  assign sent_blocksize = (sent_message == block_addr_limit) ? 1'b 1 : 1'b 0;

  // `keccak_ack` indicates the request is accepted in keccak_round
  logic keccak_ack;

  assign keccak_ack = keccak_valid_o & keccak_ready_i ;

  // msg_partial indicates the incoming message is partial write or not.
  // This is used to check if the incoming message need to be latched inside or
  // not. If no partial message is at the end, msg_buf doesn't have to latch
  // msg_data_i. It is assumed that the partial message is permitted only at
  // the end of the message. So if (msg_valid_i && msg_partial && msg_ready_o),
  // there will be no msg_valid_i till process_latched.
  // Shall be used with msg_valid_i together.
  logic msg_partial;
  assign msg_partial = (&msg_strb_i != 1'b 1);


  // `process_latched` latches the `process_i` input before it is seen in the
  // FSM. `process_i` may follow `start_i` too fast so that the FSM may not
  // see it fast enought in case of cSHAKE mode. cSHAKE needs to process the
  // prefix prior to see the process indicator.
  logic process_latched;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      process_latched <= 1'b 0;
    end else if (process_i) begin
      process_latched <= 1'b 1;
    end else if (prim_mubi_pkg::mubi4_test_true_strict(done_i)) begin
      process_latched <= 1'b0;
    end
  end

  // State Register ===========================================================
  pad_st_e st, st_d;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, st_d, st, pad_st_e, StPadIdle)

  // `end_of_block` indicates current beat is end of the block
  // It shall set when the address reaches to the end of the block. End address
  // is set by the strength_i, which is `block_addr_limit`.
  logic end_of_block;

  assign end_of_block = ((sent_message + 1'b1) == block_addr_limit) ? 1'b 1 : 1'b 0;


  // Next logic and output logic ==============================================
  // SEC_CM: ABSORBED.CTRL.MUBI
  prim_mubi_pkg::mubi4_t absorbed_d;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) absorbed_o <= prim_mubi_pkg::MuBi4False;
    else         absorbed_o <= absorbed_d;
  end

  always_comb begin
    st_d = st;

    // FSM output : default values
    keccak_run_o = 1'b 0;
    sel_mux      = MuxNone;

    fsm_keccak_valid = 1'b 0;

    hold_msg = 1'b 0;
    clr_sentmsg = 1'b 0;

    en_msgbuf = 1'b 0;
    clr_msgbuf = 1'b 0;

    absorbed_d = prim_mubi_pkg::MuBi4False;

    sparse_fsm_error_o = 1'b 0;

    unique case (st)

      // In Idle state, the FSM checks if the software (or upper FSM) initiates
      // the hash process. If `start_i` is asserted (assume it is pulse), FSM
      // starts to push the data into the keccak round logic. Depending on the
      // hashing mode, FSM may push additional prefex in front of the actual
      // message. It means, the message could be back-pressured until the first
      // prefix is processed.
      StPadIdle: begin
        if (start_i) begin
          // If cSHAKE, move to Prefix state
          if (mode_eq_cshake) begin
            st_d = StPrefix;
          end else begin
            st_d = StMessage;
          end
        end else begin
          st_d = StPadIdle;
        end
      end

      // At Prefix state, FSM pushes
      // `bytepad(encode_string(N)||encode_string(S), 168or136)`. The software
      // already prepared `encode_string(N) || encode_string(S)` in the regs.
      // So, the FSM adds 2Byte in front of ns_data_i, which is an encoded
      // block size (see `encoded_bytepad` below)
      // After pushing the prefix, it initiates the hash process and move to
      // Message state.
      StPrefix: begin
        sel_mux = MuxPrefix;

        if (sent_blocksize) begin
          st_d = StPrefixWait;

          keccak_run_o = 1'b 1;
          fsm_keccak_valid = 1'b 0;
          clr_sentmsg = 1'b 1;
        end else begin
          st_d = StPrefix;

          fsm_keccak_valid = 1'b 1;
        end
      end

      StPrefixWait: begin
        sel_mux = MuxPrefix;

        if (keccak_complete_i) begin
          st_d = StMessage;
        end else begin
          st_d = StPrefixWait;
        end
      end

      // Message state pushes the incoming message into keccak round logic.
      // It forwards the message while counting the data and if it reaches
      // the block size, it triggers the keccak round to run. If `process` is
      // set, it moves to Pad state.
      StMessage: begin
        sel_mux = MuxFifo;

        if (msg_valid_i && msg_partial) begin
          st_d = StMessage;

          en_msgbuf = 1'b 1;
        end else if (sent_blocksize) begin
          // Check block completion first even process is set.
          st_d = StMessageWait;

          keccak_run_o = 1'b 1;
          clr_sentmsg = 1'b 1;
          hold_msg = 1'b 1;
        end else if (process_latched || process_i) begin
          st_d = StPad;

          // Not asserting the msg_ready_o
          hold_msg = 1'b 1;
        end else begin
          st_d = StMessage;

        end
      end

      StMessageWait: begin
        hold_msg = 1'b 1;

        if (keccak_complete_i) begin
          st_d = StMessage;
        end else begin
          st_d = StMessageWait;
        end
      end

      // Pad state just pushes the ending suffix. Depending on the mode, the
      // padding value is unique. SHA3 adds 2'b10, SHAKE adds 4'b1111, and
      // cSHAKE adds 2'b 00. Refer `function_pad`. The signal has one more bit
      // defined to accomodate first 1 bit of `pad10*1()` function.
      StPad: begin
        sel_mux = MuxFuncPad;

        fsm_keccak_valid = 1'b 1;

        if (keccak_ack && end_of_block) begin
          // If padding is the last block, don't have to move to StPad01, just
          // run Keccak and complete
          st_d = StPadRun;

          // always clear the latched msgbuf
          clr_msgbuf = 1'b 1;
          clr_sentmsg = 1'b 1;
        end else if (keccak_ack) begin
          st_d = StPad01;
          clr_msgbuf = 1'b 1;
        end else begin
          st_d = StPad;
        end
      end

      StPadRun: begin
        st_d = StPadFlush;

        keccak_run_o = 1'b 1;
        clr_sentmsg = 1'b 1;
      end

      // Pad01 pushes the end bit of pad10*1() function. As keccak accepts byte
      // size only, StPad always pushes partial (5bits). So at this state, it
      // pushes rest of 3bits. If the data pushed in StPad is the last byte of
      // the block, then Pad01 pushes to the same byte, if not, it first
      // zero-fill the block then pad 1 to the end.
      StPad01: begin
        sel_mux = MuxZeroEnd;

        // There's no chance StPad01 can be a start of the block. So can be
        // discard that the sent_blocksize is set at the beginning.
        if (sent_blocksize) begin
          st_d = StPadFlush;

          fsm_keccak_valid = 1'b 0;
          keccak_run_o = 1'b 1;
          clr_sentmsg = 1'b 1;
        end else begin
          st_d = StPad01;

          fsm_keccak_valid = 1'b 1;
        end
      end

      StPadFlush: begin
        // Wait completion from keccak_round or wait SW indicator.
        clr_sentmsg = 1'b 1;
        clr_msgbuf = 1'b 1;

        if (keccak_complete_i) begin
          st_d = StPadIdle;

          absorbed_d = prim_mubi_pkg::MuBi4True;
        end else begin
          st_d = StPadFlush;
        end
      end

      StTerminalError: begin
        // this state is terminal
        st_d = st;
        sparse_fsm_error_o = 1'b 1;
      end

      default: begin
        // this state is terminal
        st_d = StTerminalError;
        sparse_fsm_error_o = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      st_d = StTerminalError;
    end
  end

  //////////////
  // Datapath //
  //////////////

  // `encode_bytepad` represents the first two bytes of bytepad()
  // It depends on the block size. We can reuse KeccakRate
  // 10000000 || 00010101 // 168
  // 10000000 || 00010001 // 136
  logic [15:0] encode_bytepad;

  assign encode_bytepad = encode_bytepad_len(strength_i);

  // Prefix size ==============================================================
  // Prefix represents bytepad(encode_string(N) || encode_string(S), 168 or 136)
  // encode_string(N) || encode_string(S) is prepared by the software and given
  // through `ns_data_i`. The first part of bytepad is determined by the
  // `strength_i` and stored into `encode_bytepad`.

  // It is assumed that the prefix always smaller than the block size.
  logic [PrefixSize*8-1:0] prefix;

  assign prefix = {ns_data_i, encode_bytepad};

  logic [MsgWidth-1:0] prefix_sliced;
  logic [MsgWidth-1:0] prefix_data [Share];

  prim_slicer #(
    .InW (PrefixSize*8),
    .IndexW(KeccakMsgAddrW),
    .OutW(MsgWidth)
  ) u_prefix_slicer (
    .sel_i  (prefix_index),
    .data_i (prefix),
    .data_o (prefix_sliced)
  );

  if (EnMasking) begin : gen_prefix_masked
    // If Masking is enabled, prefix is two share.
    assign prefix_data[0] = '0;
    assign prefix_data[1] = prefix_sliced;
  end else begin : gen_prefix_unmasked
    // If Unmasked, only one share exists.
    assign prefix_data[0] = prefix_sliced;
  end

  // ==========================================================================
  // function_pad is the unique value padded at the end of the message based on
  // the function among SHA3, SHAKE, cSHAKE. The standard mentioned that SHA3
  // pads `01` , SHAKE pads `1111`, and cSHAKE pads `00`.
  //
  // Then pad10*1() function follows. It adds `1` first then fill 0 until it
  // reaches the block size -1, then adds `1`.
  //
  // It means always `1` is followed by the function pad.
  logic [4:0] funcpad;

  logic [MsgWidth-1:0] funcpad_data [Share];

  always_comb begin
    unique case (mode_i)
      Sha3:   funcpad = 5'b 00110;
      Shake:  funcpad = 5'b 11111;
      CShake: funcpad = 5'b 00100;

      default: begin
        // Just create non-padding but pad10*1 only
        funcpad = 5'b 00001;
      end
    endcase
  end

  // ==========================================================================
  // `zero_with_endbit` contains all zero unless the message is for the last
  // MsgWidth beat in the block. If it is the end of the block, the last bit
  // will be set to complete pad10*1() functionality.
  logic [MsgWidth-1:0] zero_with_endbit [Share];

  if (EnMasking) begin : gen_zeroend_masked
    assign zero_with_endbit[0]               = '0;
    assign zero_with_endbit[1][MsgWidth-1]   = end_of_block;
    assign zero_with_endbit[1][MsgWidth-2:0] = '0;
  end else begin : gen_zeroend_unmasked
    assign zero_with_endbit[0][MsgWidth-1]   = end_of_block;
    assign zero_with_endbit[0][MsgWidth-2:0] = '0;
  end

  // ==========================================================================
  // Data mux for output data

  assign keccak_addr_o = (sent_message < block_addr_limit) ? sent_message : '0;

  always_comb begin
    unique case (sel_mux)
      MuxFifo:    keccak_data_o = msg_data_i;
      MuxPrefix:  keccak_data_o = prefix_data;
      MuxFuncPad: keccak_data_o = funcpad_data;
      MuxZeroEnd: keccak_data_o = zero_with_endbit;

      // MuxNone
      default:  keccak_data_o = '{default:'0};
    endcase
  end

  always_comb begin
    unique case (sel_mux)
      MuxFifo:    keccak_valid_o = msg_valid_i & ~hold_msg & ~en_msgbuf;
      MuxPrefix:  keccak_valid_o = fsm_keccak_valid;
      MuxFuncPad: keccak_valid_o = fsm_keccak_valid;
      MuxZeroEnd: keccak_valid_o = fsm_keccak_valid;

      // MuxNone
      default:  keccak_valid_o = 1'b 0;
    endcase
  end

  always_comb begin
    unique case (sel_mux)
      MuxFifo:    msg_ready_o = en_msgbuf | (keccak_ready_i & ~hold_msg);
      MuxPrefix:  msg_ready_o = 1'b 0;
      MuxFuncPad: msg_ready_o = 1'b 0;
      MuxZeroEnd: msg_ready_o = 1'b 0;

      // MuxNone
      default: msg_ready_o = 1'b 0;
    endcase
  end

  // prim_packer : packing to 64bit to update keccak storage
  // two prim_packer in this module are used to pack the data received from
  // upper layer (KMAC core) and also the 5bit padding bits.
  // It is assumed that the message from upper layer could be partial at the
  // end of the message. Then the 2 or 4bit padding is required. It can be
  // handled by some custom logic or could be done by prim_packer.
  // If packer is used, the MSG_FIFO doesn't have to have another prim_packer
  // in front of the FIFO. This logic can handle the partial writes from the
  // software.
  //
  // If a custom logic is implemented here, prim_packer is necessary in front
  // of the FIFO, as this logic only appends at the end of the message when
  // `process_i` is asserted. Also, in this case, even prim_packer is not
  // needed, still 64bit registers to latch the partial write is required.
  // If not, the logic has to delay the acceptance of the incoming write
  // accesses. It may trigger the back-pressuring in some case which may result
  // that the software(or upper layer) may not set process_i.
  //
  // For custom logic, it could be implemented by the 8 mux selection.
  // for instance: (subject to be changed)
  //   unique case (sent_byte[2:0]) // generated from msg_strb_i
  //     3'b 000: funcpad_merged = {end_of_block, 63'(function_pad)                  };
  //     3'b 001: funcpad_merged = {end_of_block, 55'(function_pad), msg_data_i[ 7:0]};
  //     3'b 010: funcpad_merged = {end_of_block, 47'(function_pad), msg_data_i[15:0]};
  //     3'b 011: funcpad_merged = {end_of_block, 39'(function_pad), msg_data_i[23:0]};
  //     3'b 100: funcpad_merged = {end_of_block, 31'(function_pad), msg_data_i[31:0]};
  //     3'b 101: funcpad_merged = {end_of_block, 23'(function_pad), msg_data_i[39:0]};
  //     3'b 110: funcpad_merged = {end_of_block, 15'(function_pad), msg_data_i[47:0]};
  //     3'b 111: funcpad_merged = {end_of_block,  7'(function_pad), msg_data_i[55:0]};
  //     default: funcpad_merged = '0;
  //   endcase

  // internal buffer to store partial write. It doesn't have to store last byte as it
  // stores only when partial write.
  logic [MsgWidth-8-1:0] msg_buf [Share];
  logic [MsgStrbW-1-1:0] msg_strb;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      msg_buf  <= '{default:'0};
      msg_strb <= '0;
    end else if (en_msgbuf) begin
      for (int i = 0 ; i < Share ; i++) begin
        msg_buf[i]  <= msg_data_i[i][0+:(MsgWidth-8)];
      end
      msg_strb <= msg_strb_i[0+:(MsgStrbW-1)];
    end else if (clr_msgbuf) begin
      msg_buf  <= '{default:'0};
      msg_strb <= '0;
    end
  end

  if (EnMasking) begin : gen_funcpad_data_masked
    always_comb begin
      unique case (msg_strb)
        7'b 000_0000: begin
          funcpad_data[0] = '0;
          funcpad_data[1] = {end_of_block, 63'(funcpad)                  };
        end
        7'b 000_0001: begin
          funcpad_data[0] = {56'h0,                      msg_buf[0][ 7:0]};
          funcpad_data[1] = {end_of_block, 55'(funcpad), msg_buf[1][ 7:0]};
        end
        7'b 000_0011: begin
          funcpad_data[0] = {48'h0,                      msg_buf[0][15:0]};
          funcpad_data[1] = {end_of_block, 47'(funcpad), msg_buf[1][15:0]};
        end
        7'b 000_0111: begin
          funcpad_data[0] = {40'h0,                      msg_buf[0][23:0]};
          funcpad_data[1] = {end_of_block, 39'(funcpad), msg_buf[1][23:0]};
        end
        7'b 000_1111: begin
          funcpad_data[0] = {32'h0,                      msg_buf[0][31:0]};
          funcpad_data[1] = {end_of_block, 31'(funcpad), msg_buf[1][31:0]};
        end
        7'b 001_1111: begin
          funcpad_data[0] = {24'h0,                      msg_buf[0][39:0]};
          funcpad_data[1] = {end_of_block, 23'(funcpad), msg_buf[1][39:0]};
        end
        7'b 011_1111: begin
          funcpad_data[0] = {16'h0,                      msg_buf[0][47:0]};
          funcpad_data[1] = {end_of_block, 15'(funcpad), msg_buf[1][47:0]};
        end
        7'b 111_1111: begin
          funcpad_data[0] = { 8'h0,                      msg_buf[0][55:0]};
          funcpad_data[1] = {end_of_block,  7'(funcpad), msg_buf[1][55:0]};
        end

        default: funcpad_data = '{default:'0};
      endcase
    end
  end else begin : gen_funcpad_data_unmasked
    always_comb begin
      unique case (msg_strb)
        7'b 000_0000: funcpad_data[0] = {end_of_block, 63'(funcpad)                  };
        7'b 000_0001: funcpad_data[0] = {end_of_block, 55'(funcpad), msg_buf[0][ 7:0]};
        7'b 000_0011: funcpad_data[0] = {end_of_block, 47'(funcpad), msg_buf[0][15:0]};
        7'b 000_0111: funcpad_data[0] = {end_of_block, 39'(funcpad), msg_buf[0][23:0]};
        7'b 000_1111: funcpad_data[0] = {end_of_block, 31'(funcpad), msg_buf[0][31:0]};
        7'b 001_1111: funcpad_data[0] = {end_of_block, 23'(funcpad), msg_buf[0][39:0]};
        7'b 011_1111: funcpad_data[0] = {end_of_block, 15'(funcpad), msg_buf[0][47:0]};
        7'b 111_1111: funcpad_data[0] = {end_of_block,  7'(funcpad), msg_buf[0][55:0]};

        default: funcpad_data = '{default:'0};
      endcase
    end
  end

  ////////////////
  // Assertions //
  ////////////////

  // Prefix size is smaller than the smallest Keccak Block Size, which is 72 bytes.
  `ASSERT_INIT(PrefixLessThanBlock_A, PrefixSize/8 < KeccakRate[4])

  // Some part of datapath in sha3pad assumes Data width as 64bit.
  // If data width need to be changed, funcpad_data part should be changed too.
  // Also, The blocksize shall be divided by MsgWidth, which means, MsgWidth
  // can be {16, 32, 64} even funcpad_data mux is fully flexible.
  `ASSERT_INIT(MsgWidthidth_A, MsgWidth == 64)

  // Assume pulse signals: start, process, done
  `ASSUME(StartPulse_A, start_i |=> !start_i)
  `ASSUME(ProcessPulse_A, process_i |=> !process_i)
  `ASSUME(DonePulse_A,
    prim_mubi_pkg::mubi4_test_true_strict(done_i) |=>
      prim_mubi_pkg::mubi4_test_false_strict(done_i))

  // ASSERT output pulse signals: absorbed_o, keccak_run_o
  `ASSERT(AbsorbedPulse_A,
    prim_mubi_pkg::mubi4_test_true_strict(absorbed_o) |=>
      prim_mubi_pkg::mubi4_test_false_strict(absorbed_o))
  `ASSERT(KeccakRunPulse_A, keccak_run_o |=> !keccak_run_o)

  // start_i, done_i, process_i cannot set high at the same time
  `ASSUME(StartProcessDoneMutex_a,
    $onehot0({
      start_i,
      process_i,
      prim_mubi_pkg::mubi4_test_true_loose(done_i)
    }))

  // Sequence, start_i --> process_i --> absorbed_o --> done_i
  //`ASSUME(Sequence_a, start_i ##[1:$] process_i ##[1:$] ##[1:$] absorbed_o ##[1:$] done_i)

`ifndef SYNTHESIS
  // Process only asserts after start and all message are fed.
  // These valid signals are qualifier of FPV to trigger the control signal
  // It is a little bit hard to specify these criteria in SVA property so creating
  // qualifiers in RTL form is easier.
  logic start_valid, process_valid, absorb_valid, done_valid;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      start_valid <= 1'b 1;
    end else if (start_i) begin
      start_valid <= 1'b 0;
    end else if (prim_mubi_pkg::mubi4_test_true_strict(done_i)) begin
      start_valid <= 1'b 1;
    end
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      process_valid <= 1'b 0;
    end else if (start_i) begin
      process_valid <= 1'b 1;
    end else if (process_i) begin
      process_valid <= 1'b 0;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      done_valid <= 1'b 0;
    end else if (prim_mubi_pkg::mubi4_test_true_strict(absorbed_o)) begin
      done_valid <= 1'b 1;
    end else if (prim_mubi_pkg::mubi4_test_true_strict(done_i)) begin
      done_valid <= 1'b 0;
    end
  end

  // Message can be fed in between start_i and process_i.
  `ASSUME(MessageCondition_M, msg_valid_i && msg_ready_o |-> process_valid && !process_i)

  // Message ready should be asserted only in between start_i and process_i
  `ASSERT(MsgReadyCondition_A, msg_ready_o |-> process_valid && !process_i)

  `ASSUME(ProcessCondition_M, process_i |-> process_valid)
  `ASSUME(StartCondition_M, start_i |-> start_valid)
  `ASSUME(DoneCondition_M,
    prim_mubi_pkg::mubi4_test_true_strict(done_i) |-> done_valid)

  // Assume mode_i and strength_i are stable during the operation
  // This will be guarded at the kmac top level
  `ASSUME(ModeStableDuringOp_M,
    $changed(mode_i) |-> start_valid)
  `ASSUME(StrengthStableDuringOp_M,
    $changed(strength_i) |-> start_valid)

`endif // SYNTHESIS

  // If not full block is written, the pad shall send message to keccak_round
  // If it is end of the message, the state moves to StPad and send the request
  `ASSERT(CompleteBlockWhenProcess_A,
    $rose(process_latched) && (!end_of_block && !sent_blocksize )
    && !(st inside {StPrefixWait, StMessageWait}) |-> ##[1:5] keccak_valid_o,
    clk_i, !rst_ni || lc_escalate_en_i != lc_ctrl_pkg::Off)

  // If process_i asserted, completion shall be asserted shall be asserted
  //`ASSERT(ProcessToAbsorbed_A, process_i |=> strong(##[24*Share:$] absorbed_o))


  // Assumption of input mode_i and strength_i
  // SHA3 variants: SHA3-224, SHA3-256, SHA3-384, SHA3-512
  // SHAKE, cSHAKE variants: SHAKE128, SHAKE256, cSHAKE128, cSHAKE256
  `ASSUME_FPV(ModeStrengthCombinations_M,
    start_i |->
      (mode_i == Sha3 && (strength_i inside {L224, L256, L384, L512})) ||
      ((mode_i == Shake || mode_i == CShake) && (strength_i inside {L128, L256})),
    clk_i, !rst_ni)

  // No partial write is allowed for Message FIFO interface
  `ASSUME(NoPartialMsgFifo_M,
    keccak_valid_o && (sel_mux == MuxFifo) |-> (&msg_strb_i) == 1'b1,
    clk_i, !rst_ni)

  // When transaction is stored into msg_buf, it shall be partial write.
  `ASSUME(AlwaysPartialMsgBuf_M,
    en_msgbuf |-> msg_valid_i && (msg_strb_i[MsgStrbW-1] == 1'b0),
    clk_i, !rst_ni)

  // if partial write comes and is acked, then no more msg_valid_i until
  // next message
  `ASSUME(PartialEndOfMsg_M,
    msg_valid_i && msg_ready_o && msg_partial |=>
      !msg_valid_i ##[1:$] $stable(msg_valid_i) ##1 process_latched,
    clk_i, !rst_ni)

  // At the first clock in StPad01 state, sent_blocksize shall not be set
  `ASSERT(Pad01NotAttheEndOfBlock_A,
    (st == StPad && st_d == StPad01) |-> !end_of_block,
    clk_i, !rst_ni)

  // When data sent to the keccak_round, the address should be in the range
  `ASSERT(KeccakAddrInRange_A,
    keccak_valid_o |-> keccak_addr_o < KeccakRate[strength_i],
    clk_i, !rst_ni)

  // NS data shall be stable during the operation.
  //`ASSUME(NsStableInProcess_A,
  //  $stable(ns_data_i) throughout(start_i ##[1:$] process_i ##[1:$] absorbed_o),
  //  clk_i, !rst_ni)

  // Functional Coverage
  `COVER(StMessageFeed_C, st == StMessage)
  `COVER(StPad_C, st == StPad01 && sent_blocksize)
  `COVER(StPadSendMsg_C, st == StPad01 && keccak_ack)
  `COVER(StComplete_C, st == StPadFlush)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// SHA3 core is a fully functional SHA3/SHAKE/cSHAKE hashing module.
//
// It instantiates a keccak_round with 1600 bits of the state.

`include "prim_assert.sv"

module sha3
  import sha3_pkg::*;
#(
  // Enable Masked Keccak if 1
  parameter  bit EnMasking = 0,
  // derived parameter
  localparam int Share = (EnMasking) ? 2 : 1
) (
  input clk_i,
  input rst_ni,

  // MSG interface
  input                       msg_valid_i,
  input        [MsgWidth-1:0] msg_data_i [Share],
  input        [MsgStrbW-1:0] msg_strb_i,         // one strobe for shares
  output logic                msg_ready_o,

  // Entropy interface
  input                     rand_valid_i,
  input                     rand_early_i,
  input      [StateW/2-1:0] rand_data_i,
  input                     rand_aux_i,
  output logic              rand_consumed_o,

  // N, S: Used in cSHAKE mode only
  input [NSRegisterSize*8-1:0] ns_data_i, // See sha3_pkg for details

  // configurations
  input sha3_mode_e       mode_i,     // see sha3pad for details
  input keccak_strength_e strength_i, // see sha3pad for details

  // controls
  input start_i,   // see sha3pad for details
  input process_i, // see sha3pad for details

  // run_i is a pulse signal to trigger the keccak_round manually by SW.
  // It is used to run additional keccak_f after sponge absorbing is completed.
  // See `keccak_run` signal
  input                        run_i,
  input prim_mubi_pkg::mubi4_t done_i,    // see sha3pad for details

  output prim_mubi_pkg::mubi4_t absorbed_o,
  output logic                  squeezing_o,

  // Indicate of one block processed. KMAC main state tracks the progression
  // based on this signal.
  output logic block_processed_o,

  output sha3_st_e sha3_fsm_o,

  // digest output
  // This value is valid only after all absorbing process is completed.
  // In invalid state, the output `state` will be zero to prevent information
  // leakage.
  output logic              state_valid_o,
  output logic [StateW-1:0] state_o [Share],

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  // error_o value is pushed to Error FIFO at KMAC/SHA3 top and reported to SW
  output err_t error_o,

  // sparse_fsm_alert
  output logic sparse_fsm_error_o,

  // counter error
  output logic count_error_o,

  // error on rst_storage in Keccak
  output logic keccak_storage_rst_error_o

);
  /////////////////
  // Definitions //
  /////////////////

  typedef enum logic[2:0] {
    MuxGuard   = 3'b 010,
    MuxRelease = 3'b 101
  } state_mux_sel_e;

  /////////////
  // Signals //
  /////////////

  // State --> Digest
  // State is exposed to the outside if the hashing process is completed.
  logic              state_valid;
  logic [StateW-1:0] state [Share];
  logic [StateW-1:0] state_guarded [Share];

  // State --> digest mux select signal
  state_mux_sel_e mux_sel;

  // absorbed is a pulse signal that indicates sponge absorbing is done.
  // After this, sha3 core allows software to manually run until squeezing
  // is completed, which is the `done_i` pulse signal.
  prim_mubi_pkg::mubi4_t absorbed;

  // `squeezing` is a status indicator that SHA3 core is in sponge squeezing
  // stage. In this stage, the state output is valid, and software can manually
  // trigger keccak_round logic to get more digest outputs in case the output
  // length is bigger than the block limit.
  logic squeezing;

  // If process_i is received, the logic initiates the final absorbing process.
  // While absorbing, the processing inticator is turned on. This signal is used
  // to check if multiple process_i is received or not.
  logic processing;

  // FSM variable
  sha3_st_sparse_e st, st_d;

  // Keccak control signal (filtered by State Machine)
  logic keccak_start, keccak_process;
  prim_mubi_pkg::mubi4_t keccak_done;

  // alert signals
  logic round_count_error, msg_count_error;
  assign count_error_o =  round_count_error | msg_count_error;

  logic sha3_state_error;
  logic keccak_round_state_error;
  logic sha3pad_state_error;

  assign sparse_fsm_error_o = sha3_state_error | keccak_round_state_error | sha3pad_state_error;

  // Keccak rst_storage is asserted unexpectedly
  logic keccak_storage_rst_error;
  assign keccak_storage_rst_error_o = keccak_storage_rst_error;

  /////////////////
  // Connections //
  /////////////////

  logic                       keccak_valid;
  logic [KeccakMsgAddrW-1:0]  keccak_addr;
  logic [MsgWidth-1:0]        keccak_data [Share];
  logic                       keccak_ready;

  // Keccak round run signal can be controlled by sha3pad and also by software
  // after all message feeding is done. it is mainly used for sponge squeezing
  // operation after absorbing is completed when output length is longer than
  // the block size.
  logic keccak_run, sha3pad_keccak_run, sw_keccak_run;
  logic keccak_complete;

  assign keccak_run = sha3pad_keccak_run | sw_keccak_run;

  // Absorb pulse output : used to generate interrupts
  // Latch absorbed signal as kmac_keymgr asserts `CmdDone` when it sees
  // `absorbed` signal. When this signal goes out, the state is still in
  // `StAbsorb`. Next state is `StSqueeze`.
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) absorbed_o <= prim_mubi_pkg::MuBi4False;
    else         absorbed_o <= absorbed;
  end

  // Squeezing output
  assign squeezing_o = squeezing;

  // processing
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)        processing <= 1'b 0;
    else if (process_i) processing <= 1'b 1;
    else if (prim_mubi_pkg::mubi4_test_true_strict(absorbed)) begin
      processing <= 1'b 0;
    end
  end

  assign block_processed_o = keccak_complete;

  // State connection
  assign state_valid_o = state_valid;
  assign state_o = state_guarded;

  assign sha3_fsm_o = sparse2logic(st);

  ///////////////////
  // State Machine //
  ///////////////////

  // State Register
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, st_d, st, sha3_st_sparse_e, StIdle_sparse)


  // Next State and Output Logic
  // Mainly the FSM controls the input signal access
  // StIdle:    only start_i signal is allowed
  // StAbsorb:  only process_i signal is allowed
  // StSqueeze: only run_i, done_i signal is allowed

  always_comb begin
    st_d = st;

    // default output values
    keccak_start = 1'b 0;
    keccak_process = 1'b 0;
    sw_keccak_run = 1'b 0;
    keccak_done = prim_mubi_pkg::MuBi4False;

    squeezing = 1'b 0;

    state_valid = 1'b 0;
    mux_sel = MuxGuard ;

    sha3_state_error = 1'b 0;

    unique case (st)
      StIdle_sparse: begin
        if (start_i) begin
          st_d = StAbsorb_sparse;

          keccak_start = 1'b 1;
        end else begin
          st_d = StIdle_sparse;
        end
      end

      StAbsorb_sparse: begin
        if (process_i && !processing) begin
          st_d = StAbsorb_sparse;

          keccak_process = 1'b 1;
        end else if (prim_mubi_pkg::mubi4_test_true_strict(absorbed)) begin
          st_d = StSqueeze_sparse;
        end else begin
          st_d = StAbsorb_sparse;
        end
      end

      StSqueeze_sparse: begin
        state_valid = 1'b 1;
        mux_sel = MuxRelease; // Expose state to register interface

        squeezing = 1'b 1;

        if (run_i) begin
          st_d = StManualRun_sparse;

          sw_keccak_run = 1'b 1;
        end else if (prim_mubi_pkg::mubi4_test_true_strict(done_i)) begin
          st_d = StFlush_sparse;

          keccak_done = done_i;
        end else begin
          st_d = StSqueeze_sparse;
        end
      end

      StManualRun_sparse: begin
        if (keccak_complete) begin
          st_d = StSqueeze_sparse;
        end else begin
          st_d = StManualRun_sparse;
        end
      end

      StFlush_sparse: begin
        st_d = StIdle_sparse;
      end

      StTerminalError_sparse: begin
        //this state is terminal
        st_d = StTerminalError_sparse;
        sha3_state_error = 1'b 1;
      end

      default: begin
        st_d = StTerminalError_sparse;
        sha3_state_error = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      st_d = StTerminalError_sparse;
    end
  end

  //////////////
  // Datapath //
  //////////////

  // State --> Digest output
  always_comb begin : state_guarded_mux
    unique case (mux_sel)
      MuxGuard:   state_guarded = '{default: '0};
      MuxRelease: state_guarded = state;
      default:    state_guarded = '{default: '0}; // a valid, safe output
    endcase
  end


  // Error Detecting
  // ErrSha3SwControl:
  //   info[ 0]: start_i set
  //   info[ 1]: process_i set
  //   info[ 2]: run_i set
  //   info[ 3]: done_i set
  //  - Sw set process_i, run_i, done_i without start_i

  always_comb begin
    error_o = '{valid: 1'b0, code: ErrNone, info: '0};

    unique case (st)
      StIdle_sparse: begin
        if (process_i || run_i ||
          prim_mubi_pkg::mubi4_test_true_loose(done_i)) begin
          error_o = '{
            valid: 1'b 1,
            code: ErrSha3SwControl,
            info: 24'({done_i, run_i, process_i, start_i})
          };
        end
      end

      StAbsorb_sparse: begin
        if (start_i || run_i || prim_mubi_pkg::mubi4_test_true_loose(done_i)
          || (process_i && processing)) begin
          error_o = '{
            valid: 1'b 1,
            code: ErrSha3SwControl,
            info: 24'({done_i, run_i, process_i, start_i})
          };
        end
      end

      StSqueeze_sparse: begin
        if (start_i || process_i) begin
          error_o = '{
            valid: 1'b 1,
            code: ErrSha3SwControl,
            info: 24'({done_i, run_i, process_i, start_i})
          };
        end
      end

      StManualRun_sparse: begin
        if (start_i || process_i || run_i ||
          prim_mubi_pkg::mubi4_test_true_loose(done_i)) begin
          error_o = '{
            valid: 1'b 1,
            code: ErrSha3SwControl,
            info: 24'({done_i, run_i, process_i, start_i})
          };
        end
      end

      StFlush_sparse: begin
        if (start_i || process_i || run_i ||
          prim_mubi_pkg::mubi4_test_true_loose(done_i)) begin
          error_o = '{
            valid: 1'b 1,
            code: ErrSha3SwControl,
            info: 24'({done_i, run_i, process_i, start_i})
          };
        end
      end

      default: begin
      end
    endcase
  end
  ///////////////
  // Instances //
  ///////////////

  // SHA3 pad logic
  sha3pad #(
    .EnMasking (EnMasking)
  ) u_pad (
    .clk_i,
    .rst_ni,

    // MSG_FIFO (or from KMAC core)
    .msg_valid_i,
    .msg_data_i, // [Share]
    .msg_strb_i,
    .msg_ready_o,

    // Encoded N, S
    .ns_data_i,

    // output to keccak_round: message path
    .keccak_valid_o (keccak_valid),
    .keccak_addr_o  (keccak_addr ),
    .keccak_data_o  (keccak_data ), // [Share]
    .keccak_ready_i (keccak_ready),

    .keccak_run_o      (sha3pad_keccak_run),
    .keccak_complete_i (keccak_complete   ),

    // configurations
    .mode_i,
    .strength_i,

    // LC
    .lc_escalate_en_i (lc_escalate_en_i),

    // controls
    .start_i   (keccak_start),
    .process_i (keccak_process),
    .done_i    (keccak_done),

    // output
    .absorbed_o         (absorbed),
    .sparse_fsm_error_o (sha3pad_state_error),
    .msg_count_error_o  (msg_count_error)
  );

  // Keccak round logic
  keccak_round #(
    .Width    (sha3_pkg::StateW),
    .DInWidth (sha3_pkg::MsgWidth),

    .EnMasking  (EnMasking)
  ) u_keccak (
    .clk_i,
    .rst_ni,

    .valid_i (keccak_valid),
    .addr_i  (keccak_addr ),
    .data_i  (keccak_data ),
    .ready_o (keccak_ready),

    .rand_valid_i,
    .rand_early_i,
    .rand_data_i,
    .rand_aux_i,
    .rand_consumed_o,

    .run_i      (keccak_run     ),
    .complete_o (keccak_complete),

    .state_o    (state),

    // LC
    .lc_escalate_en_i (lc_escalate_en_i),

    .sparse_fsm_error_o  (keccak_round_state_error),
    .round_count_error_o (round_count_error),
    .rst_storage_error_o (keccak_storage_rst_error),

    .clear_i    (keccak_done)
  );

  ////////////////
  // Assertions //
  ////////////////

  // Unknown check for case statement
  `ASSERT(MuxSelKnown_A, mux_sel inside {MuxGuard, MuxRelease})
  `ASSERT(FsmKnown_A, st inside {StIdle_sparse, StAbsorb_sparse, StSqueeze_sparse,
                                 StManualRun_sparse, StFlush_sparse, StTerminalError_sparse})

  // `state` shall be 0 in invalid
  if (EnMasking) begin: gen_chk_digest_masked
    `ASSERT(StateZeroInvalid_A, !state_valid_o |-> ((|state_o[0]) | (|state_o[1])) == 1'b 0)
  end else begin : gen_chk_digest_unmasked
    `ASSERT(StateZeroInvalid_A, !state_valid_o |-> (|state_o[0]) == 1'b 0)
  end

  // `state_valid_o` asserts only in between the completion and done
  //`ASSERT(StateValidPeriod_A, state_valid_o |-> )

  // skip the msg interface assertions as they are in sha3pad.sv

  // Software run signal happens in Squeezing stage
  `ASSUME(SwRunInSqueezing_a, run_i |-> error_o.valid || (st == StSqueeze_sparse))

  // If control received but not propagated into submodules, it is error condition
  `ASSERT(ErrDetection_A, error_o.valid
    |-> {start_i,      process_i,      run_i,         done_i}
     != {keccak_start, keccak_process, sw_keccak_run, keccak_done})

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module csrng_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output csrng_reg_pkg::csrng_reg2hw_t reg2hw, // Write
  input  csrng_reg_pkg::csrng_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import csrng_reg_pkg::* ;

  localparam int AW = 7;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [16:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(17)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_cs_cmd_req_done_qs;
  logic intr_state_cs_cmd_req_done_wd;
  logic intr_state_cs_entropy_req_qs;
  logic intr_state_cs_entropy_req_wd;
  logic intr_state_cs_hw_inst_exc_qs;
  logic intr_state_cs_hw_inst_exc_wd;
  logic intr_state_cs_fatal_err_qs;
  logic intr_state_cs_fatal_err_wd;
  logic intr_enable_we;
  logic intr_enable_cs_cmd_req_done_qs;
  logic intr_enable_cs_cmd_req_done_wd;
  logic intr_enable_cs_entropy_req_qs;
  logic intr_enable_cs_entropy_req_wd;
  logic intr_enable_cs_hw_inst_exc_qs;
  logic intr_enable_cs_hw_inst_exc_wd;
  logic intr_enable_cs_fatal_err_qs;
  logic intr_enable_cs_fatal_err_wd;
  logic intr_test_we;
  logic intr_test_cs_cmd_req_done_wd;
  logic intr_test_cs_entropy_req_wd;
  logic intr_test_cs_hw_inst_exc_wd;
  logic intr_test_cs_fatal_err_wd;
  logic alert_test_we;
  logic alert_test_recov_alert_wd;
  logic alert_test_fatal_alert_wd;
  logic regwen_we;
  logic regwen_qs;
  logic regwen_wd;
  logic ctrl_we;
  logic [3:0] ctrl_enable_qs;
  logic [3:0] ctrl_enable_wd;
  logic [3:0] ctrl_sw_app_enable_qs;
  logic [3:0] ctrl_sw_app_enable_wd;
  logic [3:0] ctrl_read_int_state_qs;
  logic [3:0] ctrl_read_int_state_wd;
  logic cmd_req_we;
  logic [31:0] cmd_req_wd;
  logic sw_cmd_sts_cmd_rdy_qs;
  logic sw_cmd_sts_cmd_sts_qs;
  logic genbits_vld_re;
  logic genbits_vld_genbits_vld_qs;
  logic genbits_vld_genbits_fips_qs;
  logic genbits_re;
  logic [31:0] genbits_qs;
  logic int_state_num_we;
  logic [3:0] int_state_num_qs;
  logic [3:0] int_state_num_wd;
  logic int_state_val_re;
  logic [31:0] int_state_val_qs;
  logic hw_exc_sts_we;
  logic [15:0] hw_exc_sts_qs;
  logic [15:0] hw_exc_sts_wd;
  logic recov_alert_sts_we;
  logic recov_alert_sts_enable_field_alert_qs;
  logic recov_alert_sts_enable_field_alert_wd;
  logic recov_alert_sts_sw_app_enable_field_alert_qs;
  logic recov_alert_sts_sw_app_enable_field_alert_wd;
  logic recov_alert_sts_read_int_state_field_alert_qs;
  logic recov_alert_sts_read_int_state_field_alert_wd;
  logic recov_alert_sts_acmd_flag0_field_alert_qs;
  logic recov_alert_sts_acmd_flag0_field_alert_wd;
  logic recov_alert_sts_cs_bus_cmp_alert_qs;
  logic recov_alert_sts_cs_bus_cmp_alert_wd;
  logic recov_alert_sts_cs_main_sm_alert_qs;
  logic recov_alert_sts_cs_main_sm_alert_wd;
  logic err_code_sfifo_cmd_err_qs;
  logic err_code_sfifo_genbits_err_qs;
  logic err_code_sfifo_cmdreq_err_qs;
  logic err_code_sfifo_rcstage_err_qs;
  logic err_code_sfifo_keyvrc_err_qs;
  logic err_code_sfifo_updreq_err_qs;
  logic err_code_sfifo_bencreq_err_qs;
  logic err_code_sfifo_bencack_err_qs;
  logic err_code_sfifo_pdata_err_qs;
  logic err_code_sfifo_final_err_qs;
  logic err_code_sfifo_gbencack_err_qs;
  logic err_code_sfifo_grcstage_err_qs;
  logic err_code_sfifo_ggenreq_err_qs;
  logic err_code_sfifo_gadstage_err_qs;
  logic err_code_sfifo_ggenbits_err_qs;
  logic err_code_sfifo_blkenc_err_qs;
  logic err_code_cmd_stage_sm_err_qs;
  logic err_code_main_sm_err_qs;
  logic err_code_drbg_gen_sm_err_qs;
  logic err_code_drbg_updbe_sm_err_qs;
  logic err_code_drbg_updob_sm_err_qs;
  logic err_code_aes_cipher_sm_err_qs;
  logic err_code_cmd_gen_cnt_err_qs;
  logic err_code_fifo_write_err_qs;
  logic err_code_fifo_read_err_qs;
  logic err_code_fifo_state_err_qs;
  logic err_code_test_we;
  logic [4:0] err_code_test_qs;
  logic [4:0] err_code_test_wd;
  logic [7:0] main_sm_state_qs;

  // Register instances
  // R[intr_state]: V(False)
  //   F[cs_cmd_req_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_cs_cmd_req_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_cs_cmd_req_done_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.cs_cmd_req_done.de),
    .d      (hw2reg.intr_state.cs_cmd_req_done.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.cs_cmd_req_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_cs_cmd_req_done_qs)
  );

  //   F[cs_entropy_req]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_cs_entropy_req (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_cs_entropy_req_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.cs_entropy_req.de),
    .d      (hw2reg.intr_state.cs_entropy_req.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.cs_entropy_req.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_cs_entropy_req_qs)
  );

  //   F[cs_hw_inst_exc]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_cs_hw_inst_exc (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_cs_hw_inst_exc_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.cs_hw_inst_exc.de),
    .d      (hw2reg.intr_state.cs_hw_inst_exc.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.cs_hw_inst_exc.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_cs_hw_inst_exc_qs)
  );

  //   F[cs_fatal_err]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_cs_fatal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_cs_fatal_err_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.cs_fatal_err.de),
    .d      (hw2reg.intr_state.cs_fatal_err.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.cs_fatal_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_cs_fatal_err_qs)
  );


  // R[intr_enable]: V(False)
  //   F[cs_cmd_req_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_cs_cmd_req_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_cs_cmd_req_done_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.cs_cmd_req_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_cs_cmd_req_done_qs)
  );

  //   F[cs_entropy_req]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_cs_entropy_req (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_cs_entropy_req_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.cs_entropy_req.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_cs_entropy_req_qs)
  );

  //   F[cs_hw_inst_exc]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_cs_hw_inst_exc (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_cs_hw_inst_exc_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.cs_hw_inst_exc.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_cs_hw_inst_exc_qs)
  );

  //   F[cs_fatal_err]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_cs_fatal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_cs_fatal_err_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.cs_fatal_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_cs_fatal_err_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [3:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  //   F[cs_cmd_req_done]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_cs_cmd_req_done (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_cs_cmd_req_done_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.cs_cmd_req_done.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.cs_cmd_req_done.qe = intr_test_qe;

  //   F[cs_entropy_req]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_cs_entropy_req (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_cs_entropy_req_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[1]),
    .q      (reg2hw.intr_test.cs_entropy_req.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.cs_entropy_req.qe = intr_test_qe;

  //   F[cs_hw_inst_exc]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_cs_hw_inst_exc (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_cs_hw_inst_exc_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[2]),
    .q      (reg2hw.intr_test.cs_hw_inst_exc.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.cs_hw_inst_exc.qe = intr_test_qe;

  //   F[cs_fatal_err]: 3:3
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_cs_fatal_err (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_cs_fatal_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[3]),
    .q      (reg2hw.intr_test.cs_fatal_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.cs_fatal_err.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[recov_alert]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov_alert (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_alert_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.recov_alert.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov_alert.qe = alert_test_qe;

  //   F[fatal_alert]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal_alert (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_alert_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.fatal_alert.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal_alert.qe = alert_test_qe;


  // R[regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (regwen_we),
    .wd     (regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (regwen_qs)
  );


  // R[ctrl]: V(False)
  // Create REGWEN-gated WE signal
  logic ctrl_gated_we;
  assign ctrl_gated_we = ctrl_we & regwen_qs;
  //   F[enable]: 3:0
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_enable_qs)
  );

  //   F[sw_app_enable]: 7:4
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_sw_app_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_sw_app_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.sw_app_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_sw_app_enable_qs)
  );

  //   F[read_int_state]: 11:8
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_ctrl_read_int_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_gated_we),
    .wd     (ctrl_read_int_state_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.read_int_state.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_read_int_state_qs)
  );


  // R[cmd_req]: V(False)
  logic cmd_req_qe;
  logic [0:0] cmd_req_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_cmd_req0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&cmd_req_flds_we),
    .q_o(cmd_req_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (32'h0)
  ) u_cmd_req (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (cmd_req_we),
    .wd     (cmd_req_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cmd_req_flds_we[0]),
    .q      (reg2hw.cmd_req.q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );
  assign reg2hw.cmd_req.qe = cmd_req_qe;


  // R[sw_cmd_sts]: V(False)
  //   F[cmd_rdy]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h1)
  ) u_sw_cmd_sts_cmd_rdy (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.sw_cmd_sts.cmd_rdy.de),
    .d      (hw2reg.sw_cmd_sts.cmd_rdy.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_cmd_sts_cmd_rdy_qs)
  );

  //   F[cmd_sts]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_sw_cmd_sts_cmd_sts (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.sw_cmd_sts.cmd_sts.de),
    .d      (hw2reg.sw_cmd_sts.cmd_sts.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_cmd_sts_cmd_sts_qs)
  );


  // R[genbits_vld]: V(True)
  //   F[genbits_vld]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_genbits_vld_genbits_vld (
    .re     (genbits_vld_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.genbits_vld.genbits_vld.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (genbits_vld_genbits_vld_qs)
  );

  //   F[genbits_fips]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_genbits_vld_genbits_fips (
    .re     (genbits_vld_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.genbits_vld.genbits_fips.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (genbits_vld_genbits_fips_qs)
  );


  // R[genbits]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_genbits (
    .re     (genbits_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.genbits.d),
    .qre    (reg2hw.genbits.re),
    .qe     (),
    .q      (reg2hw.genbits.q),
    .ds     (),
    .qs     (genbits_qs)
  );


  // R[int_state_num]: V(False)
  logic int_state_num_qe;
  logic [0:0] int_state_num_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_int_state_num0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&int_state_num_flds_we),
    .q_o(int_state_num_qe)
  );
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h0)
  ) u_int_state_num (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (int_state_num_we),
    .wd     (int_state_num_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (int_state_num_flds_we[0]),
    .q      (reg2hw.int_state_num.q),
    .ds     (),

    // to register interface (read)
    .qs     (int_state_num_qs)
  );
  assign reg2hw.int_state_num.qe = int_state_num_qe;


  // R[int_state_val]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_int_state_val (
    .re     (int_state_val_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.int_state_val.d),
    .qre    (reg2hw.int_state_val.re),
    .qe     (),
    .q      (reg2hw.int_state_val.q),
    .ds     (),
    .qs     (int_state_val_qs)
  );


  // R[hw_exc_sts]: V(False)
  prim_subreg #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (16'h0)
  ) u_hw_exc_sts (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (hw_exc_sts_we),
    .wd     (hw_exc_sts_wd),

    // from internal hardware
    .de     (hw2reg.hw_exc_sts.de),
    .d      (hw2reg.hw_exc_sts.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (hw_exc_sts_qs)
  );


  // R[recov_alert_sts]: V(False)
  //   F[enable_field_alert]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_enable_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_enable_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.enable_field_alert.de),
    .d      (hw2reg.recov_alert_sts.enable_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_enable_field_alert_qs)
  );

  //   F[sw_app_enable_field_alert]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_sw_app_enable_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_sw_app_enable_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.sw_app_enable_field_alert.de),
    .d      (hw2reg.recov_alert_sts.sw_app_enable_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_sw_app_enable_field_alert_qs)
  );

  //   F[read_int_state_field_alert]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_read_int_state_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_read_int_state_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.read_int_state_field_alert.de),
    .d      (hw2reg.recov_alert_sts.read_int_state_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_read_int_state_field_alert_qs)
  );

  //   F[acmd_flag0_field_alert]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_acmd_flag0_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_acmd_flag0_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.acmd_flag0_field_alert.de),
    .d      (hw2reg.recov_alert_sts.acmd_flag0_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_acmd_flag0_field_alert_qs)
  );

  //   F[cs_bus_cmp_alert]: 12:12
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_cs_bus_cmp_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_cs_bus_cmp_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.cs_bus_cmp_alert.de),
    .d      (hw2reg.recov_alert_sts.cs_bus_cmp_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_cs_bus_cmp_alert_qs)
  );

  //   F[cs_main_sm_alert]: 13:13
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_cs_main_sm_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_cs_main_sm_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.cs_main_sm_alert.de),
    .d      (hw2reg.recov_alert_sts.cs_main_sm_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_cs_main_sm_alert_qs)
  );


  // R[err_code]: V(False)
  //   F[sfifo_cmd_err]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_cmd_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_cmd_err.de),
    .d      (hw2reg.err_code.sfifo_cmd_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_cmd_err_qs)
  );

  //   F[sfifo_genbits_err]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_genbits_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_genbits_err.de),
    .d      (hw2reg.err_code.sfifo_genbits_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_genbits_err_qs)
  );

  //   F[sfifo_cmdreq_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_cmdreq_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_cmdreq_err.de),
    .d      (hw2reg.err_code.sfifo_cmdreq_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_cmdreq_err_qs)
  );

  //   F[sfifo_rcstage_err]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_rcstage_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_rcstage_err.de),
    .d      (hw2reg.err_code.sfifo_rcstage_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_rcstage_err_qs)
  );

  //   F[sfifo_keyvrc_err]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_keyvrc_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_keyvrc_err.de),
    .d      (hw2reg.err_code.sfifo_keyvrc_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_keyvrc_err_qs)
  );

  //   F[sfifo_updreq_err]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_updreq_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_updreq_err.de),
    .d      (hw2reg.err_code.sfifo_updreq_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_updreq_err_qs)
  );

  //   F[sfifo_bencreq_err]: 6:6
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_bencreq_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_bencreq_err.de),
    .d      (hw2reg.err_code.sfifo_bencreq_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_bencreq_err_qs)
  );

  //   F[sfifo_bencack_err]: 7:7
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_bencack_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_bencack_err.de),
    .d      (hw2reg.err_code.sfifo_bencack_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_bencack_err_qs)
  );

  //   F[sfifo_pdata_err]: 8:8
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_pdata_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_pdata_err.de),
    .d      (hw2reg.err_code.sfifo_pdata_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_pdata_err_qs)
  );

  //   F[sfifo_final_err]: 9:9
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_final_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_final_err.de),
    .d      (hw2reg.err_code.sfifo_final_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_final_err_qs)
  );

  //   F[sfifo_gbencack_err]: 10:10
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_gbencack_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_gbencack_err.de),
    .d      (hw2reg.err_code.sfifo_gbencack_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_gbencack_err_qs)
  );

  //   F[sfifo_grcstage_err]: 11:11
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_grcstage_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_grcstage_err.de),
    .d      (hw2reg.err_code.sfifo_grcstage_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_grcstage_err_qs)
  );

  //   F[sfifo_ggenreq_err]: 12:12
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_ggenreq_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_ggenreq_err.de),
    .d      (hw2reg.err_code.sfifo_ggenreq_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_ggenreq_err_qs)
  );

  //   F[sfifo_gadstage_err]: 13:13
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_gadstage_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_gadstage_err.de),
    .d      (hw2reg.err_code.sfifo_gadstage_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_gadstage_err_qs)
  );

  //   F[sfifo_ggenbits_err]: 14:14
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_ggenbits_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_ggenbits_err.de),
    .d      (hw2reg.err_code.sfifo_ggenbits_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_ggenbits_err_qs)
  );

  //   F[sfifo_blkenc_err]: 15:15
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_blkenc_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_blkenc_err.de),
    .d      (hw2reg.err_code.sfifo_blkenc_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_blkenc_err_qs)
  );

  //   F[cmd_stage_sm_err]: 20:20
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_cmd_stage_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.cmd_stage_sm_err.de),
    .d      (hw2reg.err_code.cmd_stage_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_cmd_stage_sm_err_qs)
  );

  //   F[main_sm_err]: 21:21
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_main_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.main_sm_err.de),
    .d      (hw2reg.err_code.main_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_main_sm_err_qs)
  );

  //   F[drbg_gen_sm_err]: 22:22
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_drbg_gen_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.drbg_gen_sm_err.de),
    .d      (hw2reg.err_code.drbg_gen_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_drbg_gen_sm_err_qs)
  );

  //   F[drbg_updbe_sm_err]: 23:23
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_drbg_updbe_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.drbg_updbe_sm_err.de),
    .d      (hw2reg.err_code.drbg_updbe_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_drbg_updbe_sm_err_qs)
  );

  //   F[drbg_updob_sm_err]: 24:24
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_drbg_updob_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.drbg_updob_sm_err.de),
    .d      (hw2reg.err_code.drbg_updob_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_drbg_updob_sm_err_qs)
  );

  //   F[aes_cipher_sm_err]: 25:25
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_aes_cipher_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.aes_cipher_sm_err.de),
    .d      (hw2reg.err_code.aes_cipher_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_aes_cipher_sm_err_qs)
  );

  //   F[cmd_gen_cnt_err]: 26:26
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_cmd_gen_cnt_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.cmd_gen_cnt_err.de),
    .d      (hw2reg.err_code.cmd_gen_cnt_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_cmd_gen_cnt_err_qs)
  );

  //   F[fifo_write_err]: 28:28
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_write_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_write_err.de),
    .d      (hw2reg.err_code.fifo_write_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_write_err_qs)
  );

  //   F[fifo_read_err]: 29:29
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_read_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_read_err.de),
    .d      (hw2reg.err_code.fifo_read_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_read_err_qs)
  );

  //   F[fifo_state_err]: 30:30
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_state_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_state_err.de),
    .d      (hw2reg.err_code.fifo_state_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_state_err_qs)
  );


  // R[err_code_test]: V(False)
  logic err_code_test_qe;
  logic [0:0] err_code_test_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_err_code_test0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&err_code_test_flds_we),
    .q_o(err_code_test_qe)
  );
  // Create REGWEN-gated WE signal
  logic err_code_test_gated_we;
  assign err_code_test_gated_we = err_code_test_we & regwen_qs;
  prim_subreg #(
    .DW      (5),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (5'h0)
  ) u_err_code_test (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (err_code_test_gated_we),
    .wd     (err_code_test_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (err_code_test_flds_we[0]),
    .q      (reg2hw.err_code_test.q),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_test_qs)
  );
  assign reg2hw.err_code_test.qe = err_code_test_qe;


  // R[main_sm_state]: V(False)
  prim_subreg #(
    .DW      (8),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (8'h4e)
  ) u_main_sm_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.main_sm_state.de),
    .d      (hw2reg.main_sm_state.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (main_sm_state_qs)
  );



  logic [16:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == CSRNG_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == CSRNG_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == CSRNG_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == CSRNG_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == CSRNG_REGWEN_OFFSET);
    addr_hit[ 5] = (reg_addr == CSRNG_CTRL_OFFSET);
    addr_hit[ 6] = (reg_addr == CSRNG_CMD_REQ_OFFSET);
    addr_hit[ 7] = (reg_addr == CSRNG_SW_CMD_STS_OFFSET);
    addr_hit[ 8] = (reg_addr == CSRNG_GENBITS_VLD_OFFSET);
    addr_hit[ 9] = (reg_addr == CSRNG_GENBITS_OFFSET);
    addr_hit[10] = (reg_addr == CSRNG_INT_STATE_NUM_OFFSET);
    addr_hit[11] = (reg_addr == CSRNG_INT_STATE_VAL_OFFSET);
    addr_hit[12] = (reg_addr == CSRNG_HW_EXC_STS_OFFSET);
    addr_hit[13] = (reg_addr == CSRNG_RECOV_ALERT_STS_OFFSET);
    addr_hit[14] = (reg_addr == CSRNG_ERR_CODE_OFFSET);
    addr_hit[15] = (reg_addr == CSRNG_ERR_CODE_TEST_OFFSET);
    addr_hit[16] = (reg_addr == CSRNG_MAIN_SM_STATE_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(CSRNG_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(CSRNG_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(CSRNG_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(CSRNG_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(CSRNG_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(CSRNG_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(CSRNG_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(CSRNG_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(CSRNG_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(CSRNG_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(CSRNG_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(CSRNG_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(CSRNG_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(CSRNG_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(CSRNG_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(CSRNG_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(CSRNG_PERMIT[16] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_cs_cmd_req_done_wd = reg_wdata[0];

  assign intr_state_cs_entropy_req_wd = reg_wdata[1];

  assign intr_state_cs_hw_inst_exc_wd = reg_wdata[2];

  assign intr_state_cs_fatal_err_wd = reg_wdata[3];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_cs_cmd_req_done_wd = reg_wdata[0];

  assign intr_enable_cs_entropy_req_wd = reg_wdata[1];

  assign intr_enable_cs_hw_inst_exc_wd = reg_wdata[2];

  assign intr_enable_cs_fatal_err_wd = reg_wdata[3];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_cs_cmd_req_done_wd = reg_wdata[0];

  assign intr_test_cs_entropy_req_wd = reg_wdata[1];

  assign intr_test_cs_hw_inst_exc_wd = reg_wdata[2];

  assign intr_test_cs_fatal_err_wd = reg_wdata[3];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_recov_alert_wd = reg_wdata[0];

  assign alert_test_fatal_alert_wd = reg_wdata[1];
  assign regwen_we = addr_hit[4] & reg_we & !reg_error;

  assign regwen_wd = reg_wdata[0];
  assign ctrl_we = addr_hit[5] & reg_we & !reg_error;

  assign ctrl_enable_wd = reg_wdata[3:0];

  assign ctrl_sw_app_enable_wd = reg_wdata[7:4];

  assign ctrl_read_int_state_wd = reg_wdata[11:8];
  assign cmd_req_we = addr_hit[6] & reg_we & !reg_error;

  assign cmd_req_wd = reg_wdata[31:0];
  assign genbits_vld_re = addr_hit[8] & reg_re & !reg_error;
  assign genbits_re = addr_hit[9] & reg_re & !reg_error;
  assign int_state_num_we = addr_hit[10] & reg_we & !reg_error;

  assign int_state_num_wd = reg_wdata[3:0];
  assign int_state_val_re = addr_hit[11] & reg_re & !reg_error;
  assign hw_exc_sts_we = addr_hit[12] & reg_we & !reg_error;

  assign hw_exc_sts_wd = reg_wdata[15:0];
  assign recov_alert_sts_we = addr_hit[13] & reg_we & !reg_error;

  assign recov_alert_sts_enable_field_alert_wd = reg_wdata[0];

  assign recov_alert_sts_sw_app_enable_field_alert_wd = reg_wdata[1];

  assign recov_alert_sts_read_int_state_field_alert_wd = reg_wdata[2];

  assign recov_alert_sts_acmd_flag0_field_alert_wd = reg_wdata[3];

  assign recov_alert_sts_cs_bus_cmp_alert_wd = reg_wdata[12];

  assign recov_alert_sts_cs_main_sm_alert_wd = reg_wdata[13];
  assign err_code_test_we = addr_hit[15] & reg_we & !reg_error;

  assign err_code_test_wd = reg_wdata[4:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = regwen_we;
    reg_we_check[5] = ctrl_gated_we;
    reg_we_check[6] = cmd_req_we;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = 1'b0;
    reg_we_check[9] = 1'b0;
    reg_we_check[10] = int_state_num_we;
    reg_we_check[11] = 1'b0;
    reg_we_check[12] = hw_exc_sts_we;
    reg_we_check[13] = recov_alert_sts_we;
    reg_we_check[14] = 1'b0;
    reg_we_check[15] = err_code_test_gated_we;
    reg_we_check[16] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_cs_cmd_req_done_qs;
        reg_rdata_next[1] = intr_state_cs_entropy_req_qs;
        reg_rdata_next[2] = intr_state_cs_hw_inst_exc_qs;
        reg_rdata_next[3] = intr_state_cs_fatal_err_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_cs_cmd_req_done_qs;
        reg_rdata_next[1] = intr_enable_cs_entropy_req_qs;
        reg_rdata_next[2] = intr_enable_cs_hw_inst_exc_qs;
        reg_rdata_next[3] = intr_enable_cs_fatal_err_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
        reg_rdata_next[2] = '0;
        reg_rdata_next[3] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[0] = regwen_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[3:0] = ctrl_enable_qs;
        reg_rdata_next[7:4] = ctrl_sw_app_enable_qs;
        reg_rdata_next[11:8] = ctrl_read_int_state_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[7]: begin
        reg_rdata_next[0] = sw_cmd_sts_cmd_rdy_qs;
        reg_rdata_next[1] = sw_cmd_sts_cmd_sts_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[0] = genbits_vld_genbits_vld_qs;
        reg_rdata_next[1] = genbits_vld_genbits_fips_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = genbits_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[3:0] = int_state_num_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = int_state_val_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[15:0] = hw_exc_sts_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[0] = recov_alert_sts_enable_field_alert_qs;
        reg_rdata_next[1] = recov_alert_sts_sw_app_enable_field_alert_qs;
        reg_rdata_next[2] = recov_alert_sts_read_int_state_field_alert_qs;
        reg_rdata_next[3] = recov_alert_sts_acmd_flag0_field_alert_qs;
        reg_rdata_next[12] = recov_alert_sts_cs_bus_cmp_alert_qs;
        reg_rdata_next[13] = recov_alert_sts_cs_main_sm_alert_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[0] = err_code_sfifo_cmd_err_qs;
        reg_rdata_next[1] = err_code_sfifo_genbits_err_qs;
        reg_rdata_next[2] = err_code_sfifo_cmdreq_err_qs;
        reg_rdata_next[3] = err_code_sfifo_rcstage_err_qs;
        reg_rdata_next[4] = err_code_sfifo_keyvrc_err_qs;
        reg_rdata_next[5] = err_code_sfifo_updreq_err_qs;
        reg_rdata_next[6] = err_code_sfifo_bencreq_err_qs;
        reg_rdata_next[7] = err_code_sfifo_bencack_err_qs;
        reg_rdata_next[8] = err_code_sfifo_pdata_err_qs;
        reg_rdata_next[9] = err_code_sfifo_final_err_qs;
        reg_rdata_next[10] = err_code_sfifo_gbencack_err_qs;
        reg_rdata_next[11] = err_code_sfifo_grcstage_err_qs;
        reg_rdata_next[12] = err_code_sfifo_ggenreq_err_qs;
        reg_rdata_next[13] = err_code_sfifo_gadstage_err_qs;
        reg_rdata_next[14] = err_code_sfifo_ggenbits_err_qs;
        reg_rdata_next[15] = err_code_sfifo_blkenc_err_qs;
        reg_rdata_next[20] = err_code_cmd_stage_sm_err_qs;
        reg_rdata_next[21] = err_code_main_sm_err_qs;
        reg_rdata_next[22] = err_code_drbg_gen_sm_err_qs;
        reg_rdata_next[23] = err_code_drbg_updbe_sm_err_qs;
        reg_rdata_next[24] = err_code_drbg_updob_sm_err_qs;
        reg_rdata_next[25] = err_code_aes_cipher_sm_err_qs;
        reg_rdata_next[26] = err_code_cmd_gen_cnt_err_qs;
        reg_rdata_next[28] = err_code_fifo_write_err_qs;
        reg_rdata_next[29] = err_code_fifo_read_err_qs;
        reg_rdata_next[30] = err_code_fifo_state_err_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[4:0] = err_code_test_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[7:0] = main_sm_state_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng app cmd request state machine module
//
//  - handles all app cmd requests from all requesting interfaces

module csrng_main_sm import csrng_pkg::*; #() (
  input logic                         clk_i,
  input logic                         rst_ni,

  input logic                         enable_i,
  input logic                         acmd_avail_i,
  output logic                        acmd_accept_o,
  input logic [2:0]                   acmd_i,
  input logic                         acmd_eop_i,
  input logic                         ctr_drbg_cmd_req_rdy_i,
  input logic                         flag0_i,
  output logic                        cmd_entropy_req_o,
  input logic                         cmd_entropy_avail_i,
  output logic                        instant_req_o,
  output logic                        reseed_req_o,
  output logic                        generate_req_o,
  output logic                        update_req_o,
  output logic                        uninstant_req_o,
  output logic                        clr_adata_packer_o,
  input logic                         cmd_complete_i,
  input logic                         local_escalate_i,
  output logic [MainSmStateWidth-1:0] main_sm_state_o,
  output logic                        main_sm_alert_o,
  output logic                        main_sm_err_o
);

  main_sm_state_e state_d, state_q;
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, main_sm_state_e, MainSmIdle)

  assign main_sm_state_o = {state_q};

  always_comb begin
    state_d            = state_q;
    acmd_accept_o      = 1'b0;
    cmd_entropy_req_o  = 1'b0;
    instant_req_o      = 1'b0;
    reseed_req_o       = 1'b0;
    generate_req_o     = 1'b0;
    update_req_o       = 1'b0;
    uninstant_req_o    = 1'b0;
    clr_adata_packer_o = 1'b0;
    main_sm_alert_o    = 1'b0;
    main_sm_err_o      = 1'b0;

    if (state_q == MainSmError) begin
      // In case we are in the Error state we must ignore the local escalate and enable signals.
      main_sm_err_o = 1'b1;
    end else if (local_escalate_i) begin
      // In case local escalate is high we must transition to the error state.
      state_d = MainSmError;
    end else if (!enable_i && state_q inside {MainSmIdle, MainSmParseCmd, MainSmInstantPrep,
                                              MainSmInstantReq, MainSmReseedPrep, MainSmReseedReq,
                                              MainSmGeneratePrep, MainSmGenerateReq,
                                              MainSmUpdatePrep, MainSmUpdateReq,
                                              MainSmUninstantPrep, MainSmUninstantReq,
                                              MainSmClrAData, MainSmCmdCompWait}) begin
      // In case the module is disabled and we are in a legal state we must go into idle state.
      state_d = MainSmIdle;
    end else begin
      // Otherwise do the state machine as normal.
      unique case (state_q)
        MainSmIdle: begin
          // Because of the if statement above we won't leave idle if enable is low.
          if (ctr_drbg_cmd_req_rdy_i) begin
            // Signal the arbiter to grant this request.
            if (acmd_avail_i) begin
              acmd_accept_o = 1'b1;
              state_d = MainSmParseCmd;
            end
          end
        end
        MainSmParseCmd: begin
          if (ctr_drbg_cmd_req_rdy_i) begin
            if (acmd_i == INS) begin
              if (acmd_eop_i) begin
                state_d = MainSmInstantPrep;
              end
            end else if (acmd_i == RES) begin
              if (acmd_eop_i) begin
                state_d = MainSmReseedPrep;
              end
            end else if (acmd_i == GEN) begin
              if (acmd_eop_i) begin
                state_d = MainSmGeneratePrep;
              end
            end else if (acmd_i == UPD) begin
              if (acmd_eop_i) begin
                state_d = MainSmUpdatePrep;
              end
            end else if (acmd_i == UNI) begin
              if (acmd_eop_i) begin
                state_d = MainSmUninstantPrep;
              end
            end else begin
              // Command was not supported.
              main_sm_alert_o = 1'b1;
            end
          end
        end
        MainSmInstantPrep: begin
          if (flag0_i) begin
            // Assumes all adata is present now.
            state_d = MainSmInstantReq;
          end else begin
            // Delay one clock to fix timing issue.
            cmd_entropy_req_o = 1'b1;
            if (cmd_entropy_avail_i) begin
              state_d = MainSmInstantReq;
            end
          end
        end
        MainSmInstantReq: begin
          instant_req_o = 1'b1;
          state_d = MainSmClrAData;
        end
        MainSmReseedPrep: begin
          if (flag0_i) begin
            // Assumes all adata is present now.
            state_d = MainSmReseedReq;
          end else begin
            // Delay one clock to fix timing issue.
            cmd_entropy_req_o = 1'b1;
            if (cmd_entropy_avail_i) begin
              state_d = MainSmReseedReq;
            end
          end
        end
        MainSmReseedReq: begin
          reseed_req_o = 1'b1;
          state_d = MainSmClrAData;
        end
        MainSmGeneratePrep: begin
          // Assumes all adata is present now.
          state_d = MainSmGenerateReq;
        end
        MainSmGenerateReq: begin
          generate_req_o = 1'b1;
          state_d = MainSmClrAData;
        end
        MainSmUpdatePrep: begin
          // Assumes all adata is present now.
          state_d = MainSmUpdateReq;
        end
        MainSmUpdateReq: begin
          update_req_o = 1'b1;
          state_d = MainSmClrAData;
        end
        MainSmUninstantPrep: begin
          // Assumes all adata is present now.
          state_d = MainSmUninstantReq;
        end
        MainSmUninstantReq: begin
          uninstant_req_o = 1'b1;
          state_d = MainSmClrAData;
        end
        MainSmClrAData: begin
          clr_adata_packer_o = 1'b1;
          state_d = MainSmCmdCompWait;
        end
        MainSmCmdCompWait: begin
          if (cmd_complete_i) begin
            state_d = MainSmIdle;
          end
        end
        // Error: The error state is now covered by the if statement above.
        default: begin
          state_d = MainSmError;
          main_sm_err_o = 1'b1;
        end
      endcase
    end
  end

  // Make sure that the state machine has a stable error state. This means that after the error
  // state is entered it will not exit it unless a reset signal is received.
  `ASSERT(CsrngMainErrorStStable_A, state_q == MainSmError |=> $stable(state_q))
  // If in error state, the error output must be high.
  `ASSERT(CsrngMainErrorOutput_A,   state_q == MainSmError |-> main_sm_err_o)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng state data base module
//
// This is the container for accessing the current
//    working state for a given drbg instance.

`include "prim_assert.sv"

module csrng_state_db import csrng_pkg::*; #(
  parameter int NApps = 4,
  parameter int StateId = 4,
  parameter int BlkLen = 128,
  parameter int KeyLen = 256,
  parameter int CtrLen  = 32,
  parameter int Cmd     = 3
) (
  input logic                clk_i,
  input logic                rst_ni,

   // read interface
  input logic                state_db_enable_i,
  input logic [StateId-1:0]  state_db_rd_inst_id_i,
  output logic [KeyLen-1:0]  state_db_rd_key_o,
  output logic [BlkLen-1:0]  state_db_rd_v_o,
  output logic [CtrLen-1:0]  state_db_rd_res_ctr_o,
  output logic               state_db_rd_inst_st_o,
  output logic               state_db_rd_fips_o,
  // write interface
  input logic                state_db_wr_req_i,
  output logic               state_db_wr_req_rdy_o,
  input logic [StateId-1:0]  state_db_wr_inst_id_i,
  input logic                state_db_wr_fips_i,
  input logic [Cmd-1:0]      state_db_wr_ccmd_i,
  input logic [KeyLen-1:0]   state_db_wr_key_i,
  input logic [BlkLen-1:0]   state_db_wr_v_i,
  input logic [CtrLen-1:0]   state_db_wr_res_ctr_i,
  input logic                state_db_wr_sts_i,
  // status interface
  input logic                state_db_is_dump_en_i,
  input logic                state_db_reg_rd_sel_i,
  input logic                state_db_reg_rd_id_pulse_i,
  input logic [StateId-1:0]  state_db_reg_rd_id_i,
  output logic [31:0]        state_db_reg_rd_val_o,
  output logic               state_db_sts_ack_o,
  output logic               state_db_sts_sts_o,
  output logic [StateId-1:0] state_db_sts_id_o
);

  localparam int InternalStateWidth = 2+KeyLen+BlkLen+CtrLen;
  localparam int RegInternalStateWidth = 30+InternalStateWidth;
  localparam int RegW = 32;
  localparam int StateWidth = 1+1+KeyLen+BlkLen+CtrLen+StateId+1;

  logic [StateId-1:0]              state_db_id;
  logic [KeyLen-1:0]               state_db_key;
  logic [BlkLen-1:0]               state_db_v;
  logic [CtrLen-1:0]               state_db_rc;
  logic                            state_db_fips;
  logic                            state_db_inst_st;
  logic                            state_db_sts;
  logic                            state_db_write;
  logic                            instance_status;
  logic [NApps-1:0]                int_st_out_sel;
  logic [NApps-1:0]                int_st_dump_sel;
  logic [InternalStateWidth-1:0]   internal_states_out[NApps];
  logic [InternalStateWidth-1:0]   internal_states_dump[NApps];
  logic [RegInternalStateWidth-1:0] internal_state_diag;
  logic                             reg_rd_ptr_inc;

  // flops
  logic                            state_db_sts_ack_q, state_db_sts_ack_d;
  logic                            state_db_sts_sts_q, state_db_sts_sts_d;
  logic [StateId-1:0]              state_db_sts_id_q, state_db_sts_id_d;
  logic [StateId-1:0]              reg_rd_ptr_q, reg_rd_ptr_d;
  logic [StateId-1:0]              int_st_dump_id_q, int_st_dump_id_d;

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      state_db_sts_ack_q   <= '0;
      state_db_sts_sts_q   <= '0;
      state_db_sts_id_q    <= '0;
      reg_rd_ptr_q         <= '0;
      int_st_dump_id_q     <= '0;
    end else begin
      state_db_sts_ack_q   <= state_db_sts_ack_d;
      state_db_sts_sts_q   <= state_db_sts_sts_d;
      state_db_sts_id_q    <= state_db_sts_id_d;
      reg_rd_ptr_q         <= reg_rd_ptr_d;
      int_st_dump_id_q     <= int_st_dump_id_d;
    end

  // flops - no reset
  logic [InternalStateWidth-1:0]  internal_states_q[NApps], internal_states_d[NApps];
  logic [InternalStateWidth-1:0]  internal_state_pl_q, internal_state_pl_d;
  logic [InternalStateWidth-1:0]  internal_state_pl_dump_q, internal_state_pl_dump_d;


  // no reset on state
  always_ff @(posedge clk_i)
    begin
      internal_states_q <= internal_states_d;
      internal_state_pl_q <= internal_state_pl_d;
      internal_state_pl_dump_q <= internal_state_pl_dump_d;
    end


  //--------------------------------------------
  // internal state read logic
  //--------------------------------------------
  for (genvar rd = 0; rd < NApps; rd = rd+1) begin : gen_state_rd
    assign int_st_out_sel[rd] = (state_db_rd_inst_id_i == rd);
    assign int_st_dump_sel[rd] = (int_st_dump_id_q == rd);
    assign internal_states_out[rd] = int_st_out_sel[rd] ? internal_states_q[rd] : '0;
    assign internal_states_dump[rd] = int_st_dump_sel[rd] ? internal_states_q[rd] : '0;
  end

  // since only one of the internal states is active at a time, a
  // logical "or" is made of all of the buses into one
  always_comb begin
    internal_state_pl_d = '0;
    internal_state_pl_dump_d = '0;
    for (int i = 0; i < NApps; i = i+1) begin
      internal_state_pl_d |= internal_states_out[i];
      internal_state_pl_dump_d |= internal_states_dump[i];
    end
  end

  assign {state_db_rd_fips_o,state_db_rd_inst_st_o,
          state_db_rd_key_o,state_db_rd_v_o,
          state_db_rd_res_ctr_o} = internal_state_pl_q;


  // using a copy of the internal state pipeline version for better timing
  assign internal_state_diag = {30'b0,internal_state_pl_dump_q};


  // Register access of internal state
  assign state_db_reg_rd_val_o =
         (reg_rd_ptr_q == 4'h0) ? internal_state_diag[RegW-1:0] :
         (reg_rd_ptr_q == 4'h1) ? internal_state_diag[2*RegW-1:RegW] :
         (reg_rd_ptr_q == 4'h2) ? internal_state_diag[3*RegW-1:2*RegW] :
         (reg_rd_ptr_q == 4'h3) ? internal_state_diag[4*RegW-1:3*RegW] :
         (reg_rd_ptr_q == 4'h4) ? internal_state_diag[5*RegW-1:4*RegW] :
         (reg_rd_ptr_q == 4'h5) ? internal_state_diag[6*RegW-1:5*RegW] :
         (reg_rd_ptr_q == 4'h6) ? internal_state_diag[7*RegW-1:6*RegW] :
         (reg_rd_ptr_q == 4'h7) ? internal_state_diag[8*RegW-1:7*RegW] :
         (reg_rd_ptr_q == 4'h8) ? internal_state_diag[9*RegW-1:8*RegW] :
         (reg_rd_ptr_q == 4'h9) ? internal_state_diag[10*RegW-1:9*RegW] :
         (reg_rd_ptr_q == 4'ha) ? internal_state_diag[11*RegW-1:10*RegW] :
         (reg_rd_ptr_q == 4'hb) ? internal_state_diag[12*RegW-1:11*RegW] :
         (reg_rd_ptr_q == 4'hc) ? internal_state_diag[13*RegW-1:12*RegW] :
         (reg_rd_ptr_q == 4'hd) ? internal_state_diag[14*RegW-1:13*RegW] :
         '0;

  // selects 32b fields from the internal state to be read out for diagnostics
  assign reg_rd_ptr_inc = state_db_reg_rd_sel_i;

  assign reg_rd_ptr_d =
         (!state_db_enable_i) ? 4'hf :
         (!state_db_is_dump_en_i) ? 4'hf :
         (reg_rd_ptr_q == 4'he) ? '0 :
         state_db_reg_rd_id_pulse_i ? '0 :
         reg_rd_ptr_inc ? (reg_rd_ptr_q+1) :
         reg_rd_ptr_q;


  assign int_st_dump_id_d =
         (!state_db_enable_i) ? '0 :
         state_db_reg_rd_id_pulse_i ? state_db_reg_rd_id_i :
         int_st_dump_id_q;

  //--------------------------------------------
  // write state logic
  //--------------------------------------------

  for (genvar wr = 0; wr < NApps; wr = wr+1) begin : gen_state_wr

    assign internal_states_d[wr] = !state_db_enable_i ? '0 : // better timing
                                   (state_db_write && (state_db_id == wr)) ?
                                   {state_db_fips,state_db_inst_st,state_db_key,
                                    state_db_v,state_db_rc} : internal_states_q[wr];
  end : gen_state_wr


  assign {state_db_fips,state_db_inst_st,
          state_db_key,
          state_db_v,state_db_rc,
          state_db_id,state_db_sts} = {StateWidth{state_db_enable_i}} &
                                      {state_db_wr_fips_i,instance_status,
                                       state_db_wr_key_i,
                                       state_db_wr_v_i,state_db_wr_res_ctr_i,
                                       state_db_wr_inst_id_i,state_db_wr_sts_i};

  assign instance_status =
         (state_db_wr_ccmd_i == INS) ||
         (state_db_wr_ccmd_i == RES) ||
         (state_db_wr_ccmd_i == GENU) ||
         (state_db_wr_ccmd_i == UPD);


  assign state_db_write = state_db_enable_i && state_db_wr_req_i;

  assign state_db_sts_ack_d =
         state_db_write;

  assign state_db_sts_sts_d =
         state_db_sts;

  assign state_db_sts_id_d =
         state_db_id;

  assign state_db_sts_ack_o = state_db_sts_ack_q;
  assign state_db_sts_sts_o = state_db_sts_sts_q;
  assign state_db_sts_id_o = state_db_sts_id_q;
  assign state_db_wr_req_rdy_o = 1'b1;


  // Assertions
  `ASSERT_KNOWN(IntStOutSelOneHot_A, $onehot(int_st_out_sel))

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: CSRNG command staging module.
//

module csrng_cmd_stage import csrng_pkg::*; #(
  parameter int CmdFifoWidth = 32,
  parameter int CmdFifoDepth = 16,
  parameter int StateId = 4
) (
  input logic                        clk_i,
  input logic                        rst_ni,
  // Command input.
  input logic                        cs_enable_i,
  input logic                        cmd_stage_vld_i,
  input logic [StateId-1:0]          cmd_stage_shid_i,
  input logic [CmdFifoWidth-1:0]     cmd_stage_bus_i,
  output logic                       cmd_stage_rdy_o,
  // Command to arbiter.
  output logic                       cmd_arb_req_o,
  output logic                       cmd_arb_sop_o,
  output logic                       cmd_arb_mop_o,
  output logic                       cmd_arb_eop_o,
  input logic                        cmd_arb_gnt_i,
  output logic [CmdFifoWidth-1:0]    cmd_arb_bus_o,
  // Ack from core.
  input logic                        cmd_ack_i,
  input logic                        cmd_ack_sts_i,
  // Ack to app i/f.
  output logic                       cmd_stage_ack_o,
  output logic                       cmd_stage_ack_sts_o,
  // Genbits from core.
  input logic                        genbits_vld_i,
  input logic [127:0]                genbits_bus_i,
  input logic                        genbits_fips_i,
  // Genbits to app i/f.
  output logic                       genbits_vld_o,
  input logic                        genbits_rdy_i,
  output logic [127:0]               genbits_bus_o,
  output logic                       genbits_fips_o,
  // Error indication.
  output logic [2:0]                 cmd_stage_sfifo_cmd_err_o,
  output logic [2:0]                 cmd_stage_sfifo_genbits_err_o,
  output logic                       cmd_gen_cnt_err_o,
  output logic                       cmd_stage_sm_err_o
);

  // Genbits parameters.
  localparam int GenBitsFifoWidth = 1+128;
  localparam int GenBitsFifoDepth = 1;
  localparam int GenBitsCntrWidth = 12;

  // Command FIFO.
  logic [CmdFifoWidth-1:0] sfifo_cmd_rdata;
  logic [$clog2(CmdFifoDepth):0] sfifo_cmd_depth;
  logic                    sfifo_cmd_push;
  logic [CmdFifoWidth-1:0] sfifo_cmd_wdata;
  logic                    sfifo_cmd_pop;
  logic [2:0]              sfifo_cmd_err;
  logic                    sfifo_cmd_full;
  logic                    sfifo_cmd_not_empty;

  // Genbits FIFO.
  logic [GenBitsFifoWidth-1:0] sfifo_genbits_rdata;
  logic                        sfifo_genbits_push;
  logic [GenBitsFifoWidth-1:0] sfifo_genbits_wdata;
  logic                        sfifo_genbits_pop;
  logic [2:0]                  sfifo_genbits_err;
  logic                        sfifo_genbits_full;
  logic                        sfifo_genbits_not_empty;

  // Command signals.
  logic [3:0]              cmd_len;
  logic                    cmd_fifo_zero;
  logic                    cmd_fifo_pop;
  logic                    cmd_len_dec;
  logic                    cmd_gen_cnt_dec;
  logic                    cmd_gen_1st_req;
  logic                    cmd_gen_inc_req;
  logic                    cmd_gen_cnt_last;
  logic                    cmd_final_ack;
  logic [GenBitsCntrWidth-1:0] cmd_gen_cnt;

  // Flops.
  logic                    cmd_ack_q, cmd_ack_d;
  logic                    cmd_ack_sts_q, cmd_ack_sts_d;
  logic [3:0]              cmd_len_q, cmd_len_d;
  logic                    cmd_gen_flag_q, cmd_gen_flag_d;
  logic [11:0]             cmd_gen_cmd_q, cmd_gen_cmd_d;

  logic                    local_escalate;


  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      cmd_ack_q       <= '0;
      cmd_ack_sts_q   <= '0;
      cmd_len_q       <= '0;
      cmd_gen_flag_q  <= '0;
      cmd_gen_cmd_q   <= '0;
    end else begin
      cmd_ack_q       <= cmd_ack_d;
      cmd_ack_sts_q   <= cmd_ack_sts_d;
      cmd_len_q       <= cmd_len_d;
      cmd_gen_flag_q  <= cmd_gen_flag_d;
      cmd_gen_cmd_q   <= cmd_gen_cmd_d;
    end

  assign  cmd_stage_sfifo_cmd_err_o = sfifo_cmd_err;
  assign  cmd_stage_sfifo_genbits_err_o = sfifo_genbits_err;

  //---------------------------------------------------------
  // Capture the transfer length of data behind the command.
  //---------------------------------------------------------

  prim_fifo_sync #(
    .Width(CmdFifoWidth),
    .Pass(0),
    .Depth(CmdFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_cmd (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!cs_enable_i),
    .wvalid_i       (sfifo_cmd_push),
    .wready_o       (),
    .wdata_i        (sfifo_cmd_wdata),
    .rvalid_o       (sfifo_cmd_not_empty),
    .rready_i       (sfifo_cmd_pop),
    .rdata_o        (sfifo_cmd_rdata),
    .full_o         (sfifo_cmd_full),
    .depth_o        (sfifo_cmd_depth),
    .err_o          ()
  );

  assign sfifo_cmd_wdata = cmd_stage_bus_i;

  assign sfifo_cmd_push = cs_enable_i && cmd_stage_rdy_o && cmd_stage_vld_i;

  assign sfifo_cmd_pop = cs_enable_i && cmd_fifo_pop;

  assign cmd_arb_bus_o =
         cmd_gen_inc_req ? {15'b0,cmd_gen_cnt_last,cmd_stage_shid_i,cmd_gen_cmd_q} :
        // pad,glast,id,f,clen,cmd
        cmd_gen_1st_req ? {15'b0,cmd_gen_cnt_last,cmd_stage_shid_i,sfifo_cmd_rdata[11:0]} :
        cmd_arb_mop_o   ? sfifo_cmd_rdata :
        '0;

  assign cmd_stage_rdy_o = !sfifo_cmd_full;

  assign sfifo_cmd_err =
         {(sfifo_cmd_push && sfifo_cmd_full),
          (sfifo_cmd_pop && !sfifo_cmd_not_empty),
          (sfifo_cmd_full && !sfifo_cmd_not_empty)};


  // State machine controls.
  assign cmd_fifo_zero = (sfifo_cmd_depth == '0);
  assign cmd_len = sfifo_cmd_rdata[7:4];

  // Capture the length of csrng command.
  assign cmd_len_d =
         (!cs_enable_i) ? '0 :
         cmd_arb_sop_o ? cmd_len :
         cmd_len_dec ? (cmd_len_q-1) :
         cmd_len_q;

  // For gen commands, capture information from the orignal command for use later.
  assign cmd_gen_flag_d =
         (!cs_enable_i) ? '0 :
         cmd_gen_1st_req ? (sfifo_cmd_rdata[2:0] == GEN) :
         cmd_gen_flag_q;

  assign cmd_gen_cmd_d =
         (!cs_enable_i) ? '0 :
         cmd_gen_1st_req ? {sfifo_cmd_rdata[11:0]} :
         cmd_gen_cmd_q;

  // SEC_CM: GEN_CMD.CTR.REDUN
  prim_count #(
    .Width(GenBitsCntrWidth),
    .ResetValue({GenBitsCntrWidth{1'b1}})
  ) u_prim_count_cmd_gen_cntr (
    .clk_i,
    .rst_ni,
    .clr_i(!cs_enable_i),
    .set_i(cmd_gen_1st_req),
    .set_cnt_i(sfifo_cmd_rdata[12+:GenBitsCntrWidth]),
    .incr_en_i(1'b0),
    .decr_en_i(cmd_gen_cnt_dec), // Count down.
    .step_i(GenBitsCntrWidth'(1)),
    .cnt_o(cmd_gen_cnt),
    .cnt_next_o(),
    .err_o(cmd_gen_cnt_err_o)
  );

  // For naming consistency.
  assign local_escalate = cmd_gen_cnt_err_o;

  //---------------------------------------------------------
  // state machine to process command
  //---------------------------------------------------------
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 10 -n 8 \
  //      -s 170131814 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||| (28.89%)
  //  4: |||||||||||||||||||| (35.56%)
  //  5: |||||||||||| (22.22%)
  //  6: ||||| (8.89%)
  //  7: | (2.22%)
  //  8: | (2.22%)
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 8
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 7
  //
  localparam int StateWidth = 8;
  typedef    enum logic [StateWidth-1:0] {
    Idle      = 8'b00011011, // idle
    ArbGnt    = 8'b11110101, // general arbiter request
    SendSOP   = 8'b00011100, // send sop (start of packet)
    SendMOP   = 8'b00000001, // send mop (middle of packet)
    GenCmdChk = 8'b01010110, // gen cmd check
    CmdAck    = 8'b10001101, // wait for command ack
    GenReq    = 8'b11000000, // process gen requests
    GenArbGnt = 8'b11111110, // generate subsequent arb request
    GenSOP    = 8'b10110010, // generate subsequent request
    Error     = 8'b10111001  // illegal state reached and hang
  } state_e;

  state_e state_d, state_q;
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, Idle)

  always_comb begin
    state_d = state_q;
    cmd_fifo_pop = 1'b0;
    cmd_len_dec = 1'b0;
    cmd_gen_cnt_dec = 1'b0;
    cmd_gen_1st_req = 1'b0;
    cmd_gen_inc_req = 1'b0;
    cmd_gen_cnt_last = 1'b0;
    cmd_final_ack = 1'b0;
    cmd_arb_req_o = 1'b0;
    cmd_arb_sop_o = 1'b0;
    cmd_arb_mop_o = 1'b0;
    cmd_arb_eop_o = 1'b0;
    cmd_stage_sm_err_o = 1'b0;

    if (state_q == Error) begin
      // In case we are in the Error state we must ignore the local escalate and enable signals.
      cmd_stage_sm_err_o = 1'b1;
    end else if (local_escalate) begin
      // In case local escalate is high we must transition to the error state.
      state_d = Error;
    end else if (!cs_enable_i && state_q inside {Idle, ArbGnt, SendSOP, SendMOP, GenCmdChk, CmdAck,
                                                 GenReq, GenArbGnt, GenSOP}) begin
      // In case the module is disabled and we are in a legal state we must go into idle state.
      state_d = Idle;
    end else begin
      // Otherwise do the state machine as normal.
      unique case (state_q)
        Idle: begin
          // Because of the if statement above we won't leave idle if enable is low.
          if (!cmd_fifo_zero) begin
            state_d = ArbGnt;
          end
        end
        ArbGnt: begin
          cmd_arb_req_o = 1'b1;
          if (cmd_arb_gnt_i) begin
            state_d = SendSOP;
          end
        end
        SendSOP: begin
          cmd_gen_1st_req = 1'b1;
          cmd_arb_sop_o = 1'b1;
          cmd_fifo_pop = 1'b1;
          if (sfifo_cmd_rdata[12+:GenBitsCntrWidth] == GenBitsCntrWidth'(1)) begin
            cmd_gen_cnt_last = 1'b1;
          end
          if (cmd_len == '0) begin
            cmd_arb_eop_o = 1'b1;
            state_d = GenCmdChk;
          end else begin
            state_d = SendMOP;
          end
        end
        SendMOP: begin
          if (!cmd_fifo_zero) begin
            cmd_fifo_pop = 1'b1;
            cmd_len_dec = 1'b1;
            if (cmd_len_q == 4'h1) begin
              cmd_arb_mop_o = 1'b1;
              cmd_arb_eop_o = 1'b1;
              state_d = GenCmdChk;
            end else begin
              cmd_arb_mop_o = 1'b1;
            end
          end
        end
        GenCmdChk: begin
          if (cmd_gen_flag_q) begin
            cmd_gen_cnt_dec= 1'b1;
          end
          state_d = CmdAck;
        end
        CmdAck: begin
          if (cmd_ack_i) begin
            state_d = GenReq;
          end
        end
        GenReq: begin
          // Flag set if a gen request.
          if (cmd_gen_flag_q) begin
            // Must stall if genbits fifo is not clear.
            if (!sfifo_genbits_full) begin
              if (cmd_gen_cnt == '0) begin
                cmd_final_ack = 1'b1;
                state_d = Idle;
              end else begin
                // Issue a subsequent gen request.
                state_d = GenArbGnt;
              end
            end
          end else begin
            // Ack for the non-gen request case.
            cmd_final_ack = 1'b1;
            state_d = Idle;
          end
        end
        GenArbGnt: begin
          cmd_arb_req_o = 1'b1;
          if (cmd_arb_gnt_i) begin
            state_d = GenSOP;
          end
        end
        GenSOP: begin
          cmd_arb_sop_o = 1'b1;
          cmd_arb_eop_o = 1'b1;
          cmd_gen_inc_req = 1'b1;
          state_d = GenCmdChk;
          // Check for final genbits beat.
          if (cmd_gen_cnt == GenBitsCntrWidth'(1)) begin
            cmd_gen_cnt_last = 1'b1;
          end
        end
        // Error: The error state is now covered by the if statement above.
        default: begin
          state_d = Error;
          cmd_stage_sm_err_o = 1'b1;
        end
      endcase // unique case (state_q)
    end
  end

  //---------------------------------------------------------
  // Genbits FIFO.
  //---------------------------------------------------------

  prim_fifo_sync #(
    .Width(GenBitsFifoWidth),
    .Pass(0),
    .Depth(GenBitsFifoDepth),
    .OutputZeroIfEmpty(0) // Set to 0, and let last data drive out.
  ) u_prim_fifo_genbits (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!cs_enable_i),
    .wvalid_i       (sfifo_genbits_push),
    .wready_o       (),
    .wdata_i        (sfifo_genbits_wdata),
    .rvalid_o       (sfifo_genbits_not_empty),
    .rready_i       (sfifo_genbits_pop),
    .rdata_o        (sfifo_genbits_rdata),
    .full_o         (sfifo_genbits_full),
    .depth_o        (), // sfifo_genbits_depth)
    .err_o          ()
  );

  assign sfifo_genbits_wdata = {genbits_fips_i,genbits_bus_i};

  assign sfifo_genbits_push = cs_enable_i && genbits_vld_i;

  assign sfifo_genbits_pop = genbits_vld_o && genbits_rdy_i;

  assign genbits_vld_o = cs_enable_i && sfifo_genbits_not_empty;
  assign {genbits_fips_o, genbits_bus_o} = sfifo_genbits_rdata;


  assign sfifo_genbits_err =
         {(sfifo_genbits_push && sfifo_genbits_full),
          (sfifo_genbits_pop && !sfifo_genbits_not_empty),
          (sfifo_genbits_full && !sfifo_genbits_not_empty)};

  //---------------------------------------------------------
  // Ack logic.
  //---------------------------------------------------------

  assign cmd_ack_d =
         (!cs_enable_i) ? '0 :
         cmd_final_ack;

  assign cmd_stage_ack_o = cmd_ack_q;

  assign cmd_ack_sts_d =
         (!cs_enable_i) ? '0 :
         cmd_final_ack ? cmd_ack_sts_i :
         cmd_ack_sts_q;

  assign cmd_stage_ack_sts_o = cmd_ack_sts_q;

  // Make sure that the state machine has a stable error state. This means that after the error
  // state is entered it will not exit it unless a reset signal is received.
  `ASSERT(CsrngCmdStageErrorStStable_A, state_q == Error |=> $stable(state_q))
  // If in error state, the error output must be high.
  `ASSERT(CsrngCmdStageErrorOutput_A,   state_q == Error |-> cmd_stage_sm_err_o)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng block encrypt module
//

module csrng_block_encrypt import csrng_pkg::*; #(
  parameter aes_pkg::sbox_impl_e SBoxImpl = aes_pkg::SBoxImplLut,
  parameter int Cmd = 3,
  parameter int StateId = 4,
  parameter int BlkLen = 128,
  parameter int KeyLen = 256
) (
  input logic                clk_i,
  input logic                rst_ni,

   // update interface
  input logic                block_encrypt_enable_i,
  input logic                block_encrypt_req_i,
  output logic               block_encrypt_rdy_o,
  input logic [KeyLen-1:0]   block_encrypt_key_i,
  input logic [BlkLen-1:0]   block_encrypt_v_i,
  input logic [Cmd-1:0]      block_encrypt_cmd_i,
  input logic [StateId-1:0]  block_encrypt_id_i,
  output logic               block_encrypt_ack_o,
  input logic                block_encrypt_rdy_i,
  output logic [Cmd-1:0]     block_encrypt_cmd_o,
  output logic [StateId-1:0] block_encrypt_id_o,
  output logic [BlkLen-1:0]  block_encrypt_v_o,
  output logic               block_encrypt_quiet_o,
  output logic               block_encrypt_aes_cipher_sm_err_o,
  output logic [2:0]         block_encrypt_sfifo_blkenc_err_o
);

  localparam int BlkEncFifoDepth = 1;
  localparam int BlkEncFifoWidth = StateId+Cmd;
  localparam int NumShares = 1;

  // signals
  // blk_encrypt_in fifo
  logic [BlkEncFifoWidth-1:0] sfifo_blkenc_rdata;
  logic                       sfifo_blkenc_push;
  logic [BlkEncFifoWidth-1:0] sfifo_blkenc_wdata;
  logic                       sfifo_blkenc_pop;
  logic                       sfifo_blkenc_full;
  logic                       sfifo_blkenc_not_empty;
  // breakout
  logic [Cmd-1:0]             sfifo_blkenc_cmd;
  logic [StateId-1:0]         sfifo_blkenc_id;

  aes_pkg::sp2v_e       cipher_in_valid;
  aes_pkg::sp2v_e       cipher_in_ready;
  aes_pkg::sp2v_e       cipher_out_valid;
  aes_pkg::sp2v_e       cipher_out_ready;
  aes_pkg::sp2v_e       cipher_crypt_busy;
  logic [BlkLen-1:0]    cipher_data_out;
  logic                 aes_cipher_core_enable;

  logic [aes_pkg::WidthPRDClearing-1:0] prd_clearing [NumShares];

  logic [3:0][3:0][7:0] state_init[NumShares];

  logic [7:0][31:0]     key_init[NumShares];
  logic [3:0][3:0][7:0] state_done[NumShares];
  logic [3:0][3:0][7:0] state_out;

  assign     prd_clearing[0] = '0;

  assign     state_init[0] = aes_pkg::aes_transpose({<<8{block_encrypt_v_i}});

  assign     key_init[0] = {<<8{block_encrypt_key_i}};
  assign     state_out = aes_pkg::aes_transpose(state_done[0]);
  assign     cipher_data_out = {<<8{state_out}};


  //--------------------------------------------
  // aes cipher core lifecycle enable
  //--------------------------------------------

  assign     aes_cipher_core_enable = block_encrypt_enable_i;

  //--------------------------------------------
  // aes cipher core
  //--------------------------------------------
  assign cipher_in_valid = (aes_cipher_core_enable && block_encrypt_req_i) ?
      aes_pkg::SP2V_HIGH : aes_pkg::SP2V_LOW;

  // SEC_CM: AES_CIPHER.FSM.SPARSE
  // SEC_CM: AES_CIPHER.FSM.REDUN
  // SEC_CM: AES_CIPHER.CTRL.SPARSE
  // SEC_CM: AES_CIPHER.FSM.LOCAL_ESC
  // SEC_CM: AES_CIPHER.CTR.REDUN
  // SEC_CM: AES_CIPHER.DATA_REG.LOCAL_ESC

  aes_cipher_core #(
    .AES192Enable ( 1'b0 ),  // AES192Enable disabled
    .SecMasking   ( 1'b0 ),  // Masking disable
    .SecSBoxImpl  ( SBoxImpl )
  ) u_aes_cipher_core   (
    .clk_i              (clk_i),
    .rst_ni             (rst_ni),

    .cfg_valid_i        ( 1'b1                       ),
    .in_valid_i         ( cipher_in_valid            ),
    .in_ready_o         ( cipher_in_ready            ),
    .out_valid_o        ( cipher_out_valid           ),
    .out_ready_i        ( cipher_out_ready           ),
    .op_i               ( aes_pkg::CIPH_FWD          ),
    .key_len_i          ( aes_pkg::AES_256           ),
    .crypt_i            ( aes_pkg::SP2V_HIGH         ), // Enable
    .crypt_o            ( cipher_crypt_busy          ),
    .alert_fatal_i      ( 1'b0                       ),
    .alert_o            ( block_encrypt_aes_cipher_sm_err_o),
    .dec_key_gen_i      ( aes_pkg::SP2V_LOW          ), // Disable
    .dec_key_gen_o      (                            ),
    .prng_reseed_i      ( 1'b0                       ), // Disable
    .prng_reseed_o      (                            ),
    .key_clear_i        ( 1'b0                       ), // Disable
    .key_clear_o        (                            ),
    .data_out_clear_i   ( 1'b0                       ), // Disable
    .data_out_clear_o   (                            ),
    .prd_clearing_i     ( prd_clearing               ),
    .force_masks_i      ( 1'b0                       ),
    .data_in_mask_o     (                            ),
    .entropy_req_o      (                            ),
    .entropy_ack_i      ( 1'b0                       ),
    .entropy_i          ( '0                         ),

    .state_init_i       ( state_init                 ),
    .key_init_i         ( key_init                   ),
    .state_o            ( state_done                 )
  );


  //--------------------------------------------
  // cmd / id tracking fifo
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(BlkEncFifoWidth),
    .Pass(0),
    .Depth(BlkEncFifoDepth)
  ) u_prim_fifo_sync_blkenc (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!block_encrypt_enable_i),
    .wvalid_i (sfifo_blkenc_push),
    .wready_o (),
    .wdata_i  (sfifo_blkenc_wdata),
    .rvalid_o (sfifo_blkenc_not_empty),
    .rready_i (sfifo_blkenc_pop),
    .rdata_o  (sfifo_blkenc_rdata),
    .full_o   (sfifo_blkenc_full),
    .depth_o  (),
    .err_o    ()
  );

  assign sfifo_blkenc_push = block_encrypt_req_i && !sfifo_blkenc_full;
  assign sfifo_blkenc_wdata = {block_encrypt_id_i,block_encrypt_cmd_i};

  assign block_encrypt_rdy_o = (cipher_in_ready == aes_pkg::SP2V_HIGH);

  assign sfifo_blkenc_pop = block_encrypt_ack_o;
  assign {sfifo_blkenc_id,sfifo_blkenc_cmd} = sfifo_blkenc_rdata;

  assign block_encrypt_ack_o = block_encrypt_rdy_i && (cipher_out_valid == aes_pkg::SP2V_HIGH);

  assign block_encrypt_cmd_o = sfifo_blkenc_cmd;
  assign block_encrypt_id_o = sfifo_blkenc_id;
  assign block_encrypt_v_o = cipher_data_out;

  assign cipher_out_ready = block_encrypt_rdy_i ? aes_pkg::SP2V_HIGH : aes_pkg::SP2V_LOW;

  assign block_encrypt_sfifo_blkenc_err_o =
         {(sfifo_blkenc_push && sfifo_blkenc_full),
          (sfifo_blkenc_pop && !sfifo_blkenc_not_empty),
          (sfifo_blkenc_full && !sfifo_blkenc_not_empty)};

  //--------------------------------------------
  // idle detection
  //--------------------------------------------

  // simple aes cipher activity detector
  assign block_encrypt_quiet_o =
         ((cipher_in_valid == aes_pkg::SP2V_LOW) || (cipher_in_ready == aes_pkg::SP2V_LOW)) &&
         (cipher_crypt_busy == aes_pkg::SP2V_LOW);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng ctr_drbg commands module
//
// Accepts all csrng commands

module csrng_ctr_drbg_cmd import csrng_pkg::*; #(
  parameter int Cmd = 3,
  parameter int StateId = 4,
  parameter int BlkLen = 128,
  parameter int KeyLen = 256,
  parameter int SeedLen = 384,
  parameter int CtrLen  = 32
) (
  input logic                clk_i,
  input logic                rst_ni,

   // command interface
  input logic                ctr_drbg_cmd_enable_i,
  input logic                ctr_drbg_cmd_req_i,
  output logic               ctr_drbg_cmd_rdy_o, // ready to process the req above
  input logic [Cmd-1:0]      ctr_drbg_cmd_ccmd_i,    // current command
  input logic [StateId-1:0]  ctr_drbg_cmd_inst_id_i, // instantance id
  input logic                ctr_drbg_cmd_glast_i,   // gen cmd last beat
  input logic [SeedLen-1:0]  ctr_drbg_cmd_entropy_i, // es entropy
  input logic                ctr_drbg_cmd_entropy_fips_i, // es entropy)fips
  input logic [SeedLen-1:0]  ctr_drbg_cmd_adata_i,   // additional data
  input logic [KeyLen-1:0]   ctr_drbg_cmd_key_i,
  input logic [BlkLen-1:0]   ctr_drbg_cmd_v_i,
  input logic [CtrLen-1:0]   ctr_drbg_cmd_rc_i,
  input logic                ctr_drbg_cmd_fips_i,

  output logic               ctr_drbg_cmd_ack_o, // final ack when update process has been completed
  output logic               ctr_drbg_cmd_sts_o, // final ack status
  input logic                ctr_drbg_cmd_rdy_i, // ready to process the ack above
  output logic [Cmd-1:0]     ctr_drbg_cmd_ccmd_o,
  output logic [StateId-1:0] ctr_drbg_cmd_inst_id_o,
  output logic               ctr_drbg_cmd_glast_o,
  output logic               ctr_drbg_cmd_fips_o,
  output logic [SeedLen-1:0] ctr_drbg_cmd_adata_o,
  output logic [KeyLen-1:0]  ctr_drbg_cmd_key_o,
  output logic [BlkLen-1:0]  ctr_drbg_cmd_v_o,
  output logic [CtrLen-1:0]  ctr_drbg_cmd_rc_o,

   // update interface
  output logic               cmd_upd_req_o,
  input logic                upd_cmd_rdy_i,
  output logic [Cmd-1:0]     cmd_upd_ccmd_o,
  output logic [StateId-1:0] cmd_upd_inst_id_o,
  output logic [SeedLen-1:0] cmd_upd_pdata_o,
  output logic [KeyLen-1:0]  cmd_upd_key_o,
  output logic [BlkLen-1:0]  cmd_upd_v_o,

  input logic                upd_cmd_ack_i,
  output logic               cmd_upd_rdy_o,
  input logic [Cmd-1:0]      upd_cmd_ccmd_i,
  input logic [StateId-1:0]  upd_cmd_inst_id_i,
  input logic [KeyLen-1:0]   upd_cmd_key_i,
  input logic [BlkLen-1:0]   upd_cmd_v_i,
  // misc
  output logic [2:0]         ctr_drbg_cmd_sfifo_cmdreq_err_o,
  output logic [2:0]         ctr_drbg_cmd_sfifo_rcstage_err_o,
  output logic [2:0]         ctr_drbg_cmd_sfifo_keyvrc_err_o
);

  localparam int CmdreqFifoDepth = 1;
  localparam int CmdreqFifoWidth = KeyLen+BlkLen+CtrLen+1+2*SeedLen+1+StateId+Cmd;
  localparam int RCStageFifoDepth = 1;
  localparam int RCStageFifoWidth = KeyLen+BlkLen+StateId+CtrLen+1+SeedLen+1+Cmd;
  localparam int KeyVRCFifoDepth = 1;
  localparam int KeyVRCFifoWidth = KeyLen+BlkLen+CtrLen+1+SeedLen+1+StateId+Cmd;


  // signals
  logic [Cmd-1:0]     cmdreq_ccmd;
  logic [StateId-1:0] cmdreq_id;
  logic               cmdreq_glast;
  logic [SeedLen-1:0] cmdreq_entropy;
  logic               cmdreq_entropy_fips;
  logic [SeedLen-1:0] cmdreq_adata;
  logic [KeyLen-1:0]  cmdreq_key;
  logic [BlkLen-1:0]  cmdreq_v;
  logic [CtrLen-1:0]  cmdreq_rc;

  logic [SeedLen-1:0] prep_seed_material;
  logic [KeyLen-1:0]  prep_key;
  logic [BlkLen-1:0]  prep_v;
  logic [CtrLen-1:0]  prep_rc;
  logic               prep_gen_adata_null;
  logic [KeyLen-1:0]  rcstage_key;
  logic [BlkLen-1:0]  rcstage_v;
  logic [StateId-1:0] rcstage_id;
  logic [CtrLen-1:0]  rcstage_rc;
  logic [Cmd-1:0]     rcstage_ccmd;
  logic               rcstage_glast;
  logic [SeedLen-1:0] rcstage_adata;
  logic               rcstage_fips;
  logic               fips_modified;

  // cmdreq fifo
  logic [CmdreqFifoWidth-1:0] sfifo_cmdreq_rdata;
  logic                       sfifo_cmdreq_push;
  logic [CmdreqFifoWidth-1:0] sfifo_cmdreq_wdata;
  logic                       sfifo_cmdreq_pop;
  logic                       sfifo_cmdreq_full;
  logic                       sfifo_cmdreq_not_empty;

  // rcstage fifo
  logic [RCStageFifoWidth-1:0] sfifo_rcstage_rdata;
  logic                        sfifo_rcstage_push;
  logic [RCStageFifoWidth-1:0] sfifo_rcstage_wdata;
  logic                        sfifo_rcstage_pop;
  logic                        sfifo_rcstage_full;
  logic                        sfifo_rcstage_not_empty;

  // keyvrc fifo
  logic [KeyVRCFifoWidth-1:0]  sfifo_keyvrc_rdata;
  logic                        sfifo_keyvrc_push;
  logic [KeyVRCFifoWidth-1:0]  sfifo_keyvrc_wdata;
  logic                        sfifo_keyvrc_pop;
  logic                        sfifo_keyvrc_full;
  logic                        sfifo_keyvrc_not_empty;

  // flops
  logic                        gen_adata_null_q, gen_adata_null_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      gen_adata_null_q  <= '0;
    end else begin
      gen_adata_null_q  <= gen_adata_null_d;
    end
  end

  //--------------------------------------------
  // input request fifo for staging cmd request
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(CmdreqFifoWidth),
    .Pass(0),
    .Depth(CmdreqFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_cmdreq (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_cmd_enable_i),
    .wvalid_i       (sfifo_cmdreq_push),
    .wready_o       (),
    .wdata_i        (sfifo_cmdreq_wdata),
    .rvalid_o       (sfifo_cmdreq_not_empty),
    .rready_i       (sfifo_cmdreq_pop),
    .rdata_o        (sfifo_cmdreq_rdata),
    .full_o         (sfifo_cmdreq_full),
    .depth_o        (),
    .err_o          ()
  );

  assign fips_modified = ((ctr_drbg_cmd_ccmd_i == INS) ||
                          (ctr_drbg_cmd_ccmd_i == RES)) ? ctr_drbg_cmd_entropy_fips_i :
                         ctr_drbg_cmd_fips_i;

  assign sfifo_cmdreq_wdata = {ctr_drbg_cmd_key_i,ctr_drbg_cmd_v_i,
                               ctr_drbg_cmd_rc_i,fips_modified,
                               ctr_drbg_cmd_entropy_i,ctr_drbg_cmd_adata_i,
                               ctr_drbg_cmd_glast_i,
                               ctr_drbg_cmd_inst_id_i,ctr_drbg_cmd_ccmd_i};

  assign sfifo_cmdreq_push = ctr_drbg_cmd_enable_i && ctr_drbg_cmd_req_i;

  assign sfifo_cmdreq_pop = ctr_drbg_cmd_enable_i &&
         (upd_cmd_rdy_i || gen_adata_null_q) && sfifo_cmdreq_not_empty;

  assign {cmdreq_key,cmdreq_v,cmdreq_rc,
          cmdreq_entropy_fips,cmdreq_entropy,cmdreq_adata,
          cmdreq_glast,cmdreq_id,cmdreq_ccmd} = sfifo_cmdreq_rdata;

  assign ctr_drbg_cmd_rdy_o = !sfifo_cmdreq_full;

  assign ctr_drbg_cmd_sfifo_cmdreq_err_o =
         {(sfifo_cmdreq_push && sfifo_cmdreq_full),
          (sfifo_cmdreq_pop && !sfifo_cmdreq_not_empty),
          (sfifo_cmdreq_full && !sfifo_cmdreq_not_empty)};


  //--------------------------------------------
  // prepare values for update step
  //--------------------------------------------

  assign prep_seed_material =
         (cmdreq_ccmd == INS) ? (cmdreq_entropy ^ cmdreq_adata) :
         (cmdreq_ccmd == RES) ? (cmdreq_entropy ^ cmdreq_adata) :
         (cmdreq_ccmd == GEN) ? cmdreq_adata :
         (cmdreq_ccmd == UPD) ? cmdreq_adata :
         '0;

  assign prep_key =
         (cmdreq_ccmd == INS) ? {KeyLen{1'b0}} :
         (cmdreq_ccmd == RES) ? cmdreq_key :
         (cmdreq_ccmd == GEN) ? cmdreq_key :
         (cmdreq_ccmd == UPD) ? cmdreq_key :
         '0;

  assign prep_v =
         (cmdreq_ccmd == INS) ? {BlkLen{1'b0}} :
         (cmdreq_ccmd == RES) ? cmdreq_v :
         (cmdreq_ccmd == GEN) ? cmdreq_v :
         (cmdreq_ccmd == UPD) ? cmdreq_v :
         '0;

  assign prep_rc =
         (cmdreq_ccmd == INS) ? {{(CtrLen-1){1'b0}},1'b1} :
         (cmdreq_ccmd == RES) ? {{(CtrLen-1){1'b0}},1'b1} :
         (cmdreq_ccmd == GEN) ? cmdreq_rc :
         (cmdreq_ccmd == UPD) ? cmdreq_rc :
         '0;

  assign prep_gen_adata_null = (cmdreq_ccmd == GEN) && (cmdreq_adata == '0);

  assign gen_adata_null_d = ~ctr_drbg_cmd_enable_i ? '0 : prep_gen_adata_null;

  // send to the update block
  assign cmd_upd_req_o = sfifo_cmdreq_not_empty && !prep_gen_adata_null;
  assign cmd_upd_ccmd_o = cmdreq_ccmd;
  assign cmd_upd_inst_id_o = cmdreq_id;
  assign cmd_upd_pdata_o = prep_seed_material;
  assign cmd_upd_key_o = prep_key;
  assign cmd_upd_v_o = prep_v;



  //--------------------------------------------
  // fifo to stage rc and command, waiting for update block to ack
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(RCStageFifoWidth),
    .Pass(0),
    .Depth(RCStageFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_rcstage (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_cmd_enable_i),
    .wvalid_i       (sfifo_rcstage_push),
    .wready_o       (),
    .wdata_i        (sfifo_rcstage_wdata),
    .rvalid_o       (sfifo_rcstage_not_empty),
    .rready_i       (sfifo_rcstage_pop),
    .rdata_o        (sfifo_rcstage_rdata),
    .full_o         (sfifo_rcstage_full),
    .depth_o        (),
    .err_o          ()
  );

  assign sfifo_rcstage_push = sfifo_cmdreq_pop;
  assign sfifo_rcstage_wdata = {prep_key,prep_v,cmdreq_id,prep_rc,cmdreq_entropy_fips,
                                cmdreq_adata,cmdreq_glast,cmdreq_ccmd};
  assign sfifo_rcstage_pop = sfifo_rcstage_not_empty && (upd_cmd_ack_i || gen_adata_null_q);
  assign {rcstage_key,rcstage_v,rcstage_id,rcstage_rc,rcstage_fips,
          rcstage_adata,rcstage_glast,rcstage_ccmd} = sfifo_rcstage_rdata;


  assign ctr_drbg_cmd_sfifo_rcstage_err_o =
         {(sfifo_rcstage_push && sfifo_rcstage_full),
          (sfifo_rcstage_pop && !sfifo_rcstage_not_empty),
          (sfifo_rcstage_full && !sfifo_rcstage_not_empty)};

  assign cmd_upd_rdy_o = sfifo_rcstage_not_empty && !sfifo_keyvrc_full;

  //--------------------------------------------
  // final cmd block processing
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(KeyVRCFifoWidth),
    .Pass(0),
    .Depth(KeyVRCFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_keyvrc (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_cmd_enable_i),
    .wvalid_i       (sfifo_keyvrc_push),
    .wready_o       (),
    .wdata_i        (sfifo_keyvrc_wdata),
    .rvalid_o       (sfifo_keyvrc_not_empty),
    .rready_i       (sfifo_keyvrc_pop),
    .rdata_o        (sfifo_keyvrc_rdata),
    .full_o         (sfifo_keyvrc_full),
    .depth_o        (),
    .err_o          ()
  );

  assign sfifo_keyvrc_push = sfifo_rcstage_pop;

  // if a UNI command, reset the state values
  assign sfifo_keyvrc_wdata = (rcstage_ccmd == UNI) ?
         {{(KeyLen+BlkLen+CtrLen+1+SeedLen){1'b0}},rcstage_glast,upd_cmd_inst_id_i,upd_cmd_ccmd_i} :
         gen_adata_null_q ?
         {rcstage_key,rcstage_v,rcstage_rc,rcstage_fips,
          rcstage_adata,rcstage_glast,rcstage_id,rcstage_ccmd} :
         {upd_cmd_key_i,upd_cmd_v_i,rcstage_rc,rcstage_fips,
          rcstage_adata,rcstage_glast,upd_cmd_inst_id_i,upd_cmd_ccmd_i};

  assign sfifo_keyvrc_pop = ctr_drbg_cmd_rdy_i && sfifo_keyvrc_not_empty;
  assign {ctr_drbg_cmd_key_o,ctr_drbg_cmd_v_o,ctr_drbg_cmd_rc_o,
          ctr_drbg_cmd_fips_o,ctr_drbg_cmd_adata_o,ctr_drbg_cmd_glast_o,
          ctr_drbg_cmd_inst_id_o,ctr_drbg_cmd_ccmd_o} = sfifo_keyvrc_rdata;

  assign ctr_drbg_cmd_sfifo_keyvrc_err_o =
         {(sfifo_keyvrc_push && sfifo_keyvrc_full),
          (sfifo_keyvrc_pop && !sfifo_keyvrc_not_empty),
          (sfifo_keyvrc_full && !sfifo_keyvrc_not_empty)};

  // block ack
  assign ctr_drbg_cmd_ack_o = sfifo_keyvrc_pop;

  assign ctr_drbg_cmd_sts_o = sfifo_keyvrc_pop && (ctr_drbg_cmd_ccmd_o == UNI) &&
         ((KeyLen == '0) && (BlkLen == '0) && (CtrLen == '0));


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng ctr_drbg_update module
//
// implementation using security_strength = 256

module csrng_ctr_drbg_upd #(
  parameter int Cmd = 3,
  parameter int StateId = 4,
  parameter int BlkLen = 128,
  parameter int KeyLen = 256,
  parameter int SeedLen = 384,
  parameter int CtrLen  = 32
) (
  input logic                clk_i,
  input logic                rst_ni,

   // update interface
  input logic                ctr_drbg_upd_enable_i,
  input logic                ctr_drbg_upd_req_i,
  output logic               ctr_drbg_upd_rdy_o, // ready to process the req above
  input logic [Cmd-1:0]      ctr_drbg_upd_ccmd_i,
  input logic [StateId-1:0]  ctr_drbg_upd_inst_id_i, // instantance id
  input logic [SeedLen-1:0]  ctr_drbg_upd_pdata_i, // provided_data
  input logic [KeyLen-1:0]   ctr_drbg_upd_key_i,
  input logic [BlkLen-1:0]   ctr_drbg_upd_v_i,
  output logic [Cmd-1:0]     ctr_drbg_upd_ccmd_o,
  output logic [StateId-1:0] ctr_drbg_upd_inst_id_o,
  output logic [KeyLen-1:0]  ctr_drbg_upd_key_o,
  output logic [BlkLen-1:0]  ctr_drbg_upd_v_o,
  output logic               ctr_drbg_upd_ack_o, // final ack when update process has been completed
  input logic                ctr_drbg_upd_rdy_i, // readu to process the ack above

   // es_req/ack
  input logic                ctr_drbg_upd_es_req_i,
  output logic               ctr_drbg_upd_es_ack_o,

   // block encrypt interface
  output logic               block_encrypt_req_o,
  input logic                block_encrypt_rdy_i,
  output logic [Cmd-1:0]     block_encrypt_ccmd_o,
  output logic [StateId-1:0] block_encrypt_inst_id_o,
  output logic [KeyLen-1:0]  block_encrypt_key_o,
  output logic [BlkLen-1:0]  block_encrypt_v_o,
  input logic                block_encrypt_ack_i,
  output logic               block_encrypt_rdy_o,
  input logic [Cmd-1:0]      block_encrypt_ccmd_i,
  input logic [StateId-1:0]  block_encrypt_inst_id_i,
  input logic [BlkLen-1:0]   block_encrypt_v_i,
  output logic               ctr_drbg_upd_v_ctr_err_o,
  output logic [2:0]         ctr_drbg_upd_sfifo_updreq_err_o,
  output logic [2:0]         ctr_drbg_upd_sfifo_bencreq_err_o,
  output logic [2:0]         ctr_drbg_upd_sfifo_bencack_err_o,
  output logic [2:0]         ctr_drbg_upd_sfifo_pdata_err_o,
  output logic [2:0]         ctr_drbg_upd_sfifo_final_err_o,
  output logic               ctr_drbg_updbe_sm_err_o,
  output logic               ctr_drbg_updob_sm_err_o
);

  localparam int UpdReqFifoDepth = 1;
  localparam int UpdReqFifoWidth = KeyLen+BlkLen+SeedLen+StateId+Cmd;
  localparam int BlkEncReqFifoDepth = 1;
  localparam int BlkEncReqFifoWidth = KeyLen+BlkLen+StateId+Cmd;
  localparam int BlkEncAckFifoDepth = 1;
  localparam int BlkEncAckFifoWidth = BlkLen+StateId+Cmd;
  localparam int PDataFifoDepth = 1;
  localparam int PDataFifoWidth = SeedLen;
  localparam int FinalFifoDepth = 1;
  localparam int FinalFifoWidth = KeyLen+BlkLen+StateId+Cmd;

  // signals
  logic [SeedLen-1:0] updated_key_and_v;
  logic [CtrLen-1:0]  v_inc;
  logic [BlkLen-1:0]  v_first;
  logic [BlkLen-1:0]  v_sized;

  // upd_req fifo
  logic [UpdReqFifoWidth-1:0] sfifo_updreq_rdata;
  logic                       sfifo_updreq_push;
  logic [UpdReqFifoWidth-1:0] sfifo_updreq_wdata;
  logic                       sfifo_updreq_pop;
  logic                       sfifo_updreq_full;
  logic                       sfifo_updreq_not_empty;
  // breakout
  logic [Cmd-1:0]             sfifo_updreq_ccmd;
  logic [StateId-1:0]         sfifo_updreq_inst_id;
  logic [SeedLen-1:0]         sfifo_updreq_pdata;
  logic [KeyLen-1:0]          sfifo_updreq_key;
  logic [BlkLen-1:0]          sfifo_updreq_v;

  // blk_encrypt_req fifo
  logic [BlkEncReqFifoWidth-1:0] sfifo_bencreq_rdata;
  logic                       sfifo_bencreq_push;
  logic [BlkEncReqFifoWidth-1:0] sfifo_bencreq_wdata;
  logic                       sfifo_bencreq_pop;
  logic                       sfifo_bencreq_full;
  logic                       sfifo_bencreq_not_empty;
  // breakout
  logic [Cmd-1:0]             sfifo_bencreq_ccmd;
  logic [StateId-1:0]         sfifo_bencreq_inst_id;
  logic [KeyLen-1:0]          sfifo_bencreq_key;
  logic [BlkLen-1:0]          sfifo_bencreq_v;

  // blk_encrypt_ack fifo
  logic [BlkEncAckFifoWidth-1:0] sfifo_bencack_rdata;
  logic                       sfifo_bencack_push;
  logic [BlkEncAckFifoWidth-1:0] sfifo_bencack_wdata;
  logic                       sfifo_bencack_pop;
  logic                       sfifo_bencack_full;
  logic                       sfifo_bencack_not_empty;
  // breakout
  logic [Cmd-1:0]             sfifo_bencack_ccmd;
  logic [StateId-1:0]         sfifo_bencack_inst_id;
  logic [BlkLen-1:0]          sfifo_bencack_v;

  // pdata_stage fifo
  logic [PDataFifoWidth-1:0]  sfifo_pdata_rdata;
  logic                       sfifo_pdata_push;
  logic [PDataFifoWidth-1:0]  sfifo_pdata_wdata;
  logic                       sfifo_pdata_pop;
  logic                       sfifo_pdata_full;
  logic                       sfifo_pdata_not_empty;
  logic [SeedLen-1:0]         sfifo_pdata_v;

  // key_v fifo
  logic [FinalFifoWidth-1:0]  sfifo_final_rdata;
  logic                       sfifo_final_push;
  logic [FinalFifoWidth-1:0]  sfifo_final_wdata;
  logic                       sfifo_final_pop;
  logic                       sfifo_final_full;
  logic                       sfifo_final_not_empty;
  // breakout
  logic [Cmd-1:0]             sfifo_final_ccmd;
  logic [StateId-1:0]         sfifo_final_inst_id;
  logic [KeyLen-1:0]          sfifo_final_key;
  logic [BlkLen-1:0]          sfifo_final_v;

  logic               v_ctr_load;
  logic               v_ctr_inc;
  logic               interate_ctr_done;
  logic               interate_ctr_inc;
  logic               concat_outblk_shift;
  logic               concat_ctr_done;
  logic               concat_ctr_inc;
  logic [SeedLen+BlkLen-1:0] concat_outblk_shifted_value;
  logic [CtrLen-1:0]         v_ctr;

  // flops
  logic [1:0]         interate_ctr_q, interate_ctr_d;
  logic [1:0]         concat_ctr_q, concat_ctr_d;
  logic [SeedLen-1:0] concat_outblk_q, concat_outblk_d;
  logic [Cmd-1:0]     concat_ccmd_q, concat_ccmd_d;
  logic [StateId-1:0] concat_inst_id_q, concat_inst_id_d;

// Encoding generated with:
// $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 5 \
//      -s 47328894 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (66.67%)
//  4: |||||||||| (33.33%)
//  5: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 4
// Minimum Hamming weight: 2
// Maximum Hamming weight: 3
//

  localparam int BlkEncStateWidth = 5;
  typedef enum logic [BlkEncStateWidth-1:0] {
    ReqIdle = 5'b11000,
    ReqSend = 5'b10011,
    ESHalt  = 5'b01110,
    BEError = 5'b00101
  } blk_enc_state_e;

  blk_enc_state_e blk_enc_state_d, blk_enc_state_q;

  // SEC_CM: BLK_ENC.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_blk_enc_state_regs, blk_enc_state_d,
      blk_enc_state_q, blk_enc_state_e, ReqIdle)

// Encoding generated with:
// $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 6 \
//      -s 400877681 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (66.67%)
//  4: ||||| (16.67%)
//  5: --
//  6: ||||| (16.67%)
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 6
// Minimum Hamming weight: 2
// Maximum Hamming weight: 4
//

  localparam int OutBlkStateWidth = 6;
  typedef enum logic [OutBlkStateWidth-1:0] {
    AckIdle = 6'b110110,
    Load    = 6'b110001,
    Shift   = 6'b001001,
    OBError = 6'b011100
  } outblk_state_e;

  outblk_state_e outblk_state_d, outblk_state_q;

  // SEC_CM: OUTBLK.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_outblk_state_regs, outblk_state_d,
      outblk_state_q, outblk_state_e, AckIdle)

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      interate_ctr_q     <= '0;
      concat_ctr_q       <= '0;
      concat_outblk_q    <= '0;
      concat_ccmd_q      <= '0;
      concat_inst_id_q   <= '0;
    end else begin
      interate_ctr_q     <= interate_ctr_d;
      concat_ctr_q       <= concat_ctr_d;
      concat_outblk_q    <= concat_outblk_d;
      concat_ccmd_q      <= concat_ccmd_d;
      concat_inst_id_q   <= concat_inst_id_d;
    end // else: !if(!rst_ni)


  //--------------------------------------------
  // input request fifo for staging update requests
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(UpdReqFifoWidth),
    .Pass(0),
    .Depth(UpdReqFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_updreq (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!ctr_drbg_upd_enable_i),
    .wvalid_i (sfifo_updreq_push),
    .wready_o (),
    .wdata_i  (sfifo_updreq_wdata),
    .rvalid_o (sfifo_updreq_not_empty),
    .rready_i (sfifo_updreq_pop),
    .rdata_o  (sfifo_updreq_rdata),
    .full_o   (sfifo_updreq_full),
    .depth_o  (),
    .err_o    ()
  );

  assign sfifo_updreq_push = !sfifo_updreq_full && ctr_drbg_upd_req_i;
  assign sfifo_updreq_wdata = {ctr_drbg_upd_key_i,ctr_drbg_upd_v_i,ctr_drbg_upd_pdata_i,
                               ctr_drbg_upd_inst_id_i,ctr_drbg_upd_ccmd_i};
  assign ctr_drbg_upd_rdy_o = !sfifo_updreq_full;

  assign {sfifo_updreq_key,sfifo_updreq_v,sfifo_updreq_pdata,
          sfifo_updreq_inst_id,sfifo_updreq_ccmd} = sfifo_updreq_rdata;

  assign ctr_drbg_upd_sfifo_updreq_err_o =
         {(sfifo_updreq_push && sfifo_updreq_full),
         (sfifo_updreq_pop && !sfifo_updreq_not_empty),
         (sfifo_updreq_full && !sfifo_updreq_not_empty)};

  //--------------------------------------------
  // prepare value for block_encrypt step
  //--------------------------------------------

  if (CtrLen < BlkLen) begin : g_ctrlen_sm
    // for ctr_len < blocklen
    assign v_inc = sfifo_updreq_v[CtrLen-1:0] + 1;
    assign v_first = {sfifo_updreq_v[BlkLen-1:CtrLen],v_inc};
  end else begin : g_ctrlen_lg
    assign v_first = sfifo_updreq_v + 1;
  end

  // SEC_CM: DRBG_UPD.CTR.REDUN
  prim_count #(
    .Width(CtrLen)
  ) u_prim_count_ctr_drbg (
    .clk_i,
    .rst_ni,
    .clr_i(!ctr_drbg_upd_enable_i),
    .set_i(v_ctr_load),
    .set_cnt_i(v_first[CtrLen-1:0]),
    .incr_en_i(v_ctr_inc), // count up
    .decr_en_i(1'b0),
    .step_i(CtrLen'(1)),
    .cnt_o(v_ctr),
    .cnt_next_o(),
    .err_o(ctr_drbg_upd_v_ctr_err_o)
  );

  assign     v_sized = {v_first[BlkLen-1:CtrLen],v_ctr};

  // interation counter
  assign     interate_ctr_d =
             (!ctr_drbg_upd_enable_i) ? '0 :
             interate_ctr_done ? '0 :
             interate_ctr_inc ? (interate_ctr_q + 1) :
             interate_ctr_q;

  assign interate_ctr_done = (int'(interate_ctr_q) >= SeedLen/BlkLen);

  //--------------------------------------------
  // state machine to send values to block_encrypt
  //--------------------------------------------

  always_comb begin
    blk_enc_state_d = blk_enc_state_q;
    v_ctr_load = 1'b0;
    v_ctr_inc  = 1'b0;
    interate_ctr_inc  = 1'b0;
    sfifo_pdata_push = 1'b0;
    sfifo_bencreq_push = 1'b0;
    sfifo_updreq_pop = 1'b0;
    ctr_drbg_updbe_sm_err_o = 1'b0;
    ctr_drbg_upd_es_ack_o = 1'b0;
    unique case (blk_enc_state_q)
      // ReqIdle: increment v this cycle, push in next
      ReqIdle: begin
        // Prioritize halt requests from entropy_src over disable, as CSRNG would otherwise starve
        // those requests while it is idle.
        if (ctr_drbg_upd_es_req_i) begin
          blk_enc_state_d = ESHalt;
        end else if (!ctr_drbg_upd_enable_i) begin
          blk_enc_state_d = ReqIdle;
        end else if (sfifo_updreq_not_empty && !sfifo_bencreq_full && !sfifo_pdata_full) begin
          v_ctr_load = 1'b1;
          sfifo_pdata_push = 1'b1;
          blk_enc_state_d = ReqSend;
        end
      end
      ReqSend: begin
        if (!ctr_drbg_upd_enable_i) begin
          blk_enc_state_d = ReqIdle;
        end else if (!interate_ctr_done) begin
          if (!sfifo_bencreq_full) begin
            v_ctr_inc  = 1'b1;
            interate_ctr_inc  = 1'b1;
            sfifo_bencreq_push = 1'b1;
          end
        end else begin
          sfifo_updreq_pop = 1'b1;
          blk_enc_state_d = ReqIdle;
        end
      end
      ESHalt: begin
        ctr_drbg_upd_es_ack_o = 1'b1;
        if (!ctr_drbg_upd_es_req_i) begin
          blk_enc_state_d = ReqIdle;
        end
      end
      BEError: begin
        ctr_drbg_updbe_sm_err_o = 1'b1;
      end
      default: begin
        blk_enc_state_d = BEError;
        ctr_drbg_updbe_sm_err_o = 1'b1;
      end
    endcase // case (blk_enc_state_q)
  end

  //--------------------------------------------
  // block_encrypt request fifo for staging aes requests
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(BlkEncReqFifoWidth),
    .Pass(0),
    .Depth(BlkEncReqFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_bencreq (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!ctr_drbg_upd_enable_i),
    .wvalid_i (sfifo_bencreq_push),
    .wready_o (),
    .wdata_i  (sfifo_bencreq_wdata),
    .rvalid_o (sfifo_bencreq_not_empty),
    .rready_i (sfifo_bencreq_pop),
    .rdata_o  (sfifo_bencreq_rdata),
    .full_o   (sfifo_bencreq_full),
    .depth_o  (),
    .err_o    ()
  );

  assign sfifo_bencreq_pop = block_encrypt_req_o && block_encrypt_rdy_i;
  assign block_encrypt_req_o = sfifo_bencreq_not_empty;

  assign sfifo_bencreq_wdata = {sfifo_updreq_key,v_sized,sfifo_updreq_inst_id,sfifo_updreq_ccmd};

  assign {sfifo_bencreq_key,sfifo_bencreq_v,sfifo_bencreq_inst_id,
          sfifo_bencreq_ccmd} = sfifo_bencreq_rdata;

  // set outputs
  assign block_encrypt_key_o = sfifo_bencreq_key;
  assign block_encrypt_v_o = sfifo_bencreq_v;
  assign block_encrypt_inst_id_o = sfifo_bencreq_inst_id;
  assign block_encrypt_ccmd_o = sfifo_bencreq_ccmd;

  assign ctr_drbg_upd_sfifo_bencreq_err_o =
         {(sfifo_bencreq_push && sfifo_bencreq_full),
          (sfifo_bencreq_pop && !sfifo_bencreq_not_empty),
          (sfifo_bencreq_full && !sfifo_bencreq_not_empty)};

  //--------------------------------------------
  // block_encrypt response fifo from block encrypt
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(BlkEncAckFifoWidth),
    .Pass(0),
    .Depth(BlkEncAckFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_bencack (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!ctr_drbg_upd_enable_i),
    .wvalid_i (sfifo_bencack_push),
    .wready_o (),
    .wdata_i  (sfifo_bencack_wdata),
    .rvalid_o (sfifo_bencack_not_empty),
    .rready_i (sfifo_bencack_pop),
    .rdata_o  (sfifo_bencack_rdata),
    .full_o   (sfifo_bencack_full),
    .depth_o  (),
    .err_o    ()
  );

  assign sfifo_bencack_push = !sfifo_bencack_full && block_encrypt_ack_i;
  assign sfifo_bencack_wdata = {block_encrypt_v_i,block_encrypt_inst_id_i,block_encrypt_ccmd_i};
  assign block_encrypt_rdy_o = !sfifo_bencack_full;

  assign {sfifo_bencack_v,sfifo_bencack_inst_id,sfifo_bencack_ccmd} = sfifo_bencack_rdata;

  assign ctr_drbg_upd_sfifo_bencack_err_o =
         {(sfifo_bencack_push && sfifo_bencack_full),
          (sfifo_bencack_pop && !sfifo_bencack_not_empty),
          (sfifo_bencack_full && !sfifo_bencack_not_empty)};

  //--------------------------------------------
  // fifo to stage provided_data, waiting for blk_encrypt to ack
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(PDataFifoWidth),
    .Pass(0),
    .Depth(PDataFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_pdata (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!ctr_drbg_upd_enable_i),
    .wvalid_i (sfifo_pdata_push),
    .wready_o (),
    .wdata_i  (sfifo_pdata_wdata),
    .rvalid_o (sfifo_pdata_not_empty),
    .rready_i (sfifo_pdata_pop),
    .rdata_o  (sfifo_pdata_rdata),
    .full_o   (sfifo_pdata_full),
    .depth_o  (),
    .err_o    ()
  );

  assign sfifo_pdata_wdata = sfifo_updreq_pdata;

  assign sfifo_pdata_v = sfifo_pdata_rdata;

  assign ctr_drbg_upd_sfifo_pdata_err_o =
         {(sfifo_pdata_push && sfifo_pdata_full),
          (sfifo_pdata_pop && !sfifo_pdata_not_empty),
          (sfifo_pdata_full && !sfifo_pdata_not_empty)};

  //--------------------------------------------
  // shifting logic to receive values from block_encrypt
  //--------------------------------------------

  assign concat_outblk_shifted_value = {concat_outblk_q, {BlkLen{1'b0}}};

  assign concat_outblk_d =
         (!ctr_drbg_upd_enable_i) ? '0 :
         sfifo_bencack_pop ? {concat_outblk_q[SeedLen-1:BlkLen],sfifo_bencack_v} :
         concat_outblk_shift ? concat_outblk_shifted_value[SeedLen-1:0] :
         concat_outblk_q;

  // The following signal is used to avoid possible lint errors.
  logic [BlkLen-1:0] unused_concat_outblk_shifted_value;
  assign unused_concat_outblk_shifted_value = concat_outblk_shifted_value[SeedLen+BlkLen-1:SeedLen];

  // concatination counter
  assign concat_ctr_d =
         (!ctr_drbg_upd_enable_i) ? '0 :
         concat_ctr_done ? '0 :
         concat_ctr_inc ? (concat_ctr_q + 1) :
         concat_ctr_q;

  assign concat_ctr_done = (int'(concat_ctr_q) >= (SeedLen/BlkLen));

  assign concat_inst_id_d =
         (!ctr_drbg_upd_enable_i) ? '0 :
         sfifo_bencack_pop ? sfifo_bencack_inst_id :
         concat_inst_id_q;

  assign concat_ccmd_d =
         (!ctr_drbg_upd_enable_i) ? '0 :
         sfifo_bencack_pop ? sfifo_bencack_ccmd :
         concat_ccmd_q;

  //--------------------------------------------
  // state machine to receive values from block_encrypt
  //--------------------------------------------

  always_comb begin
    outblk_state_d = outblk_state_q;
    concat_ctr_inc  = 1'b0;
    concat_outblk_shift = 1'b0;
    sfifo_pdata_pop = 1'b0;
    sfifo_bencack_pop = 1'b0;
    sfifo_final_push = 1'b0;
    ctr_drbg_updob_sm_err_o = 1'b0;
    unique case (outblk_state_q)
      // AckIdle: increment v this cycle, push in next
      AckIdle: begin
        if (!ctr_drbg_upd_enable_i) begin
          outblk_state_d = AckIdle;
        end else if (sfifo_bencack_not_empty && sfifo_pdata_not_empty && !sfifo_final_full) begin
          outblk_state_d = Load;
        end
      end
      Load: begin
        if (!ctr_drbg_upd_enable_i) begin
          outblk_state_d = AckIdle;
        end else if (sfifo_bencack_not_empty) begin
          concat_ctr_inc  = 1'b1;
          sfifo_bencack_pop = 1'b1;
          outblk_state_d = Shift;
        end
      end
      Shift: begin
        if (!ctr_drbg_upd_enable_i) begin
          outblk_state_d = AckIdle;
        end else if (concat_ctr_done) begin
          sfifo_pdata_pop = 1'b1;
          sfifo_final_push = 1'b1;
          outblk_state_d = AckIdle;
        end else begin
          concat_outblk_shift = 1'b1;
          outblk_state_d = Load;
        end
      end
      OBError: begin
        ctr_drbg_updob_sm_err_o = 1'b1;
      end
      default: begin
        outblk_state_d = OBError;
        ctr_drbg_updob_sm_err_o = 1'b1;
      end
    endcase
  end


  //--------------------------------------------
  // final update processing
  //--------------------------------------------

  // XOR the additional data with the new key and value from block encryption
  assign updated_key_and_v = concat_outblk_q ^ sfifo_pdata_v;

  prim_fifo_sync #(
    .Width(FinalFifoWidth),
    .Pass(0),
    .Depth(FinalFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_final (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!ctr_drbg_upd_enable_i),
    .wvalid_i (sfifo_final_push),
    .wready_o (),
    .wdata_i  (sfifo_final_wdata),
    .rvalid_o (sfifo_final_not_empty),
    .rready_i (sfifo_final_pop),
    .rdata_o  (sfifo_final_rdata),
    .full_o   (sfifo_final_full),
    .depth_o  (),
    .err_o    ()
  );

  assign sfifo_final_wdata = {updated_key_and_v,concat_inst_id_q,concat_ccmd_q};

  assign {sfifo_final_key,sfifo_final_v,sfifo_final_inst_id,sfifo_final_ccmd} = sfifo_final_rdata;

  assign sfifo_final_pop = ctr_drbg_upd_rdy_i && sfifo_final_not_empty;
  assign ctr_drbg_upd_ack_o = sfifo_final_pop;
  assign ctr_drbg_upd_ccmd_o = sfifo_final_ccmd;
  assign ctr_drbg_upd_inst_id_o = sfifo_final_inst_id;
  assign ctr_drbg_upd_key_o = sfifo_final_key;
  assign ctr_drbg_upd_v_o = sfifo_final_v;

  assign ctr_drbg_upd_sfifo_final_err_o =
         {(sfifo_final_push && sfifo_final_full),
          (sfifo_final_pop && !sfifo_final_not_empty),
          (sfifo_final_full && !sfifo_final_not_empty)};

  // Make sure that the two state machines have a stable error state. This means that after the
  // error state is entered it will not exit it unless a reset signal is received.
  `ASSERT(CsrngDrbgUpdBlkEncErrorStStable_A,
          blk_enc_state_q == BEError |=> $stable(blk_enc_state_q))
  `ASSERT(CsrngDrbgUpdOutBlkErrorStStable_A,
          outblk_state_q  == OBError |=> $stable(outblk_state_q))
  // If in error state, the error output must be high.
  `ASSERT(CsrngDrbgUpdBlkEncErrorOutput_A, blk_enc_state_q == BEError |-> ctr_drbg_updbe_sm_err_o)
  `ASSERT(CsrngDrbgUpdOutBlkErrorOutput_A, outblk_state_q  == OBError |-> ctr_drbg_updob_sm_err_o)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng ctr_drbg generate module
//
// This module will process the second half of the generate function.
// It takes in the key, v, and reseed counter values processed by the
// ctr_drbg cmd module.

module csrng_ctr_drbg_gen import csrng_pkg::*; #(
  parameter int NApps = 4,
  parameter int Cmd = 3,
  parameter int StateId = 4,
  parameter int BlkLen = 128,
  parameter int KeyLen = 256,
  parameter int SeedLen = 384,
  parameter int CtrLen  = 32
) (
  input logic                clk_i,
  input logic                rst_ni,

   // command interface
  input logic                ctr_drbg_gen_enable_i,
  input logic                ctr_drbg_gen_req_i,
  output logic               ctr_drbg_gen_rdy_o, // ready to process the req above
  input logic [Cmd-1:0]      ctr_drbg_gen_ccmd_i,    // current command
  input logic [StateId-1:0]  ctr_drbg_gen_inst_id_i, // instantance id
  input logic                ctr_drbg_gen_glast_i,   // gen cmd last beat
  input logic                ctr_drbg_gen_fips_i,    // fips
  input logic [SeedLen-1:0]  ctr_drbg_gen_adata_i,   // additional data
  input logic [KeyLen-1:0]   ctr_drbg_gen_key_i,
  input logic [BlkLen-1:0]   ctr_drbg_gen_v_i,
  input logic [CtrLen-1:0]   ctr_drbg_gen_rc_i,

  output logic               ctr_drbg_gen_ack_o, // final ack when update process has been completed
  output logic               ctr_drbg_gen_sts_o, // final ack status
  input logic                ctr_drbg_gen_rdy_i, // ready to process the ack above
  output logic [Cmd-1:0]     ctr_drbg_gen_ccmd_o,
  output logic [StateId-1:0] ctr_drbg_gen_inst_id_o,
  output logic [KeyLen-1:0]  ctr_drbg_gen_key_o,
  output logic [BlkLen-1:0]  ctr_drbg_gen_v_o,
  output logic [CtrLen-1:0]  ctr_drbg_gen_rc_o,
  output logic [BlkLen-1:0]  ctr_drbg_gen_bits_o,
  output logic               ctr_drbg_gen_fips_o,

   // es_req/ack
  input logic                ctr_drbg_gen_es_req_i,
  output logic               ctr_drbg_gen_es_ack_o,

  // update interface
  output logic               gen_upd_req_o,
  input logic                upd_gen_rdy_i,
  output logic [Cmd-1:0]     gen_upd_ccmd_o,
  output logic [StateId-1:0] gen_upd_inst_id_o,
  output logic [SeedLen-1:0] gen_upd_pdata_o,
  output logic [KeyLen-1:0]  gen_upd_key_o,
  output logic [BlkLen-1:0]  gen_upd_v_o,

  input logic                upd_gen_ack_i,
  output logic               gen_upd_rdy_o,
  input logic [Cmd-1:0]      upd_gen_ccmd_i,
  input logic [StateId-1:0]  upd_gen_inst_id_i,
  input logic [KeyLen-1:0]   upd_gen_key_i,
  input logic [BlkLen-1:0]   upd_gen_v_i,
  // block encrypt interface
  output logic               block_encrypt_req_o,
  input logic                block_encrypt_rdy_i,
  output logic [Cmd-1:0]     block_encrypt_ccmd_o,
  output logic [StateId-1:0] block_encrypt_inst_id_o,
  output logic [KeyLen-1:0]  block_encrypt_key_o,
  output logic [BlkLen-1:0]  block_encrypt_v_o,
  input logic                block_encrypt_ack_i,
  output logic               block_encrypt_rdy_o,
  input logic [Cmd-1:0]      block_encrypt_ccmd_i,
  input logic [StateId-1:0]  block_encrypt_inst_id_i,
  input logic [BlkLen-1:0]   block_encrypt_v_i,
  // misc
  output logic               ctr_drbg_gen_v_ctr_err_o,
  output logic [2:0]         ctr_drbg_gen_sfifo_gbencack_err_o,
  output logic [2:0]         ctr_drbg_gen_sfifo_grcstage_err_o,
  output logic [2:0]         ctr_drbg_gen_sfifo_ggenreq_err_o,
  output logic [2:0]         ctr_drbg_gen_sfifo_gadstage_err_o,
  output logic [2:0]         ctr_drbg_gen_sfifo_ggenbits_err_o,
  output logic               ctr_drbg_gen_sm_err_o
);

  localparam int GenreqFifoDepth = 1;
  localparam int GenreqFifoWidth = KeyLen+BlkLen+CtrLen+1+SeedLen+1+StateId+Cmd;
  localparam int BlkEncAckFifoDepth = 1;
  localparam int BlkEncAckFifoWidth = BlkLen+StateId+Cmd;
  localparam int AdstageFifoDepth = 1;
  localparam int AdstageFifoWidth = KeyLen+BlkLen+CtrLen+1+1;
  localparam int RCStageFifoDepth = 1;
  localparam int RCStageFifoWidth = KeyLen+BlkLen+BlkLen+CtrLen+1+1+StateId+Cmd;
  localparam int GenbitsFifoDepth = 1;
  localparam int GenbitsFifoWidth = 1+BlkLen+KeyLen+BlkLen+CtrLen+StateId+Cmd;

  // signals
  logic [Cmd-1:0]     genreq_ccmd;
  logic [StateId-1:0] genreq_id;
  logic               genreq_glast;
  logic [SeedLen-1:0] genreq_adata;
  logic               genreq_fips;
  logic [KeyLen-1:0]  genreq_key;
  logic [BlkLen-1:0]  genreq_v;
  logic [CtrLen-1:0]  genreq_rc;

  logic [KeyLen-1:0]  adstage_key;
  logic [BlkLen-1:0]  adstage_v;
  logic [CtrLen-1:0]  adstage_rc;
  logic               adstage_fips;
  logic               adstage_glast;
  logic [SeedLen-1:0] adstage_adata;

  logic [KeyLen-1:0]  rcstage_key;
  logic [BlkLen-1:0]  rcstage_v;
  logic [BlkLen-1:0]  rcstage_bits;
  logic [CtrLen-1:0]  rcstage_rc;
  logic               rcstage_glast;
  logic               rcstage_fips;
  logic [CtrLen-1:0]  rcstage_rc_plus1;
  logic [Cmd-1:0]     rcstage_ccmd;
  logic [StateId-1:0] rcstage_inst_id;

  logic [Cmd-1:0]     genreq_ccmd_modified;
  logic [Cmd-1:0]     bencack_ccmd_modified;

  // cmdreq fifo
  // logic [$clog2(CmdreqFifoDepth):0] sfifo_cmdreq_depth;
  logic [GenreqFifoWidth-1:0] sfifo_genreq_rdata;
  logic                       sfifo_genreq_push;
  logic [GenreqFifoWidth-1:0] sfifo_genreq_wdata;
  logic                       sfifo_genreq_pop;
  logic                       sfifo_genreq_full;
  logic                       sfifo_genreq_not_empty;

  // adstage fifo
  logic [AdstageFifoWidth-1:0] sfifo_adstage_rdata;
  logic                        sfifo_adstage_push;
  logic [AdstageFifoWidth-1:0] sfifo_adstage_wdata;
  logic                        sfifo_adstage_pop;
  logic                        sfifo_adstage_full;
  logic                        sfifo_adstage_not_empty;
  // blk_encrypt_ack fifo
  logic [BlkEncAckFifoWidth-1:0] sfifo_bencack_rdata;
  logic                       sfifo_bencack_push;
  logic [BlkEncAckFifoWidth-1:0] sfifo_bencack_wdata;
  logic                       sfifo_bencack_pop;
  logic                       sfifo_bencack_full;
  logic                       sfifo_bencack_not_empty;
  // breakout
  logic [Cmd-1:0]             sfifo_bencack_ccmd;
  logic [StateId-1:0]         sfifo_bencack_inst_id;
  logic [BlkLen-1:0]          sfifo_bencack_bits;

  // rcstage fifo
  logic [RCStageFifoWidth-1:0] sfifo_rcstage_rdata;
  logic                        sfifo_rcstage_push;
  logic [RCStageFifoWidth-1:0] sfifo_rcstage_wdata;
  logic                        sfifo_rcstage_pop;
  logic                        sfifo_rcstage_full;
  logic                        sfifo_rcstage_not_empty;

  // genbits fifo
  logic [GenbitsFifoWidth-1:0] sfifo_genbits_rdata;
  logic                        sfifo_genbits_push;
  logic [GenbitsFifoWidth-1:0] sfifo_genbits_wdata;
  logic                        sfifo_genbits_pop;
  logic                        sfifo_genbits_full;
  logic                        sfifo_genbits_not_empty;

  logic [CtrLen-1:0]           v_inc;
  logic [BlkLen-1:0]           v_first;
  logic [BlkLen-1:0]           v_sized;
  logic                        v_ctr_load;
  logic                        v_ctr_inc;
  logic                        interate_ctr_done;
  logic                        interate_ctr_inc;
  logic [NApps-1:0]            capt_adata;
  logic [SeedLen-1:0]          update_adata[NApps];
  logic [CtrLen-1:0]           v_ctr;

  // flops
  logic [1:0]                  interate_ctr_q, interate_ctr_d;
  logic [SeedLen-1:0]          update_adata_q[NApps], update_adata_d[NApps];
  logic [NApps-1:0]            update_adata_vld_q, update_adata_vld_d;

// Encoding generated with:
// $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 5 \
//      -s 2651202796 --language=sv
//
// Hamming distance histogram:
//
//  0: --
//  1: --
//  2: --
//  3: |||||||||||||||||||| (66.67%)
//  4: |||||||||| (33.33%)
//  5: --
//
// Minimum Hamming distance: 3
// Maximum Hamming distance: 4
// Minimum Hamming weight: 2
// Maximum Hamming weight: 3
//

  localparam int StateWidth = 5;
  typedef enum logic [StateWidth-1:0] {
    ReqIdle  = 5'b01101,
    ReqSend  = 5'b00011,
    ESHalt   = 5'b11000,
    ReqError = 5'b10110
} state_e;

  state_e state_d, state_q;

  // SEC_CM: UPDATE.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, ReqIdle)

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      interate_ctr_q     <= '0;
      update_adata_q     <= '{default:0};
      update_adata_vld_q <= '{default:0};
    end else begin
      interate_ctr_q     <= interate_ctr_d;
      update_adata_q     <= update_adata_d;
      update_adata_vld_q <= update_adata_vld_d;
    end



  //--------------------------------------------
  // input request fifo for staging gen request
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(GenreqFifoWidth),
    .Pass(0),
    .Depth(GenreqFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_genreq (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_gen_enable_i),
    .wvalid_i       (sfifo_genreq_push),
    .wready_o       (),
    .wdata_i        (sfifo_genreq_wdata),
    .rvalid_o       (sfifo_genreq_not_empty),
    .rready_i       (sfifo_genreq_pop),
    .rdata_o        (sfifo_genreq_rdata),
    .full_o         (sfifo_genreq_full),
    .depth_o        (),
    .err_o          ()
  );

  assign genreq_ccmd_modified = (ctr_drbg_gen_ccmd_i == GEN) ? GENB : INV;

  assign sfifo_genreq_wdata = {ctr_drbg_gen_key_i,ctr_drbg_gen_v_i,ctr_drbg_gen_rc_i,
                               ctr_drbg_gen_fips_i,ctr_drbg_gen_adata_i,ctr_drbg_gen_glast_i,
                               ctr_drbg_gen_inst_id_i,genreq_ccmd_modified};

  assign sfifo_genreq_push = ctr_drbg_gen_enable_i && ctr_drbg_gen_req_i;

  assign {genreq_key,genreq_v,genreq_rc,
          genreq_fips,genreq_adata,genreq_glast,
          genreq_id,genreq_ccmd} = sfifo_genreq_rdata;

  assign ctr_drbg_gen_rdy_o = !sfifo_genreq_full;

  assign ctr_drbg_gen_sfifo_ggenreq_err_o =
         {(sfifo_genreq_push && sfifo_genreq_full),
          (sfifo_genreq_pop && !sfifo_genreq_not_empty),
          (sfifo_genreq_full && !sfifo_genreq_not_empty)};



  //--------------------------------------------
  // prepare value for block_encrypt step
  //--------------------------------------------

  if (CtrLen < BlkLen) begin : gen_ctrlen_sm
    // for ctr_len < blocklen
    assign v_inc = genreq_v[CtrLen-1:0] + 1;
    assign v_first = {genreq_v[BlkLen-1:CtrLen],v_inc};
  end else begin : g_ctrlen_lg
    assign v_first = genreq_v + 1;
  end

  // SEC_CM: DRBG_GEN.CTR.REDUN
  prim_count #(
    .Width(CtrLen)
  ) u_prim_count_ctr_drbg (
    .clk_i,
    .rst_ni,
    .clr_i(!ctr_drbg_gen_enable_i),
    .set_i(v_ctr_load),
    .set_cnt_i(v_first[CtrLen-1:0]),
    .incr_en_i(v_ctr_inc), // count up
    .decr_en_i(1'b0),
    .step_i(CtrLen'(1)),
    .cnt_o(v_ctr),
    .cnt_next_o(),
    .err_o(ctr_drbg_gen_v_ctr_err_o)
  );

  assign v_sized = {v_first[BlkLen-1:CtrLen],v_ctr};

  // interation counter
  assign interate_ctr_d =
         (!ctr_drbg_gen_enable_i) ? '0 :
         interate_ctr_done ? '0 :
         interate_ctr_inc ? (interate_ctr_q + 1) :
         interate_ctr_q;

  // Supporting only 128b requests
  assign interate_ctr_done = (interate_ctr_q >= 2'(BlkLen/BlkLen));

  //--------------------------------------------
  // state machine to send values to block_encrypt
  //--------------------------------------------

  assign block_encrypt_ccmd_o = genreq_ccmd;
  assign block_encrypt_inst_id_o = genreq_id;
  assign block_encrypt_key_o = genreq_key;
  assign block_encrypt_v_o = v_sized;

  always_comb begin
    state_d = state_q;
    v_ctr_load = 1'b0;
    v_ctr_inc  = 1'b0;
    interate_ctr_inc  = 1'b0;
    sfifo_adstage_push = 1'b0;
    block_encrypt_req_o = 1'b0;
    sfifo_genreq_pop = 1'b0;
    ctr_drbg_gen_sm_err_o = 1'b0;
    ctr_drbg_gen_es_ack_o = 1'b0;
    unique case (state_q)
      // ReqIdle: increment v this cycle, push in next
      ReqIdle: begin
        // Prioritize halt requests from entropy_src over disable, as CSRNG would otherwise starve
        // those requests while it is idle.
        if (ctr_drbg_gen_es_req_i) begin
          state_d = ESHalt;
        end else if (!ctr_drbg_gen_enable_i) begin
          state_d = ReqIdle;
        end else if (sfifo_genreq_not_empty && !sfifo_adstage_full) begin
          v_ctr_load = 1'b1;
          state_d = ReqSend;
        end
      end
      ReqSend: begin
        if (!ctr_drbg_gen_enable_i) begin
          state_d = ReqIdle;
        end else if (!interate_ctr_done) begin
          block_encrypt_req_o = 1'b1;
          sfifo_adstage_push = 1'b1;
          if (block_encrypt_rdy_i) begin
            v_ctr_inc  = 1'b1;
            interate_ctr_inc  = 1'b1;
          end
        end else begin
          sfifo_genreq_pop = 1'b1;
          state_d = ReqIdle;
        end
      end
      ESHalt: begin
        ctr_drbg_gen_es_ack_o = 1'b1;
        if (!ctr_drbg_gen_es_req_i) begin
          state_d = ReqIdle;
        end
      end
      ReqError: begin
        ctr_drbg_gen_sm_err_o = 1'b1;
      end
      default: begin
        state_d = ReqError;
        ctr_drbg_gen_sm_err_o = 1'b1;
      end
    endcase
  end


  //--------------------------------------------
  // fifo to stage key, v, rc, and adata, waiting for update block to ack
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(AdstageFifoWidth),
    .Pass(0),
    .Depth(AdstageFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_adstage (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_gen_enable_i),
    .wvalid_i       (sfifo_adstage_push),
    .wready_o       (),
    .wdata_i        (sfifo_adstage_wdata),
    .rvalid_o       (sfifo_adstage_not_empty),
    .rready_i       (sfifo_adstage_pop),
    .rdata_o        (sfifo_adstage_rdata),
    .full_o         (sfifo_adstage_full),
    .depth_o        (),
    .err_o          ()
  );

  assign sfifo_adstage_wdata = {genreq_key,v_sized,genreq_rc,genreq_fips,genreq_glast};
  assign sfifo_adstage_pop = sfifo_adstage_not_empty && sfifo_bencack_pop;
  assign {adstage_key,adstage_v,adstage_rc,adstage_fips,adstage_glast} = sfifo_adstage_rdata;

  assign ctr_drbg_gen_sfifo_gadstage_err_o =
         {(sfifo_adstage_push && sfifo_adstage_full),
          (sfifo_adstage_pop && !sfifo_adstage_not_empty),
          (sfifo_adstage_full && !sfifo_adstage_not_empty)};


  // array to hold each channel's adata
  for (genvar i = 0; i < NApps; i = i+1) begin : gen_adata
    assign capt_adata[i] = (sfifo_adstage_push && (genreq_id == i));

    assign update_adata_vld_d[i] = ~ctr_drbg_gen_enable_i ? 1'b0 :
           capt_adata[i] && !update_adata_vld_q[i] ? 1'b1 :
           (gen_upd_req_o && upd_gen_rdy_i && (sfifo_bencack_inst_id == i)) ? 1'b0 :
           update_adata_vld_q[i];

    assign update_adata_d[i] = ~ctr_drbg_gen_enable_i ? '0 :
                               (capt_adata[i] && !update_adata_vld_q[i]) ? genreq_adata :
                               update_adata_q[i];
    assign update_adata[i] = update_adata_q[i] & {SeedLen{update_adata_vld_q[i] &&
                                                          (genreq_id == i)}};
  end

  always_comb begin
    adstage_adata = '0;
    for (int i = 0; i < NApps; i = i+1) begin
      // since only one bus is active at a time based on the instant id,
      // an "or" of all the buses can be done below
      adstage_adata |= update_adata[i];
    end
  end


  //--------------------------------------------
  // block_encrypt response fifo from block encrypt
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(BlkEncAckFifoWidth),
    .Pass(0),
    .Depth(BlkEncAckFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_bencack (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!ctr_drbg_gen_enable_i),
    .wvalid_i (sfifo_bencack_push),
    .wready_o (),
    .wdata_i  (sfifo_bencack_wdata),
    .rvalid_o (sfifo_bencack_not_empty),
    .rready_i (sfifo_bencack_pop),
    .rdata_o  (sfifo_bencack_rdata),
    .full_o   (sfifo_bencack_full),
    .depth_o  (),
    .err_o    ()
  );

  assign bencack_ccmd_modified = (block_encrypt_ccmd_i == GENB) ? GENU : INV;

  assign sfifo_bencack_push = !sfifo_bencack_full && block_encrypt_ack_i;
  assign sfifo_bencack_wdata = {block_encrypt_v_i,block_encrypt_inst_id_i,bencack_ccmd_modified};
  assign block_encrypt_rdy_o = !sfifo_bencack_full;

  assign sfifo_bencack_pop = !sfifo_rcstage_full && sfifo_bencack_not_empty &&
                             (upd_gen_rdy_i || !adstage_glast);

  assign {sfifo_bencack_bits,sfifo_bencack_inst_id,sfifo_bencack_ccmd} = sfifo_bencack_rdata;

  assign ctr_drbg_gen_sfifo_gbencack_err_o =
         {(sfifo_bencack_push && sfifo_bencack_full),
          (sfifo_bencack_pop && !sfifo_bencack_not_empty),
          (sfifo_bencack_full && !sfifo_bencack_not_empty)};


  //--------------------------------------------
  // prepare values for update step
  //--------------------------------------------

  // send to the update block
  assign gen_upd_req_o = sfifo_bencack_not_empty && adstage_glast;
  assign gen_upd_ccmd_o = sfifo_bencack_ccmd;
  assign gen_upd_inst_id_o = sfifo_bencack_inst_id;
  assign gen_upd_pdata_o = adstage_adata;
  assign gen_upd_key_o = adstage_key;
  assign gen_upd_v_o = adstage_v;



  //--------------------------------------------
  // fifo to stage rc, waiting for update block to ack
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(RCStageFifoWidth),
    .Pass(0),
    .Depth(RCStageFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_rcstage (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_gen_enable_i),
    .wvalid_i       (sfifo_rcstage_push),
    .wready_o       (),
    .wdata_i        (sfifo_rcstage_wdata),
    .rvalid_o       (sfifo_rcstage_not_empty),
    .rready_i       (sfifo_rcstage_pop),
    .rdata_o        (sfifo_rcstage_rdata),
    .full_o         (sfifo_rcstage_full),
    .depth_o        (),
    .err_o          ()
  );

  assign sfifo_rcstage_push = sfifo_adstage_pop;
  assign sfifo_rcstage_wdata = {adstage_key,adstage_v,sfifo_bencack_bits,
                                adstage_rc,adstage_fips,adstage_glast,
                                sfifo_bencack_inst_id,sfifo_bencack_ccmd};

  assign sfifo_rcstage_pop = sfifo_rcstage_not_empty && (upd_gen_ack_i || !rcstage_glast);

  assign {rcstage_key,rcstage_v,rcstage_bits,rcstage_rc,rcstage_fips,rcstage_glast,
          rcstage_inst_id,rcstage_ccmd} = sfifo_rcstage_rdata;


  assign ctr_drbg_gen_sfifo_grcstage_err_o =
         {(sfifo_rcstage_push && sfifo_rcstage_full),
          (sfifo_rcstage_pop && !sfifo_rcstage_not_empty),
          (sfifo_rcstage_full && !sfifo_rcstage_not_empty)};

  assign gen_upd_rdy_o = sfifo_rcstage_not_empty && !sfifo_genbits_full;


  //--------------------------------------------
  // final cmd block processing
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(GenbitsFifoWidth),
    .Pass(0),
    .Depth(GenbitsFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_genbits (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (!ctr_drbg_gen_enable_i),
    .wvalid_i       (sfifo_genbits_push),
    .wready_o       (),
    .wdata_i        (sfifo_genbits_wdata),
    .rvalid_o       (sfifo_genbits_not_empty),
    .rready_i       (sfifo_genbits_pop),
    .rdata_o        (sfifo_genbits_rdata),
    .full_o         (sfifo_genbits_full),
    .depth_o        (),
    .err_o          ()
  );

  assign sfifo_genbits_push = sfifo_rcstage_pop;

  assign rcstage_rc_plus1 = (rcstage_rc+1);

  assign sfifo_genbits_wdata = rcstage_glast ?
                               {rcstage_fips,rcstage_bits,upd_gen_key_i,upd_gen_v_i,
                                rcstage_rc_plus1,upd_gen_inst_id_i,upd_gen_ccmd_i} :
                               {rcstage_fips,rcstage_bits,rcstage_key,rcstage_v,
                                rcstage_rc,rcstage_inst_id,rcstage_ccmd};

  assign sfifo_genbits_pop = ctr_drbg_gen_rdy_i && sfifo_genbits_not_empty;
  assign {ctr_drbg_gen_fips_o,ctr_drbg_gen_bits_o,
          ctr_drbg_gen_key_o,ctr_drbg_gen_v_o,ctr_drbg_gen_rc_o,
          ctr_drbg_gen_inst_id_o,ctr_drbg_gen_ccmd_o} = sfifo_genbits_rdata;

  assign ctr_drbg_gen_sfifo_ggenbits_err_o =
         {(sfifo_genbits_push && sfifo_genbits_full),
         (sfifo_genbits_pop && !sfifo_genbits_not_empty),
         (sfifo_genbits_full && !sfifo_genbits_not_empty)};

  // block ack
  assign ctr_drbg_gen_ack_o = sfifo_genbits_pop;

  assign ctr_drbg_gen_sts_o = sfifo_genbits_pop && (
         (ctr_drbg_gen_ccmd_o == INV) ||
         (ctr_drbg_gen_ccmd_o == INS) ||
         (ctr_drbg_gen_ccmd_o == RES) ||
         (ctr_drbg_gen_ccmd_o == UPD) ||
         (ctr_drbg_gen_ccmd_o == UNI));

  // Make sure that the state machine has a stable error state. This means that after the error
  // state is entered it will not exit it unless a reset signal is received.
  `ASSERT(CsrngDrbgGenErrorStStable_A, state_q == ReqError |=> $stable(state_q))
  // If in error state, the error output must be high.
  `ASSERT(CsrngDrbgGenErrorOutput_A,
          !(state_q inside {ReqIdle, ReqSend, ESHalt}) |-> ctr_drbg_gen_sm_err_o)
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng core module
//


module csrng_core import csrng_pkg::*; #(
  parameter aes_pkg::sbox_impl_e SBoxImpl = aes_pkg::SBoxImplLut,
  parameter int NHwApps = 2,
  parameter cs_keymgr_div_t RndCnstCsKeymgrDivNonProduction = CsKeymgrDivWidth'(0),
  parameter cs_keymgr_div_t RndCnstCsKeymgrDivProduction = CsKeymgrDivWidth'(0)
) (
  input logic                                     clk_i,
  input logic                                     rst_ni,

  input  csrng_reg_pkg::csrng_reg2hw_t            reg2hw,
  output csrng_reg_pkg::csrng_hw2reg_t            hw2reg,

  // Efuse Interface
  input  prim_mubi_pkg::mubi8_t                   otp_en_csrng_sw_app_read_i,

  // Lifecycle broadcast inputs
  input  lc_ctrl_pkg::lc_tx_t                     lc_hw_debug_en_i,

  // Entropy Interface
  output entropy_src_pkg::entropy_src_hw_if_req_t entropy_src_hw_if_o,
  input  entropy_src_pkg::entropy_src_hw_if_rsp_t entropy_src_hw_if_i,

  // Entropy Interface
  input  entropy_src_pkg::cs_aes_halt_req_t       cs_aes_halt_i,
  output entropy_src_pkg::cs_aes_halt_rsp_t       cs_aes_halt_o,

  // Application Interfaces
  input  csrng_req_t [NHwApps-1:0]                csrng_cmd_i,
  output csrng_rsp_t [NHwApps-1:0]                csrng_cmd_o,

  // Alerts

  output logic                                    recov_alert_test_o,
  output logic                                    fatal_alert_test_o,
  output logic                                    recov_alert_o,
  output logic                                    fatal_alert_o,

  output logic                                    intr_cs_cmd_req_done_o,
  output logic                                    intr_cs_entropy_req_o,
  output logic                                    intr_cs_hw_inst_exc_o,
  output logic                                    intr_cs_fatal_err_o
);

  import csrng_reg_pkg::*;

  import prim_mubi_pkg::mubi4_t;
  import prim_mubi_pkg::mubi4_test_true_strict;
  import prim_mubi_pkg::mubi4_test_invalid;

  localparam int NApps = NHwApps + 1;
  localparam int AppCmdWidth = 32;
  localparam int AppCmdFifoDepth = 2;
  localparam int GenBitsWidth = 128;
  localparam int Cmd = 3;
  localparam int StateId = 4;
  localparam int KeyLen = 256;
  localparam int BlkLen = 128;
  localparam int SeedLen = 384;
  localparam int CtrLen = 32;
  localparam int NBlkEncArbReqs = 2;
  localparam int BlkEncArbWidth = KeyLen+BlkLen+StateId+Cmd;
  localparam int NUpdateArbReqs = 2;
  localparam int UpdateArbWidth = KeyLen+BlkLen+SeedLen+StateId+Cmd;
  localparam int MaxClen = 12;
  localparam int ADataDepthWidth = SeedLen/AppCmdWidth;
  localparam unsigned ADataDepthClog = $clog2(ADataDepthWidth)+1;
  localparam int CsEnableCopies = 51;
  localparam int LcHwDebugCopies = 1;
  localparam int Flag0Copies = 3;

  // signals
  // interrupt signals
  logic                        event_cs_cmd_req_done;
  logic                        event_cs_entropy_req;
  logic                        event_cs_hw_inst_exc;
  logic                        event_cs_fatal_err;
  logic [CsEnableCopies-1:1]   cs_enable_fo;
  logic [Flag0Copies-1:0]      flag0_fo;
  logic                        acmd_flag0_pfa;
  logic                        cs_enable_pfa;
  logic                        sw_app_enable;
  logic                        sw_app_enable_pfe;
  logic                        sw_app_enable_pfa;
  logic                        read_int_state;
  logic                        read_int_state_pfe;
  logic                        read_int_state_pfa;
  logic                        recov_alert_event;
  logic                        acmd_avail;
  logic                        acmd_sop;
  logic                        acmd_mop;
  logic                        acmd_eop;

  logic                        cmd_blk_select;
  logic                        gen_blk_select;
  logic                        state_db_wr_req_rdy;
  logic                        state_db_wr_req;
  logic [StateId-1:0]          state_db_wr_inst_id;
  logic [KeyLen-1:0]           state_db_wr_key;
  logic [BlkLen-1:0]           state_db_wr_v;
  logic [CtrLen-1:0]           state_db_wr_rc;
  logic                        state_db_wr_sts;
  logic                        state_db_wr_fips;
  logic [Cmd-1:0]              state_db_wr_ccmd;

  logic [AppCmdWidth-1:0]      acmd_bus;

  logic [SeedLen-1:0]          packer_adata;
  logic [ADataDepthClog-1:0]   packer_adata_depth;
  logic                        packer_adata_pop;
  logic                        packer_adata_clr;
  logic [SeedLen-1:0]          seed_diversification;

  logic                        cmd_entropy_req;
  logic                        cmd_entropy_avail;
  logic                        cmd_entropy_fips;
  logic [SeedLen-1:0]          cmd_entropy;

  logic                        cmd_result_wr_req;
  logic                        cmd_result_ack;
  logic                        cmd_result_ack_sts;
  logic [Cmd-1:0]              cmd_result_ccmd;
  logic                        cmd_result_ack_rdy;
  logic [StateId-1:0]          cmd_result_inst_id;
  logic                        cmd_result_glast;
  logic                        cmd_result_fips;
  logic [SeedLen-1:0]          cmd_result_adata;
  logic [KeyLen-1:0]           cmd_result_key;
  logic [BlkLen-1:0]           cmd_result_v;
  logic [CtrLen-1:0]           cmd_result_rc;

  logic                        state_db_sts_ack;
  logic                        state_db_sts_sts;
  logic [StateId-1:0]          state_db_sts_id;

  logic                        gen_result_wr_req;
  logic                        gen_result_ack_sts;
  logic                        gen_result_ack_rdy;
  logic [Cmd-1:0]              gen_result_ccmd;
  logic [StateId-1:0]          gen_result_inst_id;
  logic                        gen_result_fips;
  logic [KeyLen-1:0]           gen_result_key;
  logic [BlkLen-1:0]           gen_result_v;
  logic [CtrLen-1:0]           gen_result_rc;
  logic [BlkLen-1:0]           gen_result_bits;

  logic                        acmd_accept;
  logic                        instant_req;
  logic                        reseed_req;
  logic                        generate_req;
  logic                        update_req;
  logic                        uninstant_req;
  logic                        clr_adata_packer;
  logic [Cmd-1:0]              ctr_drbg_cmd_ccmd;
  logic                        ctr_drbg_cmd_req;
  logic                        ctr_drbg_gen_req;
  logic                        ctr_drbg_gen_req_rdy;
  logic                        ctr_drbg_cmd_req_rdy;
  logic                        ctr_drbg_cmd_sfifo_cmdreq_err_sum;
  logic [2:0]                  ctr_drbg_cmd_sfifo_cmdreq_err;
  logic                        ctr_drbg_cmd_sfifo_rcstage_err_sum;
  logic [2:0]                  ctr_drbg_cmd_sfifo_rcstage_err;
  logic                        ctr_drbg_cmd_sfifo_keyvrc_err_sum;
  logic [2:0]                  ctr_drbg_cmd_sfifo_keyvrc_err;
  logic                        ctr_drbg_upd_sfifo_updreq_err_sum;
  logic [2:0]                  ctr_drbg_upd_sfifo_updreq_err;
  logic                        ctr_drbg_upd_sfifo_bencreq_err_sum;
  logic [2:0]                  ctr_drbg_upd_sfifo_bencreq_err;
  logic                        ctr_drbg_upd_sfifo_bencack_err_sum;
  logic [2:0]                  ctr_drbg_upd_sfifo_bencack_err;
  logic                        ctr_drbg_upd_sfifo_pdata_err_sum;
  logic [2:0]                  ctr_drbg_upd_sfifo_pdata_err;
  logic                        ctr_drbg_upd_sfifo_final_err_sum;
  logic [2:0]                  ctr_drbg_upd_sfifo_final_err;
  logic                        ctr_drbg_gen_sfifo_gbencack_err_sum;
  logic [2:0]                  ctr_drbg_gen_sfifo_gbencack_err;
  logic                        ctr_drbg_gen_sfifo_grcstage_err_sum;
  logic [2:0]                  ctr_drbg_gen_sfifo_grcstage_err;
  logic                        ctr_drbg_gen_sfifo_ggenreq_err_sum;
  logic [2:0]                  ctr_drbg_gen_sfifo_ggenreq_err;
  logic                        ctr_drbg_gen_sfifo_gadstage_err_sum;
  logic [2:0]                  ctr_drbg_gen_sfifo_gadstage_err;
  logic                        ctr_drbg_gen_sfifo_ggenbits_err_sum;
  logic [2:0]                  ctr_drbg_gen_sfifo_ggenbits_err;
  logic                        block_encrypt_sfifo_blkenc_err_sum;
  logic [2:0]                  block_encrypt_sfifo_blkenc_err;
  logic                        cmd_gen_cnt_err_sum;
  logic                        cmd_stage_sm_err_sum;
  logic                        main_sm_err_sum;
  logic                        cs_main_sm_alert;
  logic                        cs_main_sm_err;
  logic [MainSmStateWidth-1:0] cs_main_sm_state;
  logic                        drbg_gen_sm_err_sum;
  logic                        drbg_gen_sm_err;
  logic                        drbg_updbe_sm_err_sum;
  logic                        drbg_updbe_sm_err;
  logic                        drbg_updob_sm_err_sum;
  logic                        drbg_updob_sm_err;
  logic                        aes_cipher_sm_err_sum;
  logic                        aes_cipher_sm_err;
  logic                        fifo_write_err_sum;
  logic                        fifo_read_err_sum;
  logic                        fifo_status_err_sum;

  logic [KeyLen-1:0]           state_db_rd_key;
  logic [BlkLen-1:0]           state_db_rd_v;
  logic [CtrLen-1:0]           state_db_rd_rc;
  logic                        state_db_rd_fips;
  logic [2:0]                  acmd_hold;
  logic [3:0]                  shid;
  logic                        gen_last;
  mubi4_t                      flag0;

  // blk encrypt arbiter
  logic [Cmd-1:0]              updblk_benblk_cmd_arb_din;
  logic [StateId-1:0]          updblk_benblk_id_arb_din;
  logic [BlkLen-1:0]           updblk_benblk_v_arb_din;
  logic [KeyLen-1:0]           updblk_benblk_key_arb_din;
  logic                        updblk_benblk_arb_req;
  logic                        updblk_benblk_arb_req_rdy;
  logic                        benblk_updblk_ack;
  logic                        updblk_benblk_ack_rdy;

  logic [Cmd-1:0]              genblk_benblk_cmd_arb_din;
  logic [StateId-1:0]          genblk_benblk_id_arb_din;
  logic [BlkLen-1:0]           genblk_benblk_v_arb_din;
  logic [KeyLen-1:0]           genblk_benblk_key_arb_din;
  logic                        genblk_benblk_arb_req;
  logic                        genblk_benblk_arb_req_rdy;
  logic                        benblk_genblk_ack;
  logic                        genblk_benblk_ack_rdy;

  logic [BlkEncArbWidth-1:0]   benblk_arb_din [2];
  logic [BlkEncArbWidth-1:0]   benblk_arb_data;
  logic [KeyLen-1:0]           benblk_arb_key;
  logic [BlkLen-1:0]           benblk_arb_v;
  logic [StateId-1:0]          benblk_arb_inst_id;
  logic [Cmd-1:0]              benblk_arb_cmd;
  logic                        benblk_arb_vld;
  logic                        benblk_ack;
  logic                        benblk_ack_rdy;
  logic                        benblk_arb_rdy;
  logic [Cmd-1:0]              benblk_cmd;
  logic [StateId-1:0]          benblk_inst_id;
  logic [BlkLen-1:0]           benblk_v;

  // update arbiter
  logic [Cmd-1:0]              cmdblk_updblk_ccmd_arb_din;
  logic [StateId-1:0]          cmdblk_updblk_id_arb_din;
  logic [BlkLen-1:0]           cmdblk_updblk_v_arb_din;
  logic [KeyLen-1:0]           cmdblk_updblk_key_arb_din;
  logic [SeedLen-1:0]          cmdblk_updblk_pdata_arb_din;
  logic                        cmdblk_updblk_arb_req;
  logic                        updblk_cmdblk_arb_req_rdy;
  logic                        updblk_cmdblk_ack;
  logic                        cmdblk_updblk_ack_rdy;

  logic [Cmd-1:0]              genblk_updblk_ccmd_arb_din;
  logic [StateId-1:0]          genblk_updblk_id_arb_din;
  logic [BlkLen-1:0]           genblk_updblk_v_arb_din;
  logic [KeyLen-1:0]           genblk_updblk_key_arb_din;
  logic [SeedLen-1:0]          genblk_updblk_pdata_arb_din;
  logic                        genblk_updblk_arb_req;
  logic                        updblk_genblk_arb_req_rdy;
  logic                        updblk_genblk_ack;
  logic                        genblk_updblk_ack_rdy;

  logic [UpdateArbWidth-1:0]   updblk_arb_din [2];
  logic [UpdateArbWidth-1:0]   updblk_arb_data;
  logic [KeyLen-1:0]           updblk_arb_key;
  logic [BlkLen-1:0]           updblk_arb_v;
  logic [SeedLen-1:0]          updblk_arb_pdata;
  logic [StateId-1:0]          updblk_arb_inst_id;
  logic [Cmd-1:0]              updblk_arb_ccmd;
  logic                        updblk_arb_vld;
  logic                        updblk_ack;
  logic                        updblk_ack_rdy;
  logic                        updblk_arb_rdy;
  logic [Cmd-1:0]              updblk_ccmd;
  logic [StateId-1:0]          updblk_inst_id;
  logic [KeyLen-1:0]           updblk_key;
  logic [BlkLen-1:0]           updblk_v;

  logic [2:0]                  cmd_stage_sfifo_cmd_err[NApps];
  logic [NApps-1:0]            cmd_stage_sfifo_cmd_err_sum;
  logic [NApps-1:0]            cmd_stage_sfifo_cmd_err_wr;
  logic [NApps-1:0]            cmd_stage_sfifo_cmd_err_rd;
  logic [NApps-1:0]            cmd_stage_sfifo_cmd_err_st;
  logic [2:0]                  cmd_stage_sfifo_genbits_err[NApps];
  logic [NApps-1:0]            cmd_stage_sfifo_genbits_err_sum;
  logic [NApps-1:0]            cmd_stage_sfifo_genbits_err_wr;
  logic [NApps-1:0]            cmd_stage_sfifo_genbits_err_rd;
  logic [NApps-1:0]            cmd_stage_sfifo_genbits_err_st;
  logic [NApps-1:0]            cmd_gen_cnt_err;
  logic [NApps-1:0]            cmd_stage_sm_err;
  logic                        ctr_drbg_upd_v_ctr_err;
  logic                        ctr_drbg_gen_v_ctr_err;

  logic [NApps-1:0]          cmd_stage_vld;
  logic [StateId-1:0]        cmd_stage_shid[NApps];
  logic [AppCmdWidth-1:0]    cmd_stage_bus[NApps];
  logic [NApps-1:0]          cmd_stage_rdy;
  logic [NApps-1:0]          cmd_arb_req;
  logic [NApps-1:0]          cmd_arb_gnt;
  logic [$clog2(NApps)-1:0]  cmd_arb_idx;
  logic [NApps-1:0]          cmd_arb_sop;
  logic [NApps-1:0]          cmd_arb_mop;
  logic [NApps-1:0]          cmd_arb_eop;
  logic [AppCmdWidth-1:0]    cmd_arb_bus[NApps];
  logic [NApps-1:0]          cmd_core_ack;
  logic [NApps-1:0]          cmd_core_ack_sts;
  logic [NApps-1:0]          cmd_stage_ack;
  logic [NApps-1:0]          cmd_stage_ack_sts;
  logic [NApps-1:0]          genbits_core_vld;
  logic [GenBitsWidth-1:0]   genbits_core_bus[NApps];
  logic [NApps-1:0]          genbits_core_fips;
  logic [NApps-1:0]          genbits_stage_vld;
  logic [NApps-1:0]          genbits_stage_fips;
  logic [GenBitsWidth-1:0]   genbits_stage_bus[NApps];
  logic [NApps-1:0]          genbits_stage_rdy;
  logic                      genbits_stage_vldo_sw;
  logic                      genbits_stage_bus_rd_sw;
  logic [31:0]               genbits_stage_bus_sw;
  logic                      genbits_stage_fips_sw;

  logic [15:0]               hw_exception_sts;
  logic [LcHwDebugCopies-1:0]lc_hw_debug_on_fo;
  logic                      state_db_is_dump_en;
  logic                      state_db_reg_rd_sel;
  logic                      state_db_reg_rd_id_pulse;
  logic [StateId-1:0]        state_db_reg_rd_id;
  logic [31:0]               state_db_reg_rd_val;

  logic [30:0]               err_code_test_bit;
  logic                      ctr_drbg_upd_es_ack;
  logic                      ctr_drbg_gen_es_ack;
  logic                      block_encrypt_quiet;

  logic                      cs_rdata_capt_vld;
  logic                      cs_bus_cmp_alert;
  logic                      cmd_rdy;
  logic [1:0]                efuse_sw_app_enable;

  logic                      unused_err_code_test_bit;
  logic                      unused_reg2hw_genbits;
  logic                      unused_int_state_val;

  prim_mubi_pkg::mubi8_t [1:0] en_csrng_sw_app_read;
  prim_mubi_pkg::mubi4_t [CsEnableCopies-1:0] mubi_cs_enable_fanout;
  prim_mubi_pkg::mubi4_t [Flag0Copies-1:0] mubi_flag0_fanout;

  // flops
  logic [2:0]                acmd_q, acmd_d;
  logic [3:0]                shid_q, shid_d;
  logic                      gen_last_q, gen_last_d;
  mubi4_t                    flag0_q, flag0_d;
  logic [$clog2(NApps)-1:0]  cmd_arb_idx_q, cmd_arb_idx_d;
  logic                      statedb_wr_select_q, statedb_wr_select_d;
  logic                      genbits_stage_fips_sw_q, genbits_stage_fips_sw_d;
  logic                      cmd_req_dly_q, cmd_req_dly_d;
  logic [Cmd-1:0]            cmd_req_ccmd_dly_q, cmd_req_ccmd_dly_d;
  logic                      cs_aes_halt_q, cs_aes_halt_d;
  logic [SeedLen-1:0]        entropy_src_seed_q, entropy_src_seed_d;
  logic                      entropy_src_fips_q, entropy_src_fips_d;
  logic [63:0]               cs_rdata_capt_q, cs_rdata_capt_d;
  logic                      cs_rdata_capt_vld_q, cs_rdata_capt_vld_d;
  logic                      sw_rdy_sts_q, sw_rdy_sts_d;

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      acmd_q                  <= '0;
      shid_q                  <= '0;
      gen_last_q              <= '0;
      flag0_q                 <= prim_mubi_pkg::MuBi4False;
      cmd_arb_idx_q           <= '0;
      statedb_wr_select_q     <= '0;
      genbits_stage_fips_sw_q <= '0;
      cmd_req_dly_q           <= '0;
      cmd_req_ccmd_dly_q      <= '0;
      cs_aes_halt_q           <= '0;
      entropy_src_seed_q      <= '0;
      entropy_src_fips_q      <= '0;
      cs_rdata_capt_q         <= '0;
      cs_rdata_capt_vld_q     <= '0;
      sw_rdy_sts_q            <= '0;
    end else begin
      acmd_q                  <= acmd_d;
      shid_q                  <= shid_d;
      gen_last_q              <= gen_last_d;
      flag0_q                 <= flag0_d;
      cmd_arb_idx_q           <= cmd_arb_idx_d;
      statedb_wr_select_q     <= statedb_wr_select_d;
      genbits_stage_fips_sw_q <= genbits_stage_fips_sw_d;
      cmd_req_dly_q           <= cmd_req_dly_d;
      cmd_req_ccmd_dly_q      <= cmd_req_ccmd_dly_d;
      cs_aes_halt_q           <= cs_aes_halt_d;
      entropy_src_seed_q      <= entropy_src_seed_d;
      entropy_src_fips_q      <= entropy_src_fips_d;
      cs_rdata_capt_q         <= cs_rdata_capt_d;
      cs_rdata_capt_vld_q     <= cs_rdata_capt_vld_d;
      sw_rdy_sts_q            <= sw_rdy_sts_d;
    end

  //--------------------------------------------
  // instantiate interrupt hardware primitives
  //--------------------------------------------
  // All TLUL interrupts are collect in the section.

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_cs_cmd_req_done (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_cs_cmd_req_done),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.cs_cmd_req_done.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.cs_cmd_req_done.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.cs_cmd_req_done.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.cs_cmd_req_done.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.cs_cmd_req_done.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.cs_cmd_req_done.d),
    .intr_o                 (intr_cs_cmd_req_done_o)
  );

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_cs_entropy_req (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_cs_entropy_req),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.cs_entropy_req.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.cs_entropy_req.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.cs_entropy_req.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.cs_entropy_req.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.cs_entropy_req.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.cs_entropy_req.d),
    .intr_o                 (intr_cs_entropy_req_o)
  );


  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_cs_hw_inst_exc (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_cs_hw_inst_exc),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.cs_hw_inst_exc.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.cs_hw_inst_exc.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.cs_hw_inst_exc.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.cs_hw_inst_exc.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.cs_hw_inst_exc.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.cs_hw_inst_exc.d),
    .intr_o                 (intr_cs_hw_inst_exc_o)
  );


  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_cs_fatal_err (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_cs_fatal_err),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.cs_fatal_err.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.cs_fatal_err.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.cs_fatal_err.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.cs_fatal_err.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.cs_fatal_err.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.cs_fatal_err.d),
    .intr_o                 (intr_cs_fatal_err_o)
  );

  // set the interrupt sources
  assign event_cs_fatal_err = (cs_enable_fo[1]  && (
         (|cmd_stage_sfifo_cmd_err_sum) ||
         (|cmd_stage_sfifo_genbits_err_sum) ||
         ctr_drbg_cmd_sfifo_cmdreq_err_sum ||
         ctr_drbg_cmd_sfifo_rcstage_err_sum ||
         ctr_drbg_cmd_sfifo_keyvrc_err_sum ||
         ctr_drbg_upd_sfifo_updreq_err_sum ||
         ctr_drbg_upd_sfifo_bencreq_err_sum ||
         ctr_drbg_upd_sfifo_bencack_err_sum ||
         ctr_drbg_upd_sfifo_pdata_err_sum ||
         ctr_drbg_upd_sfifo_final_err_sum ||
         ctr_drbg_gen_sfifo_gbencack_err_sum ||
         ctr_drbg_gen_sfifo_grcstage_err_sum ||
         ctr_drbg_gen_sfifo_ggenreq_err_sum ||
         ctr_drbg_gen_sfifo_gadstage_err_sum ||
         ctr_drbg_gen_sfifo_ggenbits_err_sum ||
         block_encrypt_sfifo_blkenc_err_sum ||
         fifo_write_err_sum ||
         fifo_read_err_sum ||
         fifo_status_err_sum)) ||
         // errs not gated by cs_enable
         cmd_stage_sm_err_sum ||
         main_sm_err_sum ||
         drbg_gen_sm_err_sum ||
         drbg_updbe_sm_err_sum ||
         drbg_updob_sm_err_sum ||
         aes_cipher_sm_err_sum ||
         cmd_gen_cnt_err_sum;

  // set fifo errors that are single instances of source
  assign ctr_drbg_cmd_sfifo_cmdreq_err_sum = (|ctr_drbg_cmd_sfifo_cmdreq_err) ||
         err_code_test_bit[2];
  assign ctr_drbg_cmd_sfifo_rcstage_err_sum = (|ctr_drbg_cmd_sfifo_rcstage_err) ||
         err_code_test_bit[3];
  assign ctr_drbg_cmd_sfifo_keyvrc_err_sum = (|ctr_drbg_cmd_sfifo_keyvrc_err) ||
         err_code_test_bit[4];
  assign ctr_drbg_upd_sfifo_updreq_err_sum = (|ctr_drbg_upd_sfifo_updreq_err) ||
         err_code_test_bit[5];
  assign ctr_drbg_upd_sfifo_bencreq_err_sum = (|ctr_drbg_upd_sfifo_bencreq_err) ||
         err_code_test_bit[6];
  assign ctr_drbg_upd_sfifo_bencack_err_sum = (|ctr_drbg_upd_sfifo_bencack_err) ||
         err_code_test_bit[7];
  assign ctr_drbg_upd_sfifo_pdata_err_sum = (|ctr_drbg_upd_sfifo_pdata_err) ||
         err_code_test_bit[8];
  assign ctr_drbg_upd_sfifo_final_err_sum = (|ctr_drbg_upd_sfifo_final_err) ||
         err_code_test_bit[9];
  assign ctr_drbg_gen_sfifo_gbencack_err_sum = (|ctr_drbg_gen_sfifo_gbencack_err) ||
         err_code_test_bit[10];
  assign ctr_drbg_gen_sfifo_grcstage_err_sum = (|ctr_drbg_gen_sfifo_grcstage_err) ||
         err_code_test_bit[11];
  assign ctr_drbg_gen_sfifo_ggenreq_err_sum = (|ctr_drbg_gen_sfifo_ggenreq_err) ||
         err_code_test_bit[12];
  assign ctr_drbg_gen_sfifo_gadstage_err_sum = (|ctr_drbg_gen_sfifo_gadstage_err) ||
         err_code_test_bit[13];
  assign ctr_drbg_gen_sfifo_ggenbits_err_sum = (|ctr_drbg_gen_sfifo_ggenbits_err) ||
         err_code_test_bit[14];
  assign block_encrypt_sfifo_blkenc_err_sum = (|block_encrypt_sfifo_blkenc_err) ||
         err_code_test_bit[15];
  assign cmd_stage_sm_err_sum = (|cmd_stage_sm_err) ||
         err_code_test_bit[20];
  assign main_sm_err_sum = cs_main_sm_err ||
         err_code_test_bit[21];
  assign drbg_gen_sm_err_sum = drbg_gen_sm_err ||
         err_code_test_bit[22];
  assign drbg_updbe_sm_err_sum = drbg_updbe_sm_err ||
         err_code_test_bit[23];
  assign drbg_updob_sm_err_sum = drbg_updob_sm_err ||
         err_code_test_bit[24];
  assign aes_cipher_sm_err_sum = aes_cipher_sm_err ||
         err_code_test_bit[25];
  assign cmd_gen_cnt_err_sum = (|cmd_gen_cnt_err) || ctr_drbg_gen_v_ctr_err ||
         ctr_drbg_upd_v_ctr_err || err_code_test_bit[26];
  assign fifo_write_err_sum =
         block_encrypt_sfifo_blkenc_err[2] ||
         ctr_drbg_gen_sfifo_ggenbits_err[2] ||
         ctr_drbg_gen_sfifo_gadstage_err[2] ||
         ctr_drbg_gen_sfifo_ggenreq_err[2] ||
         ctr_drbg_gen_sfifo_grcstage_err[2] ||
         ctr_drbg_gen_sfifo_gbencack_err[2] ||
         ctr_drbg_upd_sfifo_final_err[2] ||
         ctr_drbg_upd_sfifo_pdata_err[2] ||
         ctr_drbg_upd_sfifo_bencack_err[2] ||
         ctr_drbg_upd_sfifo_bencreq_err[2] ||
         ctr_drbg_upd_sfifo_updreq_err[2] ||
         ctr_drbg_cmd_sfifo_keyvrc_err[2] ||
         ctr_drbg_cmd_sfifo_rcstage_err[2] ||
         ctr_drbg_cmd_sfifo_cmdreq_err[2] ||
         (|cmd_stage_sfifo_genbits_err_wr) ||
         (|cmd_stage_sfifo_cmd_err_wr) ||
         err_code_test_bit[28];
  assign fifo_read_err_sum =
         block_encrypt_sfifo_blkenc_err[1] ||
         ctr_drbg_gen_sfifo_ggenbits_err[1] ||
         ctr_drbg_gen_sfifo_gadstage_err[1] ||
         ctr_drbg_gen_sfifo_ggenreq_err[1] ||
         ctr_drbg_gen_sfifo_grcstage_err[1] ||
         ctr_drbg_gen_sfifo_gbencack_err[1] ||
         ctr_drbg_upd_sfifo_final_err[1] ||
         ctr_drbg_upd_sfifo_pdata_err[1] ||
         ctr_drbg_upd_sfifo_bencack_err[1] ||
         ctr_drbg_upd_sfifo_bencreq_err[1] ||
         ctr_drbg_upd_sfifo_updreq_err[1] ||
         ctr_drbg_cmd_sfifo_keyvrc_err[1] ||
         ctr_drbg_cmd_sfifo_rcstage_err[1] ||
         ctr_drbg_cmd_sfifo_cmdreq_err[1] ||
         (|cmd_stage_sfifo_genbits_err_rd) ||
         (|cmd_stage_sfifo_cmd_err_rd) ||
         err_code_test_bit[29];
  assign fifo_status_err_sum =
         block_encrypt_sfifo_blkenc_err[0] ||
         ctr_drbg_gen_sfifo_ggenbits_err[0] ||
         ctr_drbg_gen_sfifo_gadstage_err[0] ||
         ctr_drbg_gen_sfifo_ggenreq_err[0] ||
         ctr_drbg_gen_sfifo_grcstage_err[0] ||
         ctr_drbg_gen_sfifo_gbencack_err[0] ||
         ctr_drbg_upd_sfifo_final_err[0] ||
         ctr_drbg_upd_sfifo_pdata_err[0] ||
         ctr_drbg_upd_sfifo_bencack_err[0] ||
         ctr_drbg_upd_sfifo_bencreq_err[0] ||
         ctr_drbg_upd_sfifo_updreq_err[0] ||
         ctr_drbg_cmd_sfifo_keyvrc_err[0] ||
         ctr_drbg_cmd_sfifo_rcstage_err[0] ||
         ctr_drbg_cmd_sfifo_cmdreq_err[0] ||
         (|cmd_stage_sfifo_genbits_err_st) ||
         (|cmd_stage_sfifo_cmd_err_st) ||
         err_code_test_bit[30];

  // set the err code source bits
  assign hw2reg.err_code.sfifo_cmd_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_cmd_err.de = cs_enable_fo[2] &&
         (|cmd_stage_sfifo_cmd_err_sum);

  assign hw2reg.err_code.sfifo_genbits_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_genbits_err.de = cs_enable_fo[3] &&
         (|cmd_stage_sfifo_genbits_err_sum);

  assign hw2reg.err_code.sfifo_cmdreq_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_cmdreq_err.de = cs_enable_fo[4] &&
         ctr_drbg_cmd_sfifo_cmdreq_err_sum;

  assign hw2reg.err_code.sfifo_rcstage_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_rcstage_err.de = cs_enable_fo[5] &&
         ctr_drbg_cmd_sfifo_rcstage_err_sum;

  assign hw2reg.err_code.sfifo_keyvrc_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_keyvrc_err.de = cs_enable_fo[6] &&
         ctr_drbg_cmd_sfifo_keyvrc_err_sum;

  assign hw2reg.err_code.sfifo_updreq_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_updreq_err.de = cs_enable_fo[7] &&
         ctr_drbg_upd_sfifo_updreq_err_sum;

  assign hw2reg.err_code.sfifo_bencreq_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_bencreq_err.de = cs_enable_fo[8] &&
         ctr_drbg_upd_sfifo_bencreq_err_sum;

  assign hw2reg.err_code.sfifo_bencack_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_bencack_err.de = cs_enable_fo[9] &&
         ctr_drbg_upd_sfifo_bencack_err_sum;

  assign hw2reg.err_code.sfifo_pdata_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_pdata_err.de = cs_enable_fo[10] &&
         ctr_drbg_upd_sfifo_pdata_err_sum;

  assign hw2reg.err_code.sfifo_final_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_final_err.de = cs_enable_fo[11] &&
         ctr_drbg_upd_sfifo_final_err_sum;

  assign hw2reg.err_code.sfifo_gbencack_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_gbencack_err.de = cs_enable_fo[12] &&
         ctr_drbg_gen_sfifo_gbencack_err_sum;

  assign hw2reg.err_code.sfifo_grcstage_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_grcstage_err.de = cs_enable_fo[13] &&
         ctr_drbg_gen_sfifo_grcstage_err_sum;

  assign hw2reg.err_code.sfifo_ggenreq_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_ggenreq_err.de = cs_enable_fo[14] &&
         ctr_drbg_gen_sfifo_ggenreq_err_sum;

  assign hw2reg.err_code.sfifo_gadstage_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_gadstage_err.de = cs_enable_fo[15] &&
         ctr_drbg_gen_sfifo_gadstage_err_sum;

  assign hw2reg.err_code.sfifo_ggenbits_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_ggenbits_err.de = cs_enable_fo[16] &&
         ctr_drbg_gen_sfifo_ggenbits_err_sum;

  assign hw2reg.err_code.sfifo_blkenc_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_blkenc_err.de = cs_enable_fo[17] &&
         block_encrypt_sfifo_blkenc_err_sum;

  assign hw2reg.err_code.cmd_stage_sm_err.d = 1'b1;
  assign hw2reg.err_code.cmd_stage_sm_err.de = cs_enable_fo[18] &&
         cmd_stage_sm_err_sum;

  assign hw2reg.err_code.main_sm_err.d = 1'b1;
  assign hw2reg.err_code.main_sm_err.de = cs_enable_fo[19] &&
         main_sm_err_sum;

  assign hw2reg.err_code.drbg_gen_sm_err.d = 1'b1;
  assign hw2reg.err_code.drbg_gen_sm_err.de = cs_enable_fo[20] &&
         drbg_gen_sm_err_sum;

  assign hw2reg.err_code.drbg_updbe_sm_err.d = 1'b1;
  assign hw2reg.err_code.drbg_updbe_sm_err.de = cs_enable_fo[21] &&
         drbg_updbe_sm_err_sum;

  assign hw2reg.err_code.drbg_updob_sm_err.d = 1'b1;
  assign hw2reg.err_code.drbg_updob_sm_err.de = cs_enable_fo[22] &&
         drbg_updob_sm_err_sum;

  assign hw2reg.err_code.aes_cipher_sm_err.d = 1'b1;
  assign hw2reg.err_code.aes_cipher_sm_err.de = cs_enable_fo[23] &&
         aes_cipher_sm_err_sum;

  assign hw2reg.err_code.cmd_gen_cnt_err.d = 1'b1;
  assign hw2reg.err_code.cmd_gen_cnt_err.de = cmd_gen_cnt_err_sum;


 // set the err code type bits
  assign hw2reg.err_code.fifo_write_err.d = 1'b1;
  assign hw2reg.err_code.fifo_write_err.de = cs_enable_fo[24] && fifo_write_err_sum;

  assign hw2reg.err_code.fifo_read_err.d = 1'b1;
  assign hw2reg.err_code.fifo_read_err.de = cs_enable_fo[25] && fifo_read_err_sum;

  assign hw2reg.err_code.fifo_state_err.d = 1'b1;
  assign hw2reg.err_code.fifo_state_err.de = cs_enable_fo[26] && fifo_status_err_sum;

  // Error forcing
  for (genvar i = 0; i < 31; i = i+1) begin : gen_err_code_test_bit
    assign err_code_test_bit[i] = (reg2hw.err_code_test.q == i) && reg2hw.err_code_test.qe;
  end : gen_err_code_test_bit

  // alert - send all interrupt sources to the alert for the fatal case
  assign fatal_alert_o = event_cs_fatal_err;

  // alert test
  assign recov_alert_test_o = {
    reg2hw.alert_test.recov_alert.q &&
    reg2hw.alert_test.recov_alert.qe
  };
  assign fatal_alert_test_o = {
    reg2hw.alert_test.fatal_alert.q &&
    reg2hw.alert_test.fatal_alert.qe
  };


  assign recov_alert_event = cs_enable_pfa ||
         sw_app_enable_pfa ||
         read_int_state_pfa ||
         acmd_flag0_pfa ||
         cs_main_sm_alert ||
         cs_bus_cmp_alert;


  prim_edge_detector #(
    .Width(1),
    .ResetValue(0),
    .EnSync(0)
  ) u_prim_edge_detector_recov_alert (
    .clk_i,
    .rst_ni,
    .d_i(recov_alert_event),
    .q_sync_o(),
    .q_posedge_pulse_o(recov_alert_o),
    .q_negedge_pulse_o()
  );


  // check for illegal enable field states, and set alert if detected

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_cs_enable;
  assign mubi_cs_enable = mubi4_t'(reg2hw.ctrl.enable.q);
  assign cs_enable_pfa = mubi4_test_invalid(mubi_cs_enable_fanout[0]);
  assign hw2reg.recov_alert_sts.enable_field_alert.de = cs_enable_pfa;
  assign hw2reg.recov_alert_sts.enable_field_alert.d  = cs_enable_pfa;

  for (genvar i = 1; i < CsEnableCopies; i = i+1) begin : gen_mubi_en_copies
    assign cs_enable_fo[i] = mubi4_test_true_strict(mubi_cs_enable_fanout[i]);
  end : gen_mubi_en_copies

  prim_mubi4_sync #(
    .NumCopies(CsEnableCopies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_cs_enable (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_cs_enable),
    .mubi_o(mubi_cs_enable_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_sw_app_enable;
  mubi4_t [1:0] mubi_sw_app_enable_fanout;
  assign mubi_sw_app_enable = mubi4_t'(reg2hw.ctrl.sw_app_enable.q);
  assign sw_app_enable_pfe = mubi4_test_true_strict(mubi_sw_app_enable_fanout[0]);
  assign sw_app_enable_pfa = mubi4_test_invalid(mubi_sw_app_enable_fanout[1]);
  assign hw2reg.recov_alert_sts.sw_app_enable_field_alert.de = sw_app_enable_pfa;
  assign hw2reg.recov_alert_sts.sw_app_enable_field_alert.d  = sw_app_enable_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_sw_app_enable (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_sw_app_enable),
    .mubi_o(mubi_sw_app_enable_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_read_int_state;
  mubi4_t [1:0] mubi_read_int_state_fanout;
  assign mubi_read_int_state = mubi4_t'(reg2hw.ctrl.read_int_state.q);
  assign read_int_state_pfe = mubi4_test_true_strict(mubi_read_int_state_fanout[0]);
  assign read_int_state_pfa = mubi4_test_invalid(mubi_read_int_state_fanout[1]);
  assign hw2reg.recov_alert_sts.read_int_state_field_alert.de = read_int_state_pfa;
  assign hw2reg.recov_alert_sts.read_int_state_field_alert.d  = read_int_state_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_read_int_state (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_read_int_state),
    .mubi_o(mubi_read_int_state_fanout)
  );


  // master module enable
  assign sw_app_enable = sw_app_enable_pfe;
  assign read_int_state = read_int_state_pfe;

  //------------------------------------------
  // application interface
  //------------------------------------------
  // Each application port has its own
  // csrng_cmd_stage block to recieve the
  // command, track the state of its completion,
  // and return any genbits if the command
  // is a generate command.

  for (genvar ai = 0; ai < NApps; ai = ai+1) begin : gen_cmd_stage

    csrng_cmd_stage #(
      .CmdFifoWidth(AppCmdWidth),
      .CmdFifoDepth(AppCmdFifoDepth),
      .StateId(StateId)
    ) u_csrng_cmd_stage (
      .clk_i                        (clk_i),
      .rst_ni                       (rst_ni),
      .cs_enable_i                  (cs_enable_fo[27]),
      .cmd_stage_vld_i              (cmd_stage_vld[ai]),
      .cmd_stage_shid_i             (cmd_stage_shid[ai]),
      .cmd_stage_bus_i              (cmd_stage_bus[ai]),
      .cmd_stage_rdy_o              (cmd_stage_rdy[ai]),
      .cmd_arb_req_o                (cmd_arb_req[ai]),
      .cmd_arb_sop_o                (cmd_arb_sop[ai]),
      .cmd_arb_mop_o                (cmd_arb_mop[ai]),
      .cmd_arb_eop_o                (cmd_arb_eop[ai]),
      .cmd_arb_gnt_i                (cmd_arb_gnt[ai]),
      .cmd_arb_bus_o                (cmd_arb_bus[ai]),
      .cmd_ack_i                    (cmd_core_ack[ai]),
      .cmd_ack_sts_i                (cmd_core_ack_sts[ai]),
      .cmd_stage_ack_o              (cmd_stage_ack[ai]),
      .cmd_stage_ack_sts_o          (cmd_stage_ack_sts[ai]),
      .genbits_vld_i                (genbits_core_vld[ai]),
      .genbits_bus_i                (genbits_core_bus[ai]),
      .genbits_fips_i               (genbits_core_fips[ai]),
      .genbits_vld_o                (genbits_stage_vld[ai]),
      .genbits_rdy_i                (genbits_stage_rdy[ai]),
      .genbits_bus_o                (genbits_stage_bus[ai]),
      .genbits_fips_o               (genbits_stage_fips[ai]),
      .cmd_stage_sfifo_cmd_err_o    (cmd_stage_sfifo_cmd_err[ai]),
      .cmd_stage_sfifo_genbits_err_o(cmd_stage_sfifo_genbits_err[ai]),
      .cmd_gen_cnt_err_o            (cmd_gen_cnt_err[ai]),
      .cmd_stage_sm_err_o           (cmd_stage_sm_err[ai])
    );

  end : gen_cmd_stage

  // SW interface connection (only 1, and must be present)
  // cmd req
  assign cmd_stage_vld[NApps-1] = reg2hw.cmd_req.qe;
  assign cmd_stage_shid[NApps-1] = StateId'(NApps-1);
  assign cmd_stage_bus[NApps-1] = reg2hw.cmd_req.q;
  assign hw2reg.sw_cmd_sts.cmd_rdy.de = 1'b1;
  assign hw2reg.sw_cmd_sts.cmd_rdy.d = cmd_rdy;
  assign cmd_rdy = !cmd_stage_vld[NApps-1] && sw_rdy_sts_q;
  assign sw_rdy_sts_d =
         !cs_enable_fo[28] ? 1'b1 :
         cmd_stage_vld[NApps-1] ? 1'b0 :
         cmd_stage_rdy[NApps-1] ? 1'b1 :
         sw_rdy_sts_q;

  // cmd ack sts
  assign hw2reg.sw_cmd_sts.cmd_sts.de = cmd_stage_ack[NApps-1];
  assign hw2reg.sw_cmd_sts.cmd_sts.d = cmd_stage_ack_sts[NApps-1];
  // genbits
  assign hw2reg.genbits_vld.genbits_vld.d = genbits_stage_vldo_sw;
  assign hw2reg.genbits_vld.genbits_fips.d = genbits_stage_fips_sw;
  assign hw2reg.genbits.d = (sw_app_enable && efuse_sw_app_enable[0]) ? genbits_stage_bus_sw : '0;
  assign genbits_stage_bus_rd_sw = reg2hw.genbits.re;

  assign efuse_sw_app_enable[0] = prim_mubi_pkg::mubi8_test_true_strict(en_csrng_sw_app_read[0]);
  assign efuse_sw_app_enable[1] = prim_mubi_pkg::mubi8_test_true_strict(en_csrng_sw_app_read[1]);

  prim_mubi8_sync #(
    .NumCopies(2),
    .AsyncOn(1)
  ) u_prim_mubi8_sync_sw_app_read (
    .clk_i,
    .rst_ni,
    .mubi_i(otp_en_csrng_sw_app_read_i),
    .mubi_o(en_csrng_sw_app_read)
  );

  // pack the gen bits into a 32 bit register sized word

  prim_packer_fifo #(
    .InW(BlkLen),
    .OutW(32),
    .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_sw_genbits (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .clr_i    (!cs_enable_fo[29]),
    .wvalid_i (genbits_stage_vld[NApps-1]),
    .wdata_i  (genbits_stage_bus[NApps-1]),
    .wready_o (genbits_stage_rdy[NApps-1]),
    .rvalid_o (genbits_stage_vldo_sw),
    .rdata_o  (genbits_stage_bus_sw),
    .rready_i (genbits_stage_bus_rd_sw),
    .depth_o  ()
  );

  // flops for SW fips status
  assign genbits_stage_fips_sw_d =
         (!cs_enable_fo[30]) ? 1'b0 :
         (genbits_stage_rdy[NApps-1] && genbits_stage_vld[NApps-1]) ? genbits_stage_fips[NApps-1] :
         genbits_stage_fips_sw_q;

  assign genbits_stage_fips_sw = genbits_stage_fips_sw_q;


  //--------------------------------------------
  // data path integrity check
  // - a countermeasure to detect entropy bus tampering attempts
  // - checks to make sure repeated data sets off
  //   an alert for sw to handle
  //--------------------------------------------

  // SEC_CM: SW_GENBITS.BUS.CONSISTENCY

  // capture a copy of the genbits data
  assign cs_rdata_capt_vld = (genbits_stage_vld[NApps-1] && genbits_stage_rdy[NApps-1]);

  assign cs_rdata_capt_d = cs_rdata_capt_vld ? genbits_stage_bus[NApps-1][63:0] : cs_rdata_capt_q;

  assign cs_rdata_capt_vld_d =
         !cs_enable_fo[31] ? 1'b0 :
         cs_rdata_capt_vld ? 1'b1 :
         cs_rdata_capt_vld_q;

  // continuous compare of the entropy data for sw port
  assign cs_bus_cmp_alert = cs_rdata_capt_vld && cs_rdata_capt_vld_q &&
         (cs_rdata_capt_q == genbits_stage_bus[NApps-1][63:0]); // only look at 64 bits

  assign hw2reg.recov_alert_sts.cs_bus_cmp_alert.de = cs_bus_cmp_alert;
  assign hw2reg.recov_alert_sts.cs_bus_cmp_alert.d  = cs_bus_cmp_alert;

  assign hw2reg.recov_alert_sts.cs_main_sm_alert.de = cs_main_sm_alert;
  assign hw2reg.recov_alert_sts.cs_main_sm_alert.d  = cs_main_sm_alert;


  // HW interface connections (up to 16, numbered 0-14)
  for (genvar hai = 0; hai < (NApps-1); hai = hai+1) begin : gen_app_if
    // cmd req
    assign cmd_stage_vld[hai] = csrng_cmd_i[hai].csrng_req_valid;
    assign cmd_stage_shid[hai] = hai;
    assign cmd_stage_bus[hai] = csrng_cmd_i[hai].csrng_req_bus;
    assign csrng_cmd_o[hai].csrng_req_ready = cmd_stage_rdy[hai];
    // cmd ack
    assign csrng_cmd_o[hai].csrng_rsp_ack = cmd_stage_ack[hai];
    assign csrng_cmd_o[hai].csrng_rsp_sts = cmd_stage_ack_sts[hai];
    // genbits
    assign csrng_cmd_o[hai].genbits_valid = genbits_stage_vld[hai];
    assign csrng_cmd_o[hai].genbits_fips = genbits_stage_fips[hai];
    assign csrng_cmd_o[hai].genbits_bus = genbits_stage_bus[hai];
    assign genbits_stage_rdy[hai] = csrng_cmd_i[hai].genbits_ready;
  end : gen_app_if

  // set ack status for configured instances
  for (genvar i = 0; i < NHwApps; i = i+1) begin : gen_app_if_sts
    assign hw_exception_sts[i] = cmd_stage_ack[i] && cmd_stage_ack_sts[i];
  end : gen_app_if_sts

  // set ack status to zero for un-configured instances
  for (genvar i = NHwApps; i < 16; i = i+1) begin : gen_app_if_zero_sts
    assign hw_exception_sts[i] = 1'b0;
  end : gen_app_if_zero_sts

  // set fifo err status bits
  for (genvar i = 0; i < NApps; i = i+1) begin : gen_fifo_sts
    assign cmd_stage_sfifo_cmd_err_sum[i] = (|cmd_stage_sfifo_cmd_err[i] ||
                                             err_code_test_bit[0]);
    assign cmd_stage_sfifo_cmd_err_wr[i] = cmd_stage_sfifo_cmd_err[i][2];
    assign cmd_stage_sfifo_cmd_err_rd[i] = cmd_stage_sfifo_cmd_err[i][1];
    assign cmd_stage_sfifo_cmd_err_st[i] = cmd_stage_sfifo_cmd_err[i][0];
    assign cmd_stage_sfifo_genbits_err_sum[i] = (|cmd_stage_sfifo_genbits_err[i] ||
                                                 err_code_test_bit[1]);
    assign cmd_stage_sfifo_genbits_err_wr[i] = cmd_stage_sfifo_genbits_err[i][2];
    assign cmd_stage_sfifo_genbits_err_rd[i] = cmd_stage_sfifo_genbits_err[i][1];
    assign cmd_stage_sfifo_genbits_err_st[i] = cmd_stage_sfifo_genbits_err[i][0];
  end : gen_fifo_sts

  //------------------------------------------
  // app command arbiter and state machine
  //------------------------------------------
  // All commands that arrive from the
  // application ports are arbitrated for
  // and processed by the main state machine
  // logic block.

  assign cmd_arb_idx_d = (acmd_avail && acmd_accept) ? cmd_arb_idx : cmd_arb_idx_q;

  assign acmd_sop = cmd_arb_sop[cmd_arb_idx_q];
  assign acmd_mop = cmd_arb_mop[cmd_arb_idx_q];
  assign acmd_eop = cmd_arb_eop[cmd_arb_idx_q];
  assign acmd_bus = cmd_arb_bus[cmd_arb_idx_q];

  prim_arbiter_ppc #(
    .EnDataPort(0),    // Ignore data port
    .N(NApps),  // Number of request ports
    .DW(1), // Data width
    .IdxW($clog2(NApps))
  ) u_prim_arbiter_ppc_acmd (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .req_chk_i(cs_enable_fo[1]),
    .req_i    (cmd_arb_req),
    .data_i   ('{default: 1'b0}),
    .gnt_o    (cmd_arb_gnt),
    .idx_o    (cmd_arb_idx),
    .valid_o  (acmd_avail), // 1 req
    .data_o   (), //NC
    .ready_i  (acmd_accept) // 1 fsm rdy
  );

  mubi4_t mubi_acmd_flag0;
  assign mubi_acmd_flag0 = mubi4_t'(acmd_bus[11:8]);
  assign acmd_flag0_pfa = mubi4_test_invalid(flag0_q);
  assign hw2reg.recov_alert_sts.acmd_flag0_field_alert.de = acmd_flag0_pfa;
  assign hw2reg.recov_alert_sts.acmd_flag0_field_alert.d  = acmd_flag0_pfa;

  // parse the command bus
  assign acmd_hold = acmd_sop ? acmd_bus[2:0] : acmd_q;
  assign flag0 = mubi_acmd_flag0;
  assign shid = acmd_bus[15:12];
  assign gen_last = acmd_bus[16];

  assign acmd_d =
         (!cs_enable_fo[32]) ? '0 :
         acmd_sop ? acmd_bus[2:0] :
         acmd_q;

  assign shid_d =
         (!cs_enable_fo[33]) ? '0 :
         acmd_sop ? shid :
         shid_q;

  assign gen_last_d =
         (!cs_enable_fo[34]) ? '0 :
         acmd_sop ? gen_last :
         gen_last_q;

  assign flag0_d =
         (!cs_enable_fo[35]) ? prim_mubi_pkg::MuBi4False :
         (acmd_sop && ((acmd_bus[2:0] == INS) || (acmd_bus[2:0] == RES))) ? flag0 :
         flag0_q;

  // SEC_CM: CTRL.MUBI
  mubi4_t mubi_flag0;
  assign mubi_flag0 = flag0_q;

  for (genvar i = 0; i < Flag0Copies; i = i+1) begin : gen_mubi_flag0_copies
    assign flag0_fo[i] = mubi4_test_true_strict(mubi_flag0_fanout[i]);
  end : gen_mubi_flag0_copies

  prim_mubi4_sync #(
    .NumCopies(Flag0Copies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_flag0 (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_flag0),
    .mubi_o(mubi_flag0_fanout)
  );

  // sm to process all instantiation requests
  // SEC_CM: MAIN_SM.CTR.LOCAL_ESC
  // SEC_CM: MAIN_SM.FSM.SPARSE
  csrng_main_sm u_csrng_main_sm (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .enable_i               (cs_enable_fo[36]),
    .acmd_avail_i           (acmd_avail),
    .acmd_accept_o          (acmd_accept),
    .acmd_i                 (acmd_hold),
    .acmd_eop_i             (acmd_eop),
    .ctr_drbg_cmd_req_rdy_i (ctr_drbg_cmd_req_rdy),
    .flag0_i                (flag0_fo[0]),
    .cmd_entropy_req_o      (cmd_entropy_req),
    .cmd_entropy_avail_i    (cmd_entropy_avail),
    .instant_req_o          (instant_req),
    .reseed_req_o           (reseed_req),
    .generate_req_o         (generate_req),
    .update_req_o           (update_req),
    .uninstant_req_o        (uninstant_req),
    .clr_adata_packer_o     (clr_adata_packer),
    .cmd_complete_i         (state_db_wr_req),
    .local_escalate_i       (cmd_gen_cnt_err_sum),
    .main_sm_state_o        (cs_main_sm_state),
    .main_sm_alert_o        (cs_main_sm_alert),
    .main_sm_err_o          (cs_main_sm_err)
  );

  // interrupt for sw app interface only
  assign event_cs_cmd_req_done = cmd_stage_ack[NApps-1];

  // interrupt for entropy request
  assign event_cs_entropy_req = entropy_src_hw_if_o.es_req;

  // interrupt for app interface exception
  assign event_cs_hw_inst_exc = |hw_exception_sts;

  // entropy available
  assign cmd_entropy_avail = entropy_src_hw_if_i.es_ack;

  for (genvar csi = 0; csi < NApps; csi = csi+1) begin : gen_cmd_ack
    assign cmd_core_ack[csi] = state_db_sts_ack && (state_db_sts_id == csi);
    assign cmd_core_ack_sts[csi] = state_db_sts_sts;
    assign genbits_core_vld[csi] = gen_result_wr_req && (gen_result_inst_id == csi);
    assign genbits_core_bus[csi] = gen_result_bits;
    assign genbits_core_fips[csi] = gen_result_fips;
  end : gen_cmd_ack


  prim_packer_fifo #(
    .InW(32),
    .OutW(SeedLen),
    .ClearOnRead(1'b1)
  ) u_prim_packer_fifo_adata (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (!cs_enable_fo[37] || packer_adata_clr),
    .wvalid_i   (acmd_mop),
    .wdata_i    (acmd_bus),
    .wready_o   (),
    .rvalid_o   (),
    .rdata_o    (packer_adata),
    .rready_i   (packer_adata_pop),
    .depth_o    (packer_adata_depth)
  );

  assign packer_adata_pop = cs_enable_fo[38] &&
         clr_adata_packer && (packer_adata_depth == ADataDepthClog'(MaxClen));

  assign packer_adata_clr = cs_enable_fo[39] &&
         clr_adata_packer && (packer_adata_depth < ADataDepthClog'(MaxClen));

  //-------------------------------------
  // csrng_state_db nstantiation
  //-------------------------------------
  // This block holds the internal state
  // of each csrng instance. The state
  // is updated after each command.

  assign cmd_result_wr_req = cmd_result_ack && (cmd_result_ccmd != GEN);

  // register read access
  assign state_db_reg_rd_sel = reg2hw.int_state_val.re;
  assign state_db_reg_rd_id = reg2hw.int_state_num.q;
  assign state_db_reg_rd_id_pulse = reg2hw.int_state_num.qe;
  assign hw2reg.int_state_val.d = state_db_reg_rd_val;
  assign state_db_is_dump_en = cs_enable_fo[40] && read_int_state && efuse_sw_app_enable[1];


  csrng_state_db #(
    .NApps(NApps),
    .StateId(StateId),
    .BlkLen(BlkLen),
    .KeyLen(KeyLen),
    .CtrLen(CtrLen),
    .Cmd(Cmd)
  ) u_csrng_state_db (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .state_db_enable_i(cs_enable_fo[41]),
    .state_db_rd_inst_id_i(shid_q),
    .state_db_rd_key_o(state_db_rd_key),
    .state_db_rd_v_o(state_db_rd_v),
    .state_db_rd_res_ctr_o(state_db_rd_rc),
    .state_db_rd_inst_st_o(), // NC
    .state_db_rd_fips_o(state_db_rd_fips),

    .state_db_wr_req_i(state_db_wr_req),
    .state_db_wr_req_rdy_o(state_db_wr_req_rdy),
    .state_db_wr_inst_id_i(state_db_wr_inst_id),
    .state_db_wr_fips_i(state_db_wr_fips),
    .state_db_wr_ccmd_i(state_db_wr_ccmd),
    .state_db_wr_key_i(state_db_wr_key),
    .state_db_wr_v_i(state_db_wr_v),
    .state_db_wr_res_ctr_i(state_db_wr_rc),
    .state_db_wr_sts_i(state_db_wr_sts),

    .state_db_is_dump_en_i(state_db_is_dump_en),
    .state_db_reg_rd_sel_i(state_db_reg_rd_sel),
    .state_db_reg_rd_id_pulse_i(state_db_reg_rd_id_pulse),
    .state_db_reg_rd_id_i(state_db_reg_rd_id),
    .state_db_reg_rd_val_o(state_db_reg_rd_val),
    .state_db_sts_ack_o(state_db_sts_ack),
    .state_db_sts_sts_o(state_db_sts_sts),
    .state_db_sts_id_o(state_db_sts_id)
  );

  assign statedb_wr_select_d =
         (!cs_enable_fo[42]) ? '0 :
         !statedb_wr_select_q;

  assign cmd_blk_select = !statedb_wr_select_q;
  assign gen_blk_select =  statedb_wr_select_q;

  // return to requesting block
  assign cmd_result_ack_rdy = (cmd_blk_select && state_db_wr_req_rdy) && ctr_drbg_gen_req_rdy;
  assign gen_result_ack_rdy = gen_blk_select && state_db_wr_req_rdy;

  // muxes for statedb block inputs
  assign state_db_wr_req = gen_blk_select ? gen_result_wr_req : cmd_result_wr_req;
  assign state_db_wr_inst_id = gen_blk_select ? gen_result_inst_id : cmd_result_inst_id;
  assign state_db_wr_fips = gen_blk_select ? gen_result_fips : cmd_result_fips;
  assign state_db_wr_ccmd = gen_blk_select ?  gen_result_ccmd : cmd_result_ccmd;
  assign state_db_wr_key = gen_blk_select ? gen_result_key : cmd_result_key;
  assign state_db_wr_v = gen_blk_select ? gen_result_v : cmd_result_v;
  assign state_db_wr_rc = gen_blk_select ? gen_result_rc : cmd_result_rc;
  assign state_db_wr_sts = gen_blk_select ? gen_result_ack_sts : cmd_result_ack_sts;


  //--------------------------------------------
  // entropy interface
  //--------------------------------------------
  // Basic interface logic with the entropy_src block

  assign entropy_src_hw_if_o.es_req = cs_enable_fo[43] &&
         cmd_entropy_req;


  // SEC_CM: CONSTANTS.LC_GATED
  assign seed_diversification = lc_hw_debug_on_fo[0] ? RndCnstCsKeymgrDivNonProduction :
                                                       RndCnstCsKeymgrDivProduction;

  // Capture entropy from entropy_src
  assign entropy_src_seed_d =
         flag0_fo[1] ? '0 : // special case where zero is used
         cmd_entropy_req && cmd_entropy_avail ?
            (entropy_src_hw_if_i.es_bits ^ seed_diversification) :
         entropy_src_seed_q;
  assign entropy_src_fips_d =
         flag0_fo[2] ? '0 : // special case where zero is used
         cmd_entropy_req && cmd_entropy_avail ? entropy_src_hw_if_i.es_fips :
         entropy_src_fips_q;

  assign cmd_entropy = entropy_src_seed_q;

  assign cmd_entropy_fips = entropy_src_fips_q;

  //-------------------------------------
  // csrng_ctr_drbg_cmd instantiation
  //-------------------------------------
  // commands and input parameters
  // ins -> send to csrng_state_db
  //  inputs:  384b entropy, 384b adata
  //  outputs: 416b K,V,RC
  //
  // res -> send to csrng_state_db
  //  inputs:  416b K,V,RC, 384b entropy, 384b adata
  //  outputs: 416b K,V,RC
  //
  // gen -> send to csrng_ctr_drbg_gen block
  //  inputs:  416b K,V,RC, 384b adata
  //  outputs: 416b K,V,RC, 384b adata
  //
  // gen blk -> send to csrng_state_db
  //  inputs:  416b K,V,RC, 384b adata
  //  outputs: 416b K,V,RC, 128b genbits
  //
  // upd -> send to csrng_state_db
  //  inputs:  416b K,V,RC, 384b adata
  //  outputs: 416b K,V,RC



  assign cmd_req_ccmd_dly_d =
         (!cs_enable_fo[44]) ? '0 :
         acmd_hold;

  assign ctr_drbg_cmd_ccmd = cmd_req_ccmd_dly_q;


  assign cmd_req_dly_d =
         (!cs_enable_fo[45]) ? '0 :
         (instant_req || reseed_req || generate_req || update_req || uninstant_req);

  assign ctr_drbg_cmd_req = cmd_req_dly_q;

  csrng_ctr_drbg_cmd #(
    .Cmd(Cmd),
    .StateId(StateId),
    .BlkLen(BlkLen),
    .KeyLen(KeyLen),
    .SeedLen(SeedLen),
    .CtrLen(CtrLen)
  ) u_csrng_ctr_drbg_cmd (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .ctr_drbg_cmd_enable_i(cs_enable_fo[46]),
    .ctr_drbg_cmd_req_i(ctr_drbg_cmd_req),
    .ctr_drbg_cmd_rdy_o(ctr_drbg_cmd_req_rdy),
    .ctr_drbg_cmd_ccmd_i(ctr_drbg_cmd_ccmd),
    .ctr_drbg_cmd_inst_id_i(shid_q),
    .ctr_drbg_cmd_glast_i(gen_last_q),
    .ctr_drbg_cmd_entropy_i(cmd_entropy),
    .ctr_drbg_cmd_entropy_fips_i(cmd_entropy_fips), // send to state_db
    .ctr_drbg_cmd_adata_i(packer_adata),
    .ctr_drbg_cmd_key_i(state_db_rd_key),
    .ctr_drbg_cmd_v_i(state_db_rd_v),
    .ctr_drbg_cmd_rc_i(state_db_rd_rc),
    .ctr_drbg_cmd_fips_i(state_db_rd_fips), // send to genbits user

    .ctr_drbg_cmd_ack_o(cmd_result_ack),
    .ctr_drbg_cmd_sts_o(cmd_result_ack_sts),
    .ctr_drbg_cmd_rdy_i(cmd_result_ack_rdy),
    .ctr_drbg_cmd_ccmd_o(cmd_result_ccmd),
    .ctr_drbg_cmd_inst_id_o(cmd_result_inst_id),
    .ctr_drbg_cmd_glast_o(cmd_result_glast),
    .ctr_drbg_cmd_fips_o(cmd_result_fips),
    .ctr_drbg_cmd_adata_o(cmd_result_adata),
    .ctr_drbg_cmd_key_o(cmd_result_key),
    .ctr_drbg_cmd_v_o(cmd_result_v),
    .ctr_drbg_cmd_rc_o(cmd_result_rc),

    // interface to updblk from cmdblk
    .cmd_upd_req_o(cmdblk_updblk_arb_req),
    .upd_cmd_rdy_i(updblk_cmdblk_arb_req_rdy),
    .cmd_upd_ccmd_o(cmdblk_updblk_ccmd_arb_din),
    .cmd_upd_inst_id_o(cmdblk_updblk_id_arb_din),
    .cmd_upd_pdata_o(cmdblk_updblk_pdata_arb_din),
    .cmd_upd_key_o(cmdblk_updblk_key_arb_din),
    .cmd_upd_v_o(cmdblk_updblk_v_arb_din),

    .upd_cmd_ack_i(updblk_cmdblk_ack),
    .cmd_upd_rdy_o(cmdblk_updblk_ack_rdy),
    .upd_cmd_ccmd_i(updblk_ccmd),
    .upd_cmd_inst_id_i(updblk_inst_id),
    .upd_cmd_key_i(updblk_key),
    .upd_cmd_v_i(updblk_v),

    .ctr_drbg_cmd_sfifo_cmdreq_err_o(ctr_drbg_cmd_sfifo_cmdreq_err),
    .ctr_drbg_cmd_sfifo_rcstage_err_o(ctr_drbg_cmd_sfifo_rcstage_err),
    .ctr_drbg_cmd_sfifo_keyvrc_err_o(ctr_drbg_cmd_sfifo_keyvrc_err)
  );


  //-------------------------------------
  // csrng_ctr_drbg_upd instantiation
  //-------------------------------------
  // The csrng_ctr_drbg_upd is shared
  // between the csrng_ctr_drbg_cmd block
  // and the csrng_ctr_drbg_gen block.
  // The arbiter in this section will
  // route requests and responses between
  // these two blocks.


  csrng_ctr_drbg_upd #(
    .Cmd(Cmd),
    .StateId(StateId),
    .BlkLen(BlkLen),
    .KeyLen(KeyLen),
    .SeedLen(SeedLen),
    .CtrLen(CtrLen)
  ) u_csrng_ctr_drbg_upd (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .ctr_drbg_upd_enable_i(cs_enable_fo[47]),
    .ctr_drbg_upd_req_i(updblk_arb_vld),
    .ctr_drbg_upd_rdy_o(updblk_arb_rdy),
    .ctr_drbg_upd_ack_o(updblk_ack),
    .ctr_drbg_upd_rdy_i(updblk_ack_rdy),
    .ctr_drbg_upd_ccmd_i(updblk_arb_ccmd),
    .ctr_drbg_upd_inst_id_i(updblk_arb_inst_id),
    .ctr_drbg_upd_pdata_i(updblk_arb_pdata),
    .ctr_drbg_upd_key_i(updblk_arb_key),
    .ctr_drbg_upd_v_i(updblk_arb_v),
    .ctr_drbg_upd_ccmd_o(updblk_ccmd),
    .ctr_drbg_upd_inst_id_o(updblk_inst_id),
    .ctr_drbg_upd_key_o(updblk_key),
    .ctr_drbg_upd_v_o(updblk_v),

    // es halt interface
    .ctr_drbg_upd_es_req_i(cs_aes_halt_i.cs_aes_halt_req),
    .ctr_drbg_upd_es_ack_o(ctr_drbg_upd_es_ack),

    .block_encrypt_req_o(updblk_benblk_arb_req),
    .block_encrypt_rdy_i(updblk_benblk_arb_req_rdy),
    .block_encrypt_ccmd_o(updblk_benblk_cmd_arb_din),
    .block_encrypt_inst_id_o(updblk_benblk_id_arb_din),
    .block_encrypt_key_o(updblk_benblk_key_arb_din),
    .block_encrypt_v_o(updblk_benblk_v_arb_din),
    .block_encrypt_ack_i(benblk_updblk_ack),
    .block_encrypt_rdy_o(updblk_benblk_ack_rdy),
    .block_encrypt_ccmd_i(benblk_cmd),
    .block_encrypt_inst_id_i(benblk_inst_id),
    .block_encrypt_v_i(benblk_v),
    .ctr_drbg_upd_v_ctr_err_o(ctr_drbg_upd_v_ctr_err),
    .ctr_drbg_upd_sfifo_updreq_err_o(ctr_drbg_upd_sfifo_updreq_err),
    .ctr_drbg_upd_sfifo_bencreq_err_o(ctr_drbg_upd_sfifo_bencreq_err),
    .ctr_drbg_upd_sfifo_bencack_err_o(ctr_drbg_upd_sfifo_bencack_err),
    .ctr_drbg_upd_sfifo_pdata_err_o(ctr_drbg_upd_sfifo_pdata_err),
    .ctr_drbg_upd_sfifo_final_err_o(ctr_drbg_upd_sfifo_final_err),
    .ctr_drbg_updbe_sm_err_o(drbg_updbe_sm_err),
    .ctr_drbg_updob_sm_err_o(drbg_updob_sm_err)
  );

  // update block  arbiter

  prim_arbiter_ppc #(
    .N(NUpdateArbReqs), // (cmd req and gen req)
    .DW(UpdateArbWidth) // Data width
  ) u_prim_arbiter_ppc_updblk_arb (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .req_chk_i(cs_enable_fo[1]),
    .req_i({genblk_updblk_arb_req,cmdblk_updblk_arb_req}),
    .data_i(updblk_arb_din),
    .gnt_o({updblk_genblk_arb_req_rdy,updblk_cmdblk_arb_req_rdy}),
    .idx_o(),
    .valid_o(updblk_arb_vld),
    .data_o(updblk_arb_data),
    .ready_i(updblk_arb_rdy)
  );

  assign updblk_arb_din[0] = {cmdblk_updblk_key_arb_din,cmdblk_updblk_v_arb_din,
                              cmdblk_updblk_pdata_arb_din,
                              cmdblk_updblk_id_arb_din,cmdblk_updblk_ccmd_arb_din};

  assign updblk_arb_din[1] = {genblk_updblk_key_arb_din,genblk_updblk_v_arb_din,
                              genblk_updblk_pdata_arb_din,
                              genblk_updblk_id_arb_din,genblk_updblk_ccmd_arb_din};

  assign {updblk_arb_key,updblk_arb_v,updblk_arb_pdata,
          updblk_arb_inst_id,updblk_arb_ccmd} = updblk_arb_data;

  assign updblk_cmdblk_ack = (updblk_ack && (updblk_ccmd != GENU));
  assign updblk_genblk_ack = (updblk_ack && (updblk_ccmd == GENU));

  assign updblk_ack_rdy = (updblk_ccmd == GENU) ? genblk_updblk_ack_rdy : cmdblk_updblk_ack_rdy;


  //-------------------------------------
  // life cycle logic
  //-------------------------------------
  // The chip level life cycle control
  // provide control logic to determine
  // how certain debug features are controlled.

  lc_ctrl_pkg::lc_tx_t [LcHwDebugCopies-1:0] lc_hw_debug_en_out;

  prim_lc_sync #(
    .NumCopies(LcHwDebugCopies)
  ) u_prim_lc_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i(lc_hw_debug_en_i),
    .lc_en_o({lc_hw_debug_en_out})
  );

  for (genvar i = 0; i < LcHwDebugCopies; i = i+1) begin : gen_lc_dbg_copies
    assign lc_hw_debug_on_fo[i] = (lc_hw_debug_en_out[i] == lc_ctrl_pkg::On);
  end : gen_lc_dbg_copies


  //-------------------------------------
  // csrng_block_encrypt instantiation
  //-------------------------------------
  // The csrng_block_encrypt is shared
  // between the csrng_ctr_drbg_cmd block
  // and the csrng_ctr_drbg_gen block.
  // The arbiter in this section will
  // route requests and responses between
  // these two blocks.

  csrng_block_encrypt #(
    .SBoxImpl(SBoxImpl),
    .Cmd(Cmd),
    .StateId(StateId),
    .BlkLen(BlkLen),
    .KeyLen(KeyLen)
  ) u_csrng_block_encrypt (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .block_encrypt_enable_i(cs_enable_fo[48]),
    .block_encrypt_req_i(benblk_arb_vld),
    .block_encrypt_rdy_o(benblk_arb_rdy),
    .block_encrypt_key_i(benblk_arb_key),
    .block_encrypt_v_i(benblk_arb_v),
    .block_encrypt_cmd_i(benblk_arb_cmd),
    .block_encrypt_id_i(benblk_arb_inst_id),
    .block_encrypt_ack_o(benblk_ack),
    .block_encrypt_rdy_i(benblk_ack_rdy),
    .block_encrypt_cmd_o(benblk_cmd),
    .block_encrypt_id_o(benblk_inst_id),
    .block_encrypt_v_o(benblk_v),
    .block_encrypt_quiet_o(block_encrypt_quiet),
    .block_encrypt_aes_cipher_sm_err_o(aes_cipher_sm_err),
    .block_encrypt_sfifo_blkenc_err_o(block_encrypt_sfifo_blkenc_err)
  );


  prim_arbiter_ppc #(
    .N(NBlkEncArbReqs), // (upd req and gen req)
    .DW(BlkEncArbWidth) // Data width
  ) u_prim_arbiter_ppc_benblk_arb (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .req_chk_i(cs_enable_fo[1]),
    .req_i({genblk_benblk_arb_req,updblk_benblk_arb_req}),
    .data_i(benblk_arb_din),
    .gnt_o({genblk_benblk_arb_req_rdy,updblk_benblk_arb_req_rdy}),
    .idx_o(),
    .valid_o(benblk_arb_vld),
    .data_o(benblk_arb_data),
    .ready_i(benblk_arb_rdy)
  );

  assign benblk_arb_din[0] = {updblk_benblk_key_arb_din,updblk_benblk_v_arb_din,
                              updblk_benblk_id_arb_din,updblk_benblk_cmd_arb_din};
  assign benblk_arb_din[1] = {genblk_benblk_key_arb_din,genblk_benblk_v_arb_din,
                              genblk_benblk_id_arb_din,genblk_benblk_cmd_arb_din};

  assign benblk_updblk_ack = (benblk_ack && (benblk_cmd != GENB));
  assign benblk_genblk_ack = (benblk_ack && (benblk_cmd == GENB));

  assign benblk_ack_rdy = (benblk_cmd == GENB) ? genblk_benblk_ack_rdy : updblk_benblk_ack_rdy;

  assign {benblk_arb_key,benblk_arb_v,benblk_arb_inst_id,benblk_arb_cmd} = benblk_arb_data;


  //-------------------------------------
  // csrng_ctr_drbg_gen instantiation
  //-------------------------------------
  // this block performs the second sequence
  // of the generate command. The first part
  // of the sequence is done by the
  // csrng_ctr_drbg_cmd block.

  assign ctr_drbg_gen_req = cmd_result_ack && (cmd_result_ccmd == GEN);


  csrng_ctr_drbg_gen #(
    .NApps(NApps),
    .Cmd(Cmd),
    .StateId(StateId),
    .BlkLen(BlkLen),
    .KeyLen(KeyLen),
    .SeedLen(SeedLen),
    .CtrLen(CtrLen)
  ) u_csrng_ctr_drbg_gen (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .ctr_drbg_gen_enable_i(cs_enable_fo[49]),
    .ctr_drbg_gen_req_i(ctr_drbg_gen_req),
    .ctr_drbg_gen_rdy_o(ctr_drbg_gen_req_rdy),
    .ctr_drbg_gen_ccmd_i(cmd_result_ccmd),
    .ctr_drbg_gen_inst_id_i(cmd_result_inst_id),
    .ctr_drbg_gen_glast_i(cmd_result_glast),
    .ctr_drbg_gen_fips_i(cmd_result_fips),
    .ctr_drbg_gen_adata_i(cmd_result_adata),
    .ctr_drbg_gen_key_i(cmd_result_key),
    .ctr_drbg_gen_v_i(cmd_result_v),
    .ctr_drbg_gen_rc_i(cmd_result_rc),

    .ctr_drbg_gen_ack_o(gen_result_wr_req),
    .ctr_drbg_gen_sts_o(gen_result_ack_sts),
    .ctr_drbg_gen_rdy_i(gen_result_ack_rdy),
    .ctr_drbg_gen_ccmd_o(gen_result_ccmd),
    .ctr_drbg_gen_inst_id_o(gen_result_inst_id),
    .ctr_drbg_gen_fips_o(gen_result_fips),
    .ctr_drbg_gen_key_o(gen_result_key),
    .ctr_drbg_gen_v_o(gen_result_v),
    .ctr_drbg_gen_rc_o(gen_result_rc),
    .ctr_drbg_gen_bits_o(gen_result_bits),

    // es halt interface
    .ctr_drbg_gen_es_req_i(cs_aes_halt_i.cs_aes_halt_req),
    .ctr_drbg_gen_es_ack_o(ctr_drbg_gen_es_ack),

    // interface to updblk from genblk
    .gen_upd_req_o(genblk_updblk_arb_req),
    .upd_gen_rdy_i(updblk_genblk_arb_req_rdy),
    .gen_upd_ccmd_o(genblk_updblk_ccmd_arb_din),
    .gen_upd_inst_id_o(genblk_updblk_id_arb_din),
    .gen_upd_pdata_o(genblk_updblk_pdata_arb_din),
    .gen_upd_key_o(genblk_updblk_key_arb_din),
    .gen_upd_v_o(genblk_updblk_v_arb_din),

    .upd_gen_ack_i(updblk_genblk_ack),
    .gen_upd_rdy_o(genblk_updblk_ack_rdy),
    .upd_gen_ccmd_i(updblk_ccmd),
    .upd_gen_inst_id_i(updblk_inst_id),
    .upd_gen_key_i(updblk_key),
    .upd_gen_v_i(updblk_v),

    .block_encrypt_req_o(genblk_benblk_arb_req),
    .block_encrypt_rdy_i(genblk_benblk_arb_req_rdy),
    .block_encrypt_ccmd_o(genblk_benblk_cmd_arb_din),
    .block_encrypt_inst_id_o(genblk_benblk_id_arb_din),
    .block_encrypt_key_o(genblk_benblk_key_arb_din),
    .block_encrypt_v_o(genblk_benblk_v_arb_din),
    .block_encrypt_ack_i(benblk_genblk_ack),
    .block_encrypt_rdy_o(genblk_benblk_ack_rdy),
    .block_encrypt_ccmd_i(benblk_cmd),
    .block_encrypt_inst_id_i(benblk_inst_id),
    .block_encrypt_v_i(benblk_v),

    .ctr_drbg_gen_v_ctr_err_o(ctr_drbg_gen_v_ctr_err),
    .ctr_drbg_gen_sfifo_gbencack_err_o(ctr_drbg_gen_sfifo_gbencack_err),
    .ctr_drbg_gen_sfifo_grcstage_err_o(ctr_drbg_gen_sfifo_grcstage_err),
    .ctr_drbg_gen_sfifo_ggenreq_err_o(ctr_drbg_gen_sfifo_ggenreq_err),
    .ctr_drbg_gen_sfifo_gadstage_err_o(ctr_drbg_gen_sfifo_gadstage_err),
    .ctr_drbg_gen_sfifo_ggenbits_err_o(ctr_drbg_gen_sfifo_ggenbits_err),
    .ctr_drbg_gen_sm_err_o(drbg_gen_sm_err)
  );


  // es to cs halt request to reduce power spikes
  assign cs_aes_halt_d =
         (ctr_drbg_upd_es_ack && ctr_drbg_gen_es_ack && block_encrypt_quiet &&
          cs_aes_halt_i.cs_aes_halt_req);

  assign cs_aes_halt_o.cs_aes_halt_ack = cs_aes_halt_q;

  //--------------------------------------------
  // observe state machine
  //--------------------------------------------

  assign hw2reg.main_sm_state.de = 1'b1;
  assign hw2reg.main_sm_state.d = cs_main_sm_state;

  //--------------------------------------------
  // report csrng request summary
  //--------------------------------------------
  // Misc status

  assign hw2reg.hw_exc_sts.de = cs_enable_fo[50];
  assign hw2reg.hw_exc_sts.d  = hw_exception_sts;

  // unused signals
  assign unused_err_code_test_bit = (|err_code_test_bit[19:16]) || (|err_code_test_bit[27:26]);
  assign unused_reg2hw_genbits = (|reg2hw.genbits.q);
  assign unused_int_state_val = (|reg2hw.int_state_val.q);

  //--------------------------------------------
  // Assertions
  //--------------------------------------------
`ifdef INC_ASSERT
  // Track activity of AES.
  logic aes_active_d, aes_active_q;
  assign aes_active_d =
      (u_csrng_block_encrypt.u_aes_cipher_core.in_valid_i == aes_pkg::SP2V_HIGH &&
       u_csrng_block_encrypt.u_aes_cipher_core.in_ready_o == aes_pkg::SP2V_HIGH)  ? 1'b1 : // set
      (u_csrng_block_encrypt.u_aes_cipher_core.out_valid_o == aes_pkg::SP2V_HIGH &&
       u_csrng_block_encrypt.u_aes_cipher_core.out_ready_i == aes_pkg::SP2V_HIGH) ? 1'b0 : // clear
      aes_active_q;                                                                        // keep

  // Track state of AES Halt req/ack with entropy_src.
  logic cs_aes_halt_active;
  assign cs_aes_halt_active = cs_aes_halt_i.cs_aes_halt_req & cs_aes_halt_o.cs_aes_halt_ack;

  // Assert that when AES Halt is active, AES is not active.
  `ASSERT(AesNotActiveWhileCsAesHaltActive_A, cs_aes_halt_active |-> !aes_active_d)

  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      aes_active_q <= '0;
    end else begin
      aes_active_q <= aes_active_d;
    end
  end
`endif

endmodule // csrng_core


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: csrng top level wrapper file

`include "prim_assert.sv"

module csrng
 import csrng_pkg::*;
 import csrng_reg_pkg::*;
#(
  parameter aes_pkg::sbox_impl_e SBoxImpl = aes_pkg::SBoxImplCanright,
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},
  parameter int NHwApps = 2,
  parameter cs_keymgr_div_t RndCnstCsKeymgrDivNonProduction = CsKeymgrDivWidth'(0),
  parameter cs_keymgr_div_t RndCnstCsKeymgrDivProduction = CsKeymgrDivWidth'(0)
) (
  input logic         clk_i,
  input logic         rst_ni,

  // Tilelink Bus Interface
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

   // OTP Interface
  // SEC_CM: INTERSIG.MUBI
  input  prim_mubi_pkg::mubi8_t otp_en_csrng_sw_app_read_i,

  // Lifecycle broadcast inputs
  input  lc_ctrl_pkg::lc_tx_t  lc_hw_debug_en_i,

  // Entropy Interface
  output entropy_src_pkg::entropy_src_hw_if_req_t entropy_src_hw_if_o,
  input  entropy_src_pkg::entropy_src_hw_if_rsp_t entropy_src_hw_if_i,

  // Entropy Interface
  input  entropy_src_pkg::cs_aes_halt_req_t cs_aes_halt_i,
  output entropy_src_pkg::cs_aes_halt_rsp_t cs_aes_halt_o,

  // Application Interfaces
  input  csrng_req_t  [NHwApps-1:0] csrng_cmd_i,
  output csrng_rsp_t  [NHwApps-1:0] csrng_cmd_o,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // Interrupts
  output logic    intr_cs_cmd_req_done_o,
  output logic    intr_cs_entropy_req_o,
  output logic    intr_cs_hw_inst_exc_o,
  output logic    intr_cs_fatal_err_o
);

  csrng_reg2hw_t reg2hw;
  csrng_hw2reg_t hw2reg;

  logic [NumAlerts-1:0] alert_test;
  logic [NumAlerts-1:0] alert;

  logic [NumAlerts-1:0] intg_err_alert;
  assign intg_err_alert[0] = 1'b0;

  // SEC_CM: CONFIG.REGWEN
  // SEC_CM: TILE_LINK.BUS.INTEGRITY

  csrng_reg_top u_reg (
    .clk_i,
    .rst_ni,
    .tl_i,
    .tl_o,
    .reg2hw,
    .hw2reg,
    .intg_err_o(intg_err_alert[1]),
    .devmode_i(1'b1)
  );

  csrng_core #(
    .SBoxImpl(SBoxImpl),
    .NHwApps(NHwApps),
    .RndCnstCsKeymgrDivNonProduction(RndCnstCsKeymgrDivNonProduction),
    .RndCnstCsKeymgrDivProduction(RndCnstCsKeymgrDivProduction)
  ) u_csrng_core (
    .clk_i,
    .rst_ni,
    .reg2hw,
    .hw2reg,

    // misc inputs
    .otp_en_csrng_sw_app_read_i(otp_en_csrng_sw_app_read_i),
    .lc_hw_debug_en_i,

    // Entropy Interface
    .entropy_src_hw_if_o,
    .entropy_src_hw_if_i,

    // Entropy Interface
    .cs_aes_halt_i,
    .cs_aes_halt_o,

    // Application Interfaces
    .csrng_cmd_i,
    .csrng_cmd_o,

    // Alerts
    .recov_alert_test_o(alert_test[0]),
    .fatal_alert_test_o(alert_test[1]),
    .recov_alert_o(alert[0]),
    .fatal_alert_o(alert[1]),

    .intr_cs_cmd_req_done_o,
    .intr_cs_entropy_req_o,
    .intr_cs_hw_inst_exc_o,
    .intr_cs_fatal_err_o
  );


  ///////////////////////////
  // Alert generation
  ///////////////////////////
  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i)
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i]                 ),
      .alert_req_i   ( alert[i] || intg_err_alert[i] ),
      .alert_ack_o   (                               ),
      .alert_state_o (                               ),
      .alert_rx_i    ( alert_rx_i[i]                 ),
      .alert_tx_o    ( alert_tx_o[i]                 )
    );
  end


  // Assertions

  `ASSERT_KNOWN(TlDValidKnownO_A, tl_o.d_valid)
  `ASSERT_KNOWN(TlAReadyKnownO_A, tl_o.a_ready)
  `ASSERT_KNOWN(EsReqKnownO_A, entropy_src_hw_if_o.es_req)

  // Application Interface Asserts
  for (genvar i = 0; i < NHwApps; i = i+1) begin : gen_app_if_asserts
    `ASSERT_KNOWN(CsrngReqReadyKnownO_A, csrng_cmd_o[i].csrng_req_ready)
    `ASSERT_KNOWN(CsrngRspAckKnownO_A, csrng_cmd_o[i].csrng_rsp_ack)
    `ASSERT_KNOWN(CsrngRspStsKnownO_A, csrng_cmd_o[i].csrng_rsp_sts)
    `ASSERT_KNOWN(CsrngGenbitsValidKnownO_A, csrng_cmd_o[i].genbits_valid)
    `ASSERT_KNOWN_IF(CsrngGenbitsFipsKnownO_A, csrng_cmd_o[i].genbits_fips,
        csrng_cmd_o[i].genbits_valid)
    `ASSERT_KNOWN_IF(CsrngGenbitsBusKnownO_A, csrng_cmd_o[i].genbits_bus,
        csrng_cmd_o[i].genbits_valid)
  end : gen_app_if_asserts

  // Alerts
  `ASSERT_KNOWN(AlertTxKnownO_A, alert_tx_o)

  `ASSERT_KNOWN(IntrCsCmdReqDoneKnownO_A, intr_cs_cmd_req_done_o)
  `ASSERT_KNOWN(IntrCsEntropyReqKnownO_A, intr_cs_entropy_req_o)
  `ASSERT_KNOWN(IntrCsHwInstExcKnownO_A, intr_cs_hw_inst_exc_o)
  `ASSERT_KNOWN(IntrCsFatalErrKnownO_A, intr_cs_fatal_err_o)

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CtrDrbgUpdAlertCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_upd.u_prim_count_ctr_drbg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CtrDrbgGenAlertCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_gen.u_prim_count_ctr_drbg,
    alert_tx_o[1])

  for (genvar i = 0; i < NHwApps + 1; i++) begin : gen_cnt_asserts
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck_A,
      u_csrng_core.gen_cmd_stage[i].u_csrng_cmd_stage.u_prim_count_cmd_gen_cntr,
      alert_tx_o[1])

    `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgCmdFsmCheck_A,
      u_csrng_core.gen_cmd_stage[i].u_csrng_cmd_stage.u_state_regs,
      alert_tx_o[1])
  end

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlMainFsmCheck_A,
    u_csrng_core.u_csrng_main_sm.u_state_regs,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgGenFsmCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_gen.u_state_regs,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgUpdBlkEncFsmCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_upd.u_blk_enc_state_regs,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(DrbgUpdOutBlkFsmCheck_A,
    u_csrng_core.u_csrng_ctr_drbg_upd.u_outblk_state_regs,
    alert_tx_o[1])

  for (genvar i = 0; i < aes_pkg::Sp2VWidth; i++) begin : gen_aes_cipher_control_fsm_svas
    if (aes_pkg::SP2V_LOGIC_HIGH[i] == 1'b1) begin : gen_aes_cipher_control_fsm_svas_p
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCipherControlFsmCheck_A,
          u_csrng_core.u_csrng_block_encrypt.u_aes_cipher_core.u_aes_cipher_control.gen_fsm[i].
              gen_fsm_p.u_aes_cipher_control_fsm_i.u_aes_cipher_control_fsm.u_state_regs,
          alert_tx_o[1])
    end else begin : gen_aes_cipher_control_fsm_svas_n
      `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(AesCipherControlFsmCheck_A,
          u_csrng_core.u_csrng_block_encrypt.u_aes_cipher_core.u_aes_cipher_control.gen_fsm[i].
              gen_fsm_n.u_aes_cipher_control_fsm_i.u_aes_cipher_control_fsm.u_state_regs,
          alert_tx_o[1])
    end
  end

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package entropy_src_reg_pkg;

  // Param list
  parameter int unsigned ObserveFifoDepth = 64;
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 8;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } es_entropy_valid;
    struct packed {
      logic        q;
    } es_health_test_failed;
    struct packed {
      logic        q;
    } es_observe_fifo_ready;
    struct packed {
      logic        q;
    } es_fatal_err;
  } entropy_src_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } es_entropy_valid;
    struct packed {
      logic        q;
    } es_health_test_failed;
    struct packed {
      logic        q;
    } es_observe_fifo_ready;
    struct packed {
      logic        q;
    } es_fatal_err;
  } entropy_src_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } es_entropy_valid;
    struct packed {
      logic        q;
      logic        qe;
    } es_health_test_failed;
    struct packed {
      logic        q;
      logic        qe;
    } es_observe_fifo_ready;
    struct packed {
      logic        q;
      logic        qe;
    } es_fatal_err;
  } entropy_src_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_alert;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_alert;
  } entropy_src_reg2hw_alert_test_reg_t;

  typedef struct packed {
    logic        q;
  } entropy_src_reg2hw_sw_regupd_reg_t;

  typedef struct packed {
    logic [3:0]  q;
  } entropy_src_reg2hw_module_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } fips_enable;
    struct packed {
      logic [3:0]  q;
    } entropy_data_reg_enable;
    struct packed {
      logic [3:0]  q;
    } threshold_scope;
    struct packed {
      logic [3:0]  q;
    } rng_bit_enable;
    struct packed {
      logic [1:0]  q;
    } rng_bit_sel;
  } entropy_src_reg2hw_conf_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } es_route;
    struct packed {
      logic [3:0]  q;
    } es_type;
  } entropy_src_reg2hw_entropy_control_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        re;
  } entropy_src_reg2hw_entropy_data_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
    } fips_window;
    struct packed {
      logic [15:0] q;
    } bypass_window;
  } entropy_src_reg2hw_health_test_windows_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_repcnt_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_repcnts_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_adaptp_hi_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_adaptp_lo_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_bucket_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_markov_hi_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_markov_lo_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_extht_hi_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
      logic        qe;
    } fips_thresh;
    struct packed {
      logic [15:0] q;
      logic        qe;
    } bypass_thresh;
  } entropy_src_reg2hw_extht_lo_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] q;
    } alert_threshold;
    struct packed {
      logic [15:0] q;
    } alert_threshold_inv;
  } entropy_src_reg2hw_alert_threshold_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  q;
    } fw_ov_mode;
    struct packed {
      logic [3:0]  q;
    } fw_ov_entropy_insert;
  } entropy_src_reg2hw_fw_ov_control_reg_t;

  typedef struct packed {
    logic [3:0]  q;
  } entropy_src_reg2hw_fw_ov_sha3_start_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        re;
  } entropy_src_reg2hw_fw_ov_rd_data_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } entropy_src_reg2hw_fw_ov_wr_data_reg_t;

  typedef struct packed {
    logic [6:0]  q;
  } entropy_src_reg2hw_observe_fifo_thresh_reg_t;

  typedef struct packed {
    logic [4:0]  q;
    logic        qe;
  } entropy_src_reg2hw_err_code_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } es_entropy_valid;
    struct packed {
      logic        d;
      logic        de;
    } es_health_test_failed;
    struct packed {
      logic        d;
      logic        de;
    } es_observe_fifo_ready;
    struct packed {
      logic        d;
      logic        de;
    } es_fatal_err;
  } entropy_src_hw2reg_intr_state_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } entropy_src_hw2reg_regwen_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_entropy_data_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_repcnt_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_repcnts_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_adaptp_hi_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_adaptp_lo_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_bucket_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_markov_hi_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_markov_lo_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_extht_hi_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_thresh;
    struct packed {
      logic [15:0] d;
    } bypass_thresh;
  } entropy_src_hw2reg_extht_lo_thresholds_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_repcnt_hi_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_repcnts_hi_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_adaptp_hi_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_adaptp_lo_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_extht_hi_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_extht_lo_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_bucket_hi_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_markov_hi_watermarks_reg_t;

  typedef struct packed {
    struct packed {
      logic [15:0] d;
    } fips_watermark;
    struct packed {
      logic [15:0] d;
    } bypass_watermark;
  } entropy_src_hw2reg_markov_lo_watermarks_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_repcnt_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_repcnts_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_adaptp_hi_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_adaptp_lo_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_bucket_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_markov_hi_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_markov_lo_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_extht_hi_total_fails_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_extht_lo_total_fails_reg_t;

  typedef struct packed {
    logic [15:0] d;
  } entropy_src_hw2reg_alert_summary_fail_counts_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  d;
    } repcnt_fail_count;
    struct packed {
      logic [3:0]  d;
    } adaptp_hi_fail_count;
    struct packed {
      logic [3:0]  d;
    } adaptp_lo_fail_count;
    struct packed {
      logic [3:0]  d;
    } bucket_fail_count;
    struct packed {
      logic [3:0]  d;
    } markov_hi_fail_count;
    struct packed {
      logic [3:0]  d;
    } markov_lo_fail_count;
    struct packed {
      logic [3:0]  d;
    } repcnts_fail_count;
  } entropy_src_hw2reg_alert_fail_counts_reg_t;

  typedef struct packed {
    struct packed {
      logic [3:0]  d;
    } extht_hi_fail_count;
    struct packed {
      logic [3:0]  d;
    } extht_lo_fail_count;
  } entropy_src_hw2reg_extht_fail_counts_reg_t;

  typedef struct packed {
    logic        d;
  } entropy_src_hw2reg_fw_ov_wr_fifo_full_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } entropy_src_hw2reg_fw_ov_rd_fifo_overflow_reg_t;

  typedef struct packed {
    logic [31:0] d;
  } entropy_src_hw2reg_fw_ov_rd_data_reg_t;

  typedef struct packed {
    logic [6:0]  d;
  } entropy_src_hw2reg_observe_fifo_depth_reg_t;

  typedef struct packed {
    struct packed {
      logic [2:0]  d;
    } entropy_fifo_depth;
    struct packed {
      logic [2:0]  d;
    } sha3_fsm;
    struct packed {
      logic        d;
    } sha3_block_pr;
    struct packed {
      logic        d;
    } sha3_squeezing;
    struct packed {
      logic        d;
    } sha3_absorbed;
    struct packed {
      logic        d;
    } sha3_err;
    struct packed {
      logic        d;
    } main_sm_idle;
    struct packed {
      logic        d;
    } main_sm_boot_done;
  } entropy_src_hw2reg_debug_status_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } fips_enable_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } entropy_data_reg_en_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } module_enable_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } threshold_scope_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } rng_bit_enable_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } fw_ov_sha3_start_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } fw_ov_mode_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } fw_ov_entropy_insert_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_route_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_type_field_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_main_sm_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_bus_cmp_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_thresh_cfg_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_fw_ov_wr_alert;
    struct packed {
      logic        d;
      logic        de;
    } es_fw_ov_disable_alert;
  } entropy_src_hw2reg_recov_alert_sts_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } sfifo_esrng_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_observe_err;
    struct packed {
      logic        d;
      logic        de;
    } sfifo_esfinal_err;
    struct packed {
      logic        d;
      logic        de;
    } es_ack_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } es_main_sm_err;
    struct packed {
      logic        d;
      logic        de;
    } es_cntr_err;
    struct packed {
      logic        d;
      logic        de;
    } sha3_state_err;
    struct packed {
      logic        d;
      logic        de;
    } sha3_rst_storage_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_write_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_read_err;
    struct packed {
      logic        d;
      logic        de;
    } fifo_state_err;
  } entropy_src_hw2reg_err_code_reg_t;

  typedef struct packed {
    logic [8:0]  d;
    logic        de;
  } entropy_src_hw2reg_main_sm_state_reg_t;

  // Register -> HW type
  typedef struct packed {
    entropy_src_reg2hw_intr_state_reg_t intr_state; // [544:541]
    entropy_src_reg2hw_intr_enable_reg_t intr_enable; // [540:537]
    entropy_src_reg2hw_intr_test_reg_t intr_test; // [536:529]
    entropy_src_reg2hw_alert_test_reg_t alert_test; // [528:525]
    entropy_src_reg2hw_sw_regupd_reg_t sw_regupd; // [524:524]
    entropy_src_reg2hw_module_enable_reg_t module_enable; // [523:520]
    entropy_src_reg2hw_conf_reg_t conf; // [519:502]
    entropy_src_reg2hw_entropy_control_reg_t entropy_control; // [501:494]
    entropy_src_reg2hw_entropy_data_reg_t entropy_data; // [493:461]
    entropy_src_reg2hw_health_test_windows_reg_t health_test_windows; // [460:429]
    entropy_src_reg2hw_repcnt_thresholds_reg_t repcnt_thresholds; // [428:395]
    entropy_src_reg2hw_repcnts_thresholds_reg_t repcnts_thresholds; // [394:361]
    entropy_src_reg2hw_adaptp_hi_thresholds_reg_t adaptp_hi_thresholds; // [360:327]
    entropy_src_reg2hw_adaptp_lo_thresholds_reg_t adaptp_lo_thresholds; // [326:293]
    entropy_src_reg2hw_bucket_thresholds_reg_t bucket_thresholds; // [292:259]
    entropy_src_reg2hw_markov_hi_thresholds_reg_t markov_hi_thresholds; // [258:225]
    entropy_src_reg2hw_markov_lo_thresholds_reg_t markov_lo_thresholds; // [224:191]
    entropy_src_reg2hw_extht_hi_thresholds_reg_t extht_hi_thresholds; // [190:157]
    entropy_src_reg2hw_extht_lo_thresholds_reg_t extht_lo_thresholds; // [156:123]
    entropy_src_reg2hw_alert_threshold_reg_t alert_threshold; // [122:91]
    entropy_src_reg2hw_fw_ov_control_reg_t fw_ov_control; // [90:83]
    entropy_src_reg2hw_fw_ov_sha3_start_reg_t fw_ov_sha3_start; // [82:79]
    entropy_src_reg2hw_fw_ov_rd_data_reg_t fw_ov_rd_data; // [78:46]
    entropy_src_reg2hw_fw_ov_wr_data_reg_t fw_ov_wr_data; // [45:13]
    entropy_src_reg2hw_observe_fifo_thresh_reg_t observe_fifo_thresh; // [12:6]
    entropy_src_reg2hw_err_code_test_reg_t err_code_test; // [5:0]
  } entropy_src_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    entropy_src_hw2reg_intr_state_reg_t intr_state; // [1073:1066]
    entropy_src_hw2reg_regwen_reg_t regwen; // [1065:1064]
    entropy_src_hw2reg_entropy_data_reg_t entropy_data; // [1063:1032]
    entropy_src_hw2reg_repcnt_thresholds_reg_t repcnt_thresholds; // [1031:1000]
    entropy_src_hw2reg_repcnts_thresholds_reg_t repcnts_thresholds; // [999:968]
    entropy_src_hw2reg_adaptp_hi_thresholds_reg_t adaptp_hi_thresholds; // [967:936]
    entropy_src_hw2reg_adaptp_lo_thresholds_reg_t adaptp_lo_thresholds; // [935:904]
    entropy_src_hw2reg_bucket_thresholds_reg_t bucket_thresholds; // [903:872]
    entropy_src_hw2reg_markov_hi_thresholds_reg_t markov_hi_thresholds; // [871:840]
    entropy_src_hw2reg_markov_lo_thresholds_reg_t markov_lo_thresholds; // [839:808]
    entropy_src_hw2reg_extht_hi_thresholds_reg_t extht_hi_thresholds; // [807:776]
    entropy_src_hw2reg_extht_lo_thresholds_reg_t extht_lo_thresholds; // [775:744]
    entropy_src_hw2reg_repcnt_hi_watermarks_reg_t repcnt_hi_watermarks; // [743:712]
    entropy_src_hw2reg_repcnts_hi_watermarks_reg_t repcnts_hi_watermarks; // [711:680]
    entropy_src_hw2reg_adaptp_hi_watermarks_reg_t adaptp_hi_watermarks; // [679:648]
    entropy_src_hw2reg_adaptp_lo_watermarks_reg_t adaptp_lo_watermarks; // [647:616]
    entropy_src_hw2reg_extht_hi_watermarks_reg_t extht_hi_watermarks; // [615:584]
    entropy_src_hw2reg_extht_lo_watermarks_reg_t extht_lo_watermarks; // [583:552]
    entropy_src_hw2reg_bucket_hi_watermarks_reg_t bucket_hi_watermarks; // [551:520]
    entropy_src_hw2reg_markov_hi_watermarks_reg_t markov_hi_watermarks; // [519:488]
    entropy_src_hw2reg_markov_lo_watermarks_reg_t markov_lo_watermarks; // [487:456]
    entropy_src_hw2reg_repcnt_total_fails_reg_t repcnt_total_fails; // [455:424]
    entropy_src_hw2reg_repcnts_total_fails_reg_t repcnts_total_fails; // [423:392]
    entropy_src_hw2reg_adaptp_hi_total_fails_reg_t adaptp_hi_total_fails; // [391:360]
    entropy_src_hw2reg_adaptp_lo_total_fails_reg_t adaptp_lo_total_fails; // [359:328]
    entropy_src_hw2reg_bucket_total_fails_reg_t bucket_total_fails; // [327:296]
    entropy_src_hw2reg_markov_hi_total_fails_reg_t markov_hi_total_fails; // [295:264]
    entropy_src_hw2reg_markov_lo_total_fails_reg_t markov_lo_total_fails; // [263:232]
    entropy_src_hw2reg_extht_hi_total_fails_reg_t extht_hi_total_fails; // [231:200]
    entropy_src_hw2reg_extht_lo_total_fails_reg_t extht_lo_total_fails; // [199:168]
    entropy_src_hw2reg_alert_summary_fail_counts_reg_t alert_summary_fail_counts; // [167:152]
    entropy_src_hw2reg_alert_fail_counts_reg_t alert_fail_counts; // [151:124]
    entropy_src_hw2reg_extht_fail_counts_reg_t extht_fail_counts; // [123:116]
    entropy_src_hw2reg_fw_ov_wr_fifo_full_reg_t fw_ov_wr_fifo_full; // [115:115]
    entropy_src_hw2reg_fw_ov_rd_fifo_overflow_reg_t fw_ov_rd_fifo_overflow; // [114:113]
    entropy_src_hw2reg_fw_ov_rd_data_reg_t fw_ov_rd_data; // [112:81]
    entropy_src_hw2reg_observe_fifo_depth_reg_t observe_fifo_depth; // [80:74]
    entropy_src_hw2reg_debug_status_reg_t debug_status; // [73:62]
    entropy_src_hw2reg_recov_alert_sts_reg_t recov_alert_sts; // [61:32]
    entropy_src_hw2reg_err_code_reg_t err_code; // [31:10]
    entropy_src_hw2reg_main_sm_state_reg_t main_sm_state; // [9:0]
  } entropy_src_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] ENTROPY_SRC_INTR_STATE_OFFSET = 8'h 0;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_INTR_ENABLE_OFFSET = 8'h 4;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_INTR_TEST_OFFSET = 8'h 8;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ALERT_TEST_OFFSET = 8'h c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ME_REGWEN_OFFSET = 8'h 10;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_SW_REGUPD_OFFSET = 8'h 14;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REGWEN_OFFSET = 8'h 18;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REV_OFFSET = 8'h 1c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MODULE_ENABLE_OFFSET = 8'h 20;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_CONF_OFFSET = 8'h 24;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ENTROPY_CONTROL_OFFSET = 8'h 28;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ENTROPY_DATA_OFFSET = 8'h 2c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_HEALTH_TEST_WINDOWS_OFFSET = 8'h 30;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REPCNT_THRESHOLDS_OFFSET = 8'h 34;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REPCNTS_THRESHOLDS_OFFSET = 8'h 38;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ADAPTP_HI_THRESHOLDS_OFFSET = 8'h 3c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ADAPTP_LO_THRESHOLDS_OFFSET = 8'h 40;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_BUCKET_THRESHOLDS_OFFSET = 8'h 44;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MARKOV_HI_THRESHOLDS_OFFSET = 8'h 48;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MARKOV_LO_THRESHOLDS_OFFSET = 8'h 4c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_HI_THRESHOLDS_OFFSET = 8'h 50;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_LO_THRESHOLDS_OFFSET = 8'h 54;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REPCNT_HI_WATERMARKS_OFFSET = 8'h 58;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REPCNTS_HI_WATERMARKS_OFFSET = 8'h 5c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ADAPTP_HI_WATERMARKS_OFFSET = 8'h 60;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ADAPTP_LO_WATERMARKS_OFFSET = 8'h 64;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_HI_WATERMARKS_OFFSET = 8'h 68;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_LO_WATERMARKS_OFFSET = 8'h 6c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_BUCKET_HI_WATERMARKS_OFFSET = 8'h 70;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MARKOV_HI_WATERMARKS_OFFSET = 8'h 74;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MARKOV_LO_WATERMARKS_OFFSET = 8'h 78;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REPCNT_TOTAL_FAILS_OFFSET = 8'h 7c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_REPCNTS_TOTAL_FAILS_OFFSET = 8'h 80;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ADAPTP_HI_TOTAL_FAILS_OFFSET = 8'h 84;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ADAPTP_LO_TOTAL_FAILS_OFFSET = 8'h 88;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_BUCKET_TOTAL_FAILS_OFFSET = 8'h 8c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MARKOV_HI_TOTAL_FAILS_OFFSET = 8'h 90;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MARKOV_LO_TOTAL_FAILS_OFFSET = 8'h 94;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_HI_TOTAL_FAILS_OFFSET = 8'h 98;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_LO_TOTAL_FAILS_OFFSET = 8'h 9c;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ALERT_THRESHOLD_OFFSET = 8'h a0;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ALERT_SUMMARY_FAIL_COUNTS_OFFSET = 8'h a4;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ALERT_FAIL_COUNTS_OFFSET = 8'h a8;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_EXTHT_FAIL_COUNTS_OFFSET = 8'h ac;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_FW_OV_CONTROL_OFFSET = 8'h b0;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_FW_OV_SHA3_START_OFFSET = 8'h b4;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_FW_OV_WR_FIFO_FULL_OFFSET = 8'h b8;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_FW_OV_RD_FIFO_OVERFLOW_OFFSET = 8'h bc;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_FW_OV_RD_DATA_OFFSET = 8'h c0;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_FW_OV_WR_DATA_OFFSET = 8'h c4;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_OBSERVE_FIFO_THRESH_OFFSET = 8'h c8;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_OBSERVE_FIFO_DEPTH_OFFSET = 8'h cc;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_DEBUG_STATUS_OFFSET = 8'h d0;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_RECOV_ALERT_STS_OFFSET = 8'h d4;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ERR_CODE_OFFSET = 8'h d8;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_ERR_CODE_TEST_OFFSET = 8'h dc;
  parameter logic [BlockAw-1:0] ENTROPY_SRC_MAIN_SM_STATE_OFFSET = 8'h e0;

  // Reset values for hwext registers and their fields
  parameter logic [3:0] ENTROPY_SRC_INTR_TEST_RESVAL = 4'h 0;
  parameter logic [0:0] ENTROPY_SRC_INTR_TEST_ES_ENTROPY_VALID_RESVAL = 1'h 0;
  parameter logic [0:0] ENTROPY_SRC_INTR_TEST_ES_HEALTH_TEST_FAILED_RESVAL = 1'h 0;
  parameter logic [0:0] ENTROPY_SRC_INTR_TEST_ES_OBSERVE_FIFO_READY_RESVAL = 1'h 0;
  parameter logic [0:0] ENTROPY_SRC_INTR_TEST_ES_FATAL_ERR_RESVAL = 1'h 0;
  parameter logic [1:0] ENTROPY_SRC_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] ENTROPY_SRC_ALERT_TEST_RECOV_ALERT_RESVAL = 1'h 0;
  parameter logic [0:0] ENTROPY_SRC_ALERT_TEST_FATAL_ALERT_RESVAL = 1'h 0;
  parameter logic [31:0] ENTROPY_SRC_ENTROPY_DATA_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_REPCNT_THRESHOLDS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_REPCNT_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_REPCNT_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_REPCNTS_THRESHOLDS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_REPCNTS_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_REPCNTS_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_ADAPTP_HI_THRESHOLDS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_ADAPTP_HI_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_ADAPTP_HI_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_ADAPTP_LO_THRESHOLDS_RESVAL = 32'h 0;
  parameter logic [15:0] ENTROPY_SRC_ADAPTP_LO_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h 0;
  parameter logic [15:0] ENTROPY_SRC_ADAPTP_LO_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h 0;
  parameter logic [31:0] ENTROPY_SRC_BUCKET_THRESHOLDS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_BUCKET_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_BUCKET_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_MARKOV_HI_THRESHOLDS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_MARKOV_HI_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_MARKOV_HI_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_MARKOV_LO_THRESHOLDS_RESVAL = 32'h 0;
  parameter logic [15:0] ENTROPY_SRC_MARKOV_LO_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h 0;
  parameter logic [15:0] ENTROPY_SRC_MARKOV_LO_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h 0;
  parameter logic [31:0] ENTROPY_SRC_EXTHT_HI_THRESHOLDS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_EXTHT_HI_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_EXTHT_HI_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_EXTHT_LO_THRESHOLDS_RESVAL = 32'h 0;
  parameter logic [15:0] ENTROPY_SRC_EXTHT_LO_THRESHOLDS_FIPS_THRESH_RESVAL = 16'h 0;
  parameter logic [15:0] ENTROPY_SRC_EXTHT_LO_THRESHOLDS_BYPASS_THRESH_RESVAL = 16'h 0;
  parameter logic [31:0] ENTROPY_SRC_REPCNT_HI_WATERMARKS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_REPCNTS_HI_WATERMARKS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_ADAPTP_HI_WATERMARKS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_ADAPTP_LO_WATERMARKS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_ADAPTP_LO_WATERMARKS_FIPS_WATERMARK_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_ADAPTP_LO_WATERMARKS_BYPASS_WATERMARK_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_EXTHT_HI_WATERMARKS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_EXTHT_LO_WATERMARKS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_EXTHT_LO_WATERMARKS_FIPS_WATERMARK_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_EXTHT_LO_WATERMARKS_BYPASS_WATERMARK_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_BUCKET_HI_WATERMARKS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_MARKOV_HI_WATERMARKS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_MARKOV_LO_WATERMARKS_RESVAL = 32'h ffffffff;
  parameter logic [15:0] ENTROPY_SRC_MARKOV_LO_WATERMARKS_FIPS_WATERMARK_RESVAL = 16'h ffff;
  parameter logic [15:0] ENTROPY_SRC_MARKOV_LO_WATERMARKS_BYPASS_WATERMARK_RESVAL = 16'h ffff;
  parameter logic [31:0] ENTROPY_SRC_REPCNT_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_REPCNTS_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_ADAPTP_HI_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_ADAPTP_LO_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_BUCKET_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_MARKOV_HI_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_MARKOV_LO_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_EXTHT_HI_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_EXTHT_LO_TOTAL_FAILS_RESVAL = 32'h 0;
  parameter logic [15:0] ENTROPY_SRC_ALERT_SUMMARY_FAIL_COUNTS_RESVAL = 16'h 0;
  parameter logic [31:0] ENTROPY_SRC_ALERT_FAIL_COUNTS_RESVAL = 32'h 0;
  parameter logic [7:0] ENTROPY_SRC_EXTHT_FAIL_COUNTS_RESVAL = 8'h 0;
  parameter logic [0:0] ENTROPY_SRC_FW_OV_WR_FIFO_FULL_RESVAL = 1'h 0;
  parameter logic [31:0] ENTROPY_SRC_FW_OV_RD_DATA_RESVAL = 32'h 0;
  parameter logic [31:0] ENTROPY_SRC_FW_OV_WR_DATA_RESVAL = 32'h 0;
  parameter logic [6:0] ENTROPY_SRC_OBSERVE_FIFO_DEPTH_RESVAL = 7'h 0;
  parameter logic [17:0] ENTROPY_SRC_DEBUG_STATUS_RESVAL = 18'h 10000;
  parameter logic [0:0] ENTROPY_SRC_DEBUG_STATUS_MAIN_SM_IDLE_RESVAL = 1'h 1;

  // Register index
  typedef enum int {
    ENTROPY_SRC_INTR_STATE,
    ENTROPY_SRC_INTR_ENABLE,
    ENTROPY_SRC_INTR_TEST,
    ENTROPY_SRC_ALERT_TEST,
    ENTROPY_SRC_ME_REGWEN,
    ENTROPY_SRC_SW_REGUPD,
    ENTROPY_SRC_REGWEN,
    ENTROPY_SRC_REV,
    ENTROPY_SRC_MODULE_ENABLE,
    ENTROPY_SRC_CONF,
    ENTROPY_SRC_ENTROPY_CONTROL,
    ENTROPY_SRC_ENTROPY_DATA,
    ENTROPY_SRC_HEALTH_TEST_WINDOWS,
    ENTROPY_SRC_REPCNT_THRESHOLDS,
    ENTROPY_SRC_REPCNTS_THRESHOLDS,
    ENTROPY_SRC_ADAPTP_HI_THRESHOLDS,
    ENTROPY_SRC_ADAPTP_LO_THRESHOLDS,
    ENTROPY_SRC_BUCKET_THRESHOLDS,
    ENTROPY_SRC_MARKOV_HI_THRESHOLDS,
    ENTROPY_SRC_MARKOV_LO_THRESHOLDS,
    ENTROPY_SRC_EXTHT_HI_THRESHOLDS,
    ENTROPY_SRC_EXTHT_LO_THRESHOLDS,
    ENTROPY_SRC_REPCNT_HI_WATERMARKS,
    ENTROPY_SRC_REPCNTS_HI_WATERMARKS,
    ENTROPY_SRC_ADAPTP_HI_WATERMARKS,
    ENTROPY_SRC_ADAPTP_LO_WATERMARKS,
    ENTROPY_SRC_EXTHT_HI_WATERMARKS,
    ENTROPY_SRC_EXTHT_LO_WATERMARKS,
    ENTROPY_SRC_BUCKET_HI_WATERMARKS,
    ENTROPY_SRC_MARKOV_HI_WATERMARKS,
    ENTROPY_SRC_MARKOV_LO_WATERMARKS,
    ENTROPY_SRC_REPCNT_TOTAL_FAILS,
    ENTROPY_SRC_REPCNTS_TOTAL_FAILS,
    ENTROPY_SRC_ADAPTP_HI_TOTAL_FAILS,
    ENTROPY_SRC_ADAPTP_LO_TOTAL_FAILS,
    ENTROPY_SRC_BUCKET_TOTAL_FAILS,
    ENTROPY_SRC_MARKOV_HI_TOTAL_FAILS,
    ENTROPY_SRC_MARKOV_LO_TOTAL_FAILS,
    ENTROPY_SRC_EXTHT_HI_TOTAL_FAILS,
    ENTROPY_SRC_EXTHT_LO_TOTAL_FAILS,
    ENTROPY_SRC_ALERT_THRESHOLD,
    ENTROPY_SRC_ALERT_SUMMARY_FAIL_COUNTS,
    ENTROPY_SRC_ALERT_FAIL_COUNTS,
    ENTROPY_SRC_EXTHT_FAIL_COUNTS,
    ENTROPY_SRC_FW_OV_CONTROL,
    ENTROPY_SRC_FW_OV_SHA3_START,
    ENTROPY_SRC_FW_OV_WR_FIFO_FULL,
    ENTROPY_SRC_FW_OV_RD_FIFO_OVERFLOW,
    ENTROPY_SRC_FW_OV_RD_DATA,
    ENTROPY_SRC_FW_OV_WR_DATA,
    ENTROPY_SRC_OBSERVE_FIFO_THRESH,
    ENTROPY_SRC_OBSERVE_FIFO_DEPTH,
    ENTROPY_SRC_DEBUG_STATUS,
    ENTROPY_SRC_RECOV_ALERT_STS,
    ENTROPY_SRC_ERR_CODE,
    ENTROPY_SRC_ERR_CODE_TEST,
    ENTROPY_SRC_MAIN_SM_STATE
  } entropy_src_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] ENTROPY_SRC_PERMIT [57] = '{
    4'b 0001, // index[ 0] ENTROPY_SRC_INTR_STATE
    4'b 0001, // index[ 1] ENTROPY_SRC_INTR_ENABLE
    4'b 0001, // index[ 2] ENTROPY_SRC_INTR_TEST
    4'b 0001, // index[ 3] ENTROPY_SRC_ALERT_TEST
    4'b 0001, // index[ 4] ENTROPY_SRC_ME_REGWEN
    4'b 0001, // index[ 5] ENTROPY_SRC_SW_REGUPD
    4'b 0001, // index[ 6] ENTROPY_SRC_REGWEN
    4'b 0111, // index[ 7] ENTROPY_SRC_REV
    4'b 0001, // index[ 8] ENTROPY_SRC_MODULE_ENABLE
    4'b 1111, // index[ 9] ENTROPY_SRC_CONF
    4'b 0001, // index[10] ENTROPY_SRC_ENTROPY_CONTROL
    4'b 1111, // index[11] ENTROPY_SRC_ENTROPY_DATA
    4'b 1111, // index[12] ENTROPY_SRC_HEALTH_TEST_WINDOWS
    4'b 1111, // index[13] ENTROPY_SRC_REPCNT_THRESHOLDS
    4'b 1111, // index[14] ENTROPY_SRC_REPCNTS_THRESHOLDS
    4'b 1111, // index[15] ENTROPY_SRC_ADAPTP_HI_THRESHOLDS
    4'b 1111, // index[16] ENTROPY_SRC_ADAPTP_LO_THRESHOLDS
    4'b 1111, // index[17] ENTROPY_SRC_BUCKET_THRESHOLDS
    4'b 1111, // index[18] ENTROPY_SRC_MARKOV_HI_THRESHOLDS
    4'b 1111, // index[19] ENTROPY_SRC_MARKOV_LO_THRESHOLDS
    4'b 1111, // index[20] ENTROPY_SRC_EXTHT_HI_THRESHOLDS
    4'b 1111, // index[21] ENTROPY_SRC_EXTHT_LO_THRESHOLDS
    4'b 1111, // index[22] ENTROPY_SRC_REPCNT_HI_WATERMARKS
    4'b 1111, // index[23] ENTROPY_SRC_REPCNTS_HI_WATERMARKS
    4'b 1111, // index[24] ENTROPY_SRC_ADAPTP_HI_WATERMARKS
    4'b 1111, // index[25] ENTROPY_SRC_ADAPTP_LO_WATERMARKS
    4'b 1111, // index[26] ENTROPY_SRC_EXTHT_HI_WATERMARKS
    4'b 1111, // index[27] ENTROPY_SRC_EXTHT_LO_WATERMARKS
    4'b 1111, // index[28] ENTROPY_SRC_BUCKET_HI_WATERMARKS
    4'b 1111, // index[29] ENTROPY_SRC_MARKOV_HI_WATERMARKS
    4'b 1111, // index[30] ENTROPY_SRC_MARKOV_LO_WATERMARKS
    4'b 1111, // index[31] ENTROPY_SRC_REPCNT_TOTAL_FAILS
    4'b 1111, // index[32] ENTROPY_SRC_REPCNTS_TOTAL_FAILS
    4'b 1111, // index[33] ENTROPY_SRC_ADAPTP_HI_TOTAL_FAILS
    4'b 1111, // index[34] ENTROPY_SRC_ADAPTP_LO_TOTAL_FAILS
    4'b 1111, // index[35] ENTROPY_SRC_BUCKET_TOTAL_FAILS
    4'b 1111, // index[36] ENTROPY_SRC_MARKOV_HI_TOTAL_FAILS
    4'b 1111, // index[37] ENTROPY_SRC_MARKOV_LO_TOTAL_FAILS
    4'b 1111, // index[38] ENTROPY_SRC_EXTHT_HI_TOTAL_FAILS
    4'b 1111, // index[39] ENTROPY_SRC_EXTHT_LO_TOTAL_FAILS
    4'b 1111, // index[40] ENTROPY_SRC_ALERT_THRESHOLD
    4'b 0011, // index[41] ENTROPY_SRC_ALERT_SUMMARY_FAIL_COUNTS
    4'b 1111, // index[42] ENTROPY_SRC_ALERT_FAIL_COUNTS
    4'b 0001, // index[43] ENTROPY_SRC_EXTHT_FAIL_COUNTS
    4'b 0001, // index[44] ENTROPY_SRC_FW_OV_CONTROL
    4'b 0001, // index[45] ENTROPY_SRC_FW_OV_SHA3_START
    4'b 0001, // index[46] ENTROPY_SRC_FW_OV_WR_FIFO_FULL
    4'b 0001, // index[47] ENTROPY_SRC_FW_OV_RD_FIFO_OVERFLOW
    4'b 1111, // index[48] ENTROPY_SRC_FW_OV_RD_DATA
    4'b 1111, // index[49] ENTROPY_SRC_FW_OV_WR_DATA
    4'b 0001, // index[50] ENTROPY_SRC_OBSERVE_FIFO_THRESH
    4'b 0001, // index[51] ENTROPY_SRC_OBSERVE_FIFO_DEPTH
    4'b 0111, // index[52] ENTROPY_SRC_DEBUG_STATUS
    4'b 0111, // index[53] ENTROPY_SRC_RECOV_ALERT_STS
    4'b 1111, // index[54] ENTROPY_SRC_ERR_CODE
    4'b 0001, // index[55] ENTROPY_SRC_ERR_CODE_TEST
    4'b 0011  // index[56] ENTROPY_SRC_MAIN_SM_STATE
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module entropy_src_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output entropy_src_reg_pkg::entropy_src_reg2hw_t reg2hw, // Write
  input  entropy_src_reg_pkg::entropy_src_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import entropy_src_reg_pkg::* ;

  localparam int AW = 8;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [56:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(57)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_es_entropy_valid_qs;
  logic intr_state_es_entropy_valid_wd;
  logic intr_state_es_health_test_failed_qs;
  logic intr_state_es_health_test_failed_wd;
  logic intr_state_es_observe_fifo_ready_qs;
  logic intr_state_es_observe_fifo_ready_wd;
  logic intr_state_es_fatal_err_qs;
  logic intr_state_es_fatal_err_wd;
  logic intr_enable_we;
  logic intr_enable_es_entropy_valid_qs;
  logic intr_enable_es_entropy_valid_wd;
  logic intr_enable_es_health_test_failed_qs;
  logic intr_enable_es_health_test_failed_wd;
  logic intr_enable_es_observe_fifo_ready_qs;
  logic intr_enable_es_observe_fifo_ready_wd;
  logic intr_enable_es_fatal_err_qs;
  logic intr_enable_es_fatal_err_wd;
  logic intr_test_we;
  logic intr_test_es_entropy_valid_wd;
  logic intr_test_es_health_test_failed_wd;
  logic intr_test_es_observe_fifo_ready_wd;
  logic intr_test_es_fatal_err_wd;
  logic alert_test_we;
  logic alert_test_recov_alert_wd;
  logic alert_test_fatal_alert_wd;
  logic me_regwen_we;
  logic me_regwen_qs;
  logic me_regwen_wd;
  logic sw_regupd_we;
  logic sw_regupd_qs;
  logic sw_regupd_wd;
  logic regwen_qs;
  logic [7:0] rev_abi_revision_qs;
  logic [7:0] rev_hw_revision_qs;
  logic [7:0] rev_chip_type_qs;
  logic module_enable_we;
  logic [3:0] module_enable_qs;
  logic [3:0] module_enable_wd;
  logic conf_we;
  logic [3:0] conf_fips_enable_qs;
  logic [3:0] conf_fips_enable_wd;
  logic [3:0] conf_entropy_data_reg_enable_qs;
  logic [3:0] conf_entropy_data_reg_enable_wd;
  logic [3:0] conf_threshold_scope_qs;
  logic [3:0] conf_threshold_scope_wd;
  logic [3:0] conf_rng_bit_enable_qs;
  logic [3:0] conf_rng_bit_enable_wd;
  logic [1:0] conf_rng_bit_sel_qs;
  logic [1:0] conf_rng_bit_sel_wd;
  logic entropy_control_we;
  logic [3:0] entropy_control_es_route_qs;
  logic [3:0] entropy_control_es_route_wd;
  logic [3:0] entropy_control_es_type_qs;
  logic [3:0] entropy_control_es_type_wd;
  logic entropy_data_re;
  logic [31:0] entropy_data_qs;
  logic health_test_windows_we;
  logic [15:0] health_test_windows_fips_window_qs;
  logic [15:0] health_test_windows_fips_window_wd;
  logic [15:0] health_test_windows_bypass_window_qs;
  logic [15:0] health_test_windows_bypass_window_wd;
  logic repcnt_thresholds_re;
  logic repcnt_thresholds_we;
  logic [15:0] repcnt_thresholds_fips_thresh_qs;
  logic [15:0] repcnt_thresholds_fips_thresh_wd;
  logic [15:0] repcnt_thresholds_bypass_thresh_qs;
  logic [15:0] repcnt_thresholds_bypass_thresh_wd;
  logic repcnts_thresholds_re;
  logic repcnts_thresholds_we;
  logic [15:0] repcnts_thresholds_fips_thresh_qs;
  logic [15:0] repcnts_thresholds_fips_thresh_wd;
  logic [15:0] repcnts_thresholds_bypass_thresh_qs;
  logic [15:0] repcnts_thresholds_bypass_thresh_wd;
  logic adaptp_hi_thresholds_re;
  logic adaptp_hi_thresholds_we;
  logic [15:0] adaptp_hi_thresholds_fips_thresh_qs;
  logic [15:0] adaptp_hi_thresholds_fips_thresh_wd;
  logic [15:0] adaptp_hi_thresholds_bypass_thresh_qs;
  logic [15:0] adaptp_hi_thresholds_bypass_thresh_wd;
  logic adaptp_lo_thresholds_re;
  logic adaptp_lo_thresholds_we;
  logic [15:0] adaptp_lo_thresholds_fips_thresh_qs;
  logic [15:0] adaptp_lo_thresholds_fips_thresh_wd;
  logic [15:0] adaptp_lo_thresholds_bypass_thresh_qs;
  logic [15:0] adaptp_lo_thresholds_bypass_thresh_wd;
  logic bucket_thresholds_re;
  logic bucket_thresholds_we;
  logic [15:0] bucket_thresholds_fips_thresh_qs;
  logic [15:0] bucket_thresholds_fips_thresh_wd;
  logic [15:0] bucket_thresholds_bypass_thresh_qs;
  logic [15:0] bucket_thresholds_bypass_thresh_wd;
  logic markov_hi_thresholds_re;
  logic markov_hi_thresholds_we;
  logic [15:0] markov_hi_thresholds_fips_thresh_qs;
  logic [15:0] markov_hi_thresholds_fips_thresh_wd;
  logic [15:0] markov_hi_thresholds_bypass_thresh_qs;
  logic [15:0] markov_hi_thresholds_bypass_thresh_wd;
  logic markov_lo_thresholds_re;
  logic markov_lo_thresholds_we;
  logic [15:0] markov_lo_thresholds_fips_thresh_qs;
  logic [15:0] markov_lo_thresholds_fips_thresh_wd;
  logic [15:0] markov_lo_thresholds_bypass_thresh_qs;
  logic [15:0] markov_lo_thresholds_bypass_thresh_wd;
  logic extht_hi_thresholds_re;
  logic extht_hi_thresholds_we;
  logic [15:0] extht_hi_thresholds_fips_thresh_qs;
  logic [15:0] extht_hi_thresholds_fips_thresh_wd;
  logic [15:0] extht_hi_thresholds_bypass_thresh_qs;
  logic [15:0] extht_hi_thresholds_bypass_thresh_wd;
  logic extht_lo_thresholds_re;
  logic extht_lo_thresholds_we;
  logic [15:0] extht_lo_thresholds_fips_thresh_qs;
  logic [15:0] extht_lo_thresholds_fips_thresh_wd;
  logic [15:0] extht_lo_thresholds_bypass_thresh_qs;
  logic [15:0] extht_lo_thresholds_bypass_thresh_wd;
  logic repcnt_hi_watermarks_re;
  logic [15:0] repcnt_hi_watermarks_fips_watermark_qs;
  logic [15:0] repcnt_hi_watermarks_bypass_watermark_qs;
  logic repcnts_hi_watermarks_re;
  logic [15:0] repcnts_hi_watermarks_fips_watermark_qs;
  logic [15:0] repcnts_hi_watermarks_bypass_watermark_qs;
  logic adaptp_hi_watermarks_re;
  logic [15:0] adaptp_hi_watermarks_fips_watermark_qs;
  logic [15:0] adaptp_hi_watermarks_bypass_watermark_qs;
  logic adaptp_lo_watermarks_re;
  logic [15:0] adaptp_lo_watermarks_fips_watermark_qs;
  logic [15:0] adaptp_lo_watermarks_bypass_watermark_qs;
  logic extht_hi_watermarks_re;
  logic [15:0] extht_hi_watermarks_fips_watermark_qs;
  logic [15:0] extht_hi_watermarks_bypass_watermark_qs;
  logic extht_lo_watermarks_re;
  logic [15:0] extht_lo_watermarks_fips_watermark_qs;
  logic [15:0] extht_lo_watermarks_bypass_watermark_qs;
  logic bucket_hi_watermarks_re;
  logic [15:0] bucket_hi_watermarks_fips_watermark_qs;
  logic [15:0] bucket_hi_watermarks_bypass_watermark_qs;
  logic markov_hi_watermarks_re;
  logic [15:0] markov_hi_watermarks_fips_watermark_qs;
  logic [15:0] markov_hi_watermarks_bypass_watermark_qs;
  logic markov_lo_watermarks_re;
  logic [15:0] markov_lo_watermarks_fips_watermark_qs;
  logic [15:0] markov_lo_watermarks_bypass_watermark_qs;
  logic repcnt_total_fails_re;
  logic [31:0] repcnt_total_fails_qs;
  logic repcnts_total_fails_re;
  logic [31:0] repcnts_total_fails_qs;
  logic adaptp_hi_total_fails_re;
  logic [31:0] adaptp_hi_total_fails_qs;
  logic adaptp_lo_total_fails_re;
  logic [31:0] adaptp_lo_total_fails_qs;
  logic bucket_total_fails_re;
  logic [31:0] bucket_total_fails_qs;
  logic markov_hi_total_fails_re;
  logic [31:0] markov_hi_total_fails_qs;
  logic markov_lo_total_fails_re;
  logic [31:0] markov_lo_total_fails_qs;
  logic extht_hi_total_fails_re;
  logic [31:0] extht_hi_total_fails_qs;
  logic extht_lo_total_fails_re;
  logic [31:0] extht_lo_total_fails_qs;
  logic alert_threshold_we;
  logic [15:0] alert_threshold_alert_threshold_qs;
  logic [15:0] alert_threshold_alert_threshold_wd;
  logic [15:0] alert_threshold_alert_threshold_inv_qs;
  logic [15:0] alert_threshold_alert_threshold_inv_wd;
  logic alert_summary_fail_counts_re;
  logic [15:0] alert_summary_fail_counts_qs;
  logic alert_fail_counts_re;
  logic [3:0] alert_fail_counts_repcnt_fail_count_qs;
  logic [3:0] alert_fail_counts_adaptp_hi_fail_count_qs;
  logic [3:0] alert_fail_counts_adaptp_lo_fail_count_qs;
  logic [3:0] alert_fail_counts_bucket_fail_count_qs;
  logic [3:0] alert_fail_counts_markov_hi_fail_count_qs;
  logic [3:0] alert_fail_counts_markov_lo_fail_count_qs;
  logic [3:0] alert_fail_counts_repcnts_fail_count_qs;
  logic extht_fail_counts_re;
  logic [3:0] extht_fail_counts_extht_hi_fail_count_qs;
  logic [3:0] extht_fail_counts_extht_lo_fail_count_qs;
  logic fw_ov_control_we;
  logic [3:0] fw_ov_control_fw_ov_mode_qs;
  logic [3:0] fw_ov_control_fw_ov_mode_wd;
  logic [3:0] fw_ov_control_fw_ov_entropy_insert_qs;
  logic [3:0] fw_ov_control_fw_ov_entropy_insert_wd;
  logic fw_ov_sha3_start_we;
  logic [3:0] fw_ov_sha3_start_qs;
  logic [3:0] fw_ov_sha3_start_wd;
  logic fw_ov_wr_fifo_full_re;
  logic fw_ov_wr_fifo_full_qs;
  logic fw_ov_rd_fifo_overflow_we;
  logic fw_ov_rd_fifo_overflow_qs;
  logic fw_ov_rd_fifo_overflow_wd;
  logic fw_ov_rd_data_re;
  logic [31:0] fw_ov_rd_data_qs;
  logic fw_ov_wr_data_we;
  logic [31:0] fw_ov_wr_data_wd;
  logic observe_fifo_thresh_we;
  logic [6:0] observe_fifo_thresh_qs;
  logic [6:0] observe_fifo_thresh_wd;
  logic observe_fifo_depth_re;
  logic [6:0] observe_fifo_depth_qs;
  logic debug_status_re;
  logic [2:0] debug_status_entropy_fifo_depth_qs;
  logic [2:0] debug_status_sha3_fsm_qs;
  logic debug_status_sha3_block_pr_qs;
  logic debug_status_sha3_squeezing_qs;
  logic debug_status_sha3_absorbed_qs;
  logic debug_status_sha3_err_qs;
  logic debug_status_main_sm_idle_qs;
  logic debug_status_main_sm_boot_done_qs;
  logic recov_alert_sts_we;
  logic recov_alert_sts_fips_enable_field_alert_qs;
  logic recov_alert_sts_fips_enable_field_alert_wd;
  logic recov_alert_sts_entropy_data_reg_en_field_alert_qs;
  logic recov_alert_sts_entropy_data_reg_en_field_alert_wd;
  logic recov_alert_sts_module_enable_field_alert_qs;
  logic recov_alert_sts_module_enable_field_alert_wd;
  logic recov_alert_sts_threshold_scope_field_alert_qs;
  logic recov_alert_sts_threshold_scope_field_alert_wd;
  logic recov_alert_sts_rng_bit_enable_field_alert_qs;
  logic recov_alert_sts_rng_bit_enable_field_alert_wd;
  logic recov_alert_sts_fw_ov_sha3_start_field_alert_qs;
  logic recov_alert_sts_fw_ov_sha3_start_field_alert_wd;
  logic recov_alert_sts_fw_ov_mode_field_alert_qs;
  logic recov_alert_sts_fw_ov_mode_field_alert_wd;
  logic recov_alert_sts_fw_ov_entropy_insert_field_alert_qs;
  logic recov_alert_sts_fw_ov_entropy_insert_field_alert_wd;
  logic recov_alert_sts_es_route_field_alert_qs;
  logic recov_alert_sts_es_route_field_alert_wd;
  logic recov_alert_sts_es_type_field_alert_qs;
  logic recov_alert_sts_es_type_field_alert_wd;
  logic recov_alert_sts_es_main_sm_alert_qs;
  logic recov_alert_sts_es_main_sm_alert_wd;
  logic recov_alert_sts_es_bus_cmp_alert_qs;
  logic recov_alert_sts_es_bus_cmp_alert_wd;
  logic recov_alert_sts_es_thresh_cfg_alert_qs;
  logic recov_alert_sts_es_thresh_cfg_alert_wd;
  logic recov_alert_sts_es_fw_ov_wr_alert_qs;
  logic recov_alert_sts_es_fw_ov_wr_alert_wd;
  logic recov_alert_sts_es_fw_ov_disable_alert_qs;
  logic recov_alert_sts_es_fw_ov_disable_alert_wd;
  logic err_code_sfifo_esrng_err_qs;
  logic err_code_sfifo_observe_err_qs;
  logic err_code_sfifo_esfinal_err_qs;
  logic err_code_es_ack_sm_err_qs;
  logic err_code_es_main_sm_err_qs;
  logic err_code_es_cntr_err_qs;
  logic err_code_sha3_state_err_qs;
  logic err_code_sha3_rst_storage_err_qs;
  logic err_code_fifo_write_err_qs;
  logic err_code_fifo_read_err_qs;
  logic err_code_fifo_state_err_qs;
  logic err_code_test_we;
  logic [4:0] err_code_test_qs;
  logic [4:0] err_code_test_wd;
  logic [8:0] main_sm_state_qs;

  // Register instances
  // R[intr_state]: V(False)
  //   F[es_entropy_valid]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_es_entropy_valid (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_es_entropy_valid_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.es_entropy_valid.de),
    .d      (hw2reg.intr_state.es_entropy_valid.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.es_entropy_valid.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_es_entropy_valid_qs)
  );

  //   F[es_health_test_failed]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_es_health_test_failed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_es_health_test_failed_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.es_health_test_failed.de),
    .d      (hw2reg.intr_state.es_health_test_failed.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.es_health_test_failed.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_es_health_test_failed_qs)
  );

  //   F[es_observe_fifo_ready]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_es_observe_fifo_ready (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_es_observe_fifo_ready_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.es_observe_fifo_ready.de),
    .d      (hw2reg.intr_state.es_observe_fifo_ready.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.es_observe_fifo_ready.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_es_observe_fifo_ready_qs)
  );

  //   F[es_fatal_err]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_es_fatal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_es_fatal_err_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.es_fatal_err.de),
    .d      (hw2reg.intr_state.es_fatal_err.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.es_fatal_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_es_fatal_err_qs)
  );


  // R[intr_enable]: V(False)
  //   F[es_entropy_valid]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_es_entropy_valid (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_es_entropy_valid_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.es_entropy_valid.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_es_entropy_valid_qs)
  );

  //   F[es_health_test_failed]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_es_health_test_failed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_es_health_test_failed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.es_health_test_failed.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_es_health_test_failed_qs)
  );

  //   F[es_observe_fifo_ready]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_es_observe_fifo_ready (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_es_observe_fifo_ready_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.es_observe_fifo_ready.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_es_observe_fifo_ready_qs)
  );

  //   F[es_fatal_err]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_es_fatal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_es_fatal_err_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.es_fatal_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_es_fatal_err_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [3:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  //   F[es_entropy_valid]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_es_entropy_valid (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_es_entropy_valid_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.es_entropy_valid.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.es_entropy_valid.qe = intr_test_qe;

  //   F[es_health_test_failed]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_es_health_test_failed (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_es_health_test_failed_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[1]),
    .q      (reg2hw.intr_test.es_health_test_failed.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.es_health_test_failed.qe = intr_test_qe;

  //   F[es_observe_fifo_ready]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_es_observe_fifo_ready (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_es_observe_fifo_ready_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[2]),
    .q      (reg2hw.intr_test.es_observe_fifo_ready.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.es_observe_fifo_ready.qe = intr_test_qe;

  //   F[es_fatal_err]: 3:3
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_es_fatal_err (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_es_fatal_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[3]),
    .q      (reg2hw.intr_test.es_fatal_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.es_fatal_err.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[recov_alert]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov_alert (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_alert_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.recov_alert.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov_alert.qe = alert_test_qe;

  //   F[fatal_alert]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal_alert (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_alert_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.fatal_alert.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal_alert.qe = alert_test_qe;


  // R[me_regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_me_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (me_regwen_we),
    .wd     (me_regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (me_regwen_qs)
  );


  // R[sw_regupd]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_sw_regupd (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_regupd_we),
    .wd     (sw_regupd_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sw_regupd.q),
    .ds     (),

    // to register interface (read)
    .qs     (sw_regupd_qs)
  );


  // R[regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h1)
  ) u_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.regwen.de),
    .d      (hw2reg.regwen.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (regwen_qs)
  );


  // R[rev]: V(False)
  //   F[abi_revision]: 7:0
  // constant-only read
  assign rev_abi_revision_qs = 8'h3;

  //   F[hw_revision]: 15:8
  // constant-only read
  assign rev_hw_revision_qs = 8'h3;

  //   F[chip_type]: 23:16
  // constant-only read
  assign rev_chip_type_qs = 8'h1;


  // R[module_enable]: V(False)
  // Create REGWEN-gated WE signal
  logic module_enable_gated_we;
  assign module_enable_gated_we = module_enable_we & me_regwen_qs;
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_module_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (module_enable_gated_we),
    .wd     (module_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.module_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (module_enable_qs)
  );


  // R[conf]: V(False)
  // Create REGWEN-gated WE signal
  logic conf_gated_we;
  assign conf_gated_we = conf_we & regwen_qs;
  //   F[fips_enable]: 3:0
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_conf_fips_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (conf_gated_we),
    .wd     (conf_fips_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.conf.fips_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (conf_fips_enable_qs)
  );

  //   F[entropy_data_reg_enable]: 7:4
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_conf_entropy_data_reg_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (conf_gated_we),
    .wd     (conf_entropy_data_reg_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.conf.entropy_data_reg_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (conf_entropy_data_reg_enable_qs)
  );

  //   F[threshold_scope]: 15:12
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_conf_threshold_scope (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (conf_gated_we),
    .wd     (conf_threshold_scope_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.conf.threshold_scope.q),
    .ds     (),

    // to register interface (read)
    .qs     (conf_threshold_scope_qs)
  );

  //   F[rng_bit_enable]: 23:20
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_conf_rng_bit_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (conf_gated_we),
    .wd     (conf_rng_bit_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.conf.rng_bit_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (conf_rng_bit_enable_qs)
  );

  //   F[rng_bit_sel]: 25:24
  prim_subreg #(
    .DW      (2),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (2'h0)
  ) u_conf_rng_bit_sel (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (conf_gated_we),
    .wd     (conf_rng_bit_sel_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.conf.rng_bit_sel.q),
    .ds     (),

    // to register interface (read)
    .qs     (conf_rng_bit_sel_qs)
  );


  // R[entropy_control]: V(False)
  // Create REGWEN-gated WE signal
  logic entropy_control_gated_we;
  assign entropy_control_gated_we = entropy_control_we & regwen_qs;
  //   F[es_route]: 3:0
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_entropy_control_es_route (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (entropy_control_gated_we),
    .wd     (entropy_control_es_route_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.entropy_control.es_route.q),
    .ds     (),

    // to register interface (read)
    .qs     (entropy_control_es_route_qs)
  );

  //   F[es_type]: 7:4
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_entropy_control_es_type (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (entropy_control_gated_we),
    .wd     (entropy_control_es_type_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.entropy_control.es_type.q),
    .ds     (),

    // to register interface (read)
    .qs     (entropy_control_es_type_qs)
  );


  // R[entropy_data]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_entropy_data (
    .re     (entropy_data_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.entropy_data.d),
    .qre    (reg2hw.entropy_data.re),
    .qe     (),
    .q      (reg2hw.entropy_data.q),
    .ds     (),
    .qs     (entropy_data_qs)
  );


  // R[health_test_windows]: V(False)
  // Create REGWEN-gated WE signal
  logic health_test_windows_gated_we;
  assign health_test_windows_gated_we = health_test_windows_we & regwen_qs;
  //   F[fips_window]: 15:0
  prim_subreg #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h200)
  ) u_health_test_windows_fips_window (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (health_test_windows_gated_we),
    .wd     (health_test_windows_fips_window_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.health_test_windows.fips_window.q),
    .ds     (),

    // to register interface (read)
    .qs     (health_test_windows_fips_window_qs)
  );

  //   F[bypass_window]: 31:16
  prim_subreg #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h60)
  ) u_health_test_windows_bypass_window (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (health_test_windows_gated_we),
    .wd     (health_test_windows_bypass_window_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.health_test_windows.bypass_window.q),
    .ds     (),

    // to register interface (read)
    .qs     (health_test_windows_bypass_window_qs)
  );


  // R[repcnt_thresholds]: V(True)
  logic repcnt_thresholds_qe;
  logic [1:0] repcnt_thresholds_flds_we;
  assign repcnt_thresholds_qe = &repcnt_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic repcnt_thresholds_gated_we;
  assign repcnt_thresholds_gated_we = repcnt_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnt_thresholds_fips_thresh (
    .re     (repcnt_thresholds_re),
    .we     (repcnt_thresholds_gated_we),
    .wd     (repcnt_thresholds_fips_thresh_wd),
    .d      (hw2reg.repcnt_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (repcnt_thresholds_flds_we[0]),
    .q      (reg2hw.repcnt_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (repcnt_thresholds_fips_thresh_qs)
  );
  assign reg2hw.repcnt_thresholds.fips_thresh.qe = repcnt_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnt_thresholds_bypass_thresh (
    .re     (repcnt_thresholds_re),
    .we     (repcnt_thresholds_gated_we),
    .wd     (repcnt_thresholds_bypass_thresh_wd),
    .d      (hw2reg.repcnt_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (repcnt_thresholds_flds_we[1]),
    .q      (reg2hw.repcnt_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (repcnt_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.repcnt_thresholds.bypass_thresh.qe = repcnt_thresholds_qe;


  // R[repcnts_thresholds]: V(True)
  logic repcnts_thresholds_qe;
  logic [1:0] repcnts_thresholds_flds_we;
  assign repcnts_thresholds_qe = &repcnts_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic repcnts_thresholds_gated_we;
  assign repcnts_thresholds_gated_we = repcnts_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnts_thresholds_fips_thresh (
    .re     (repcnts_thresholds_re),
    .we     (repcnts_thresholds_gated_we),
    .wd     (repcnts_thresholds_fips_thresh_wd),
    .d      (hw2reg.repcnts_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (repcnts_thresholds_flds_we[0]),
    .q      (reg2hw.repcnts_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (repcnts_thresholds_fips_thresh_qs)
  );
  assign reg2hw.repcnts_thresholds.fips_thresh.qe = repcnts_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnts_thresholds_bypass_thresh (
    .re     (repcnts_thresholds_re),
    .we     (repcnts_thresholds_gated_we),
    .wd     (repcnts_thresholds_bypass_thresh_wd),
    .d      (hw2reg.repcnts_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (repcnts_thresholds_flds_we[1]),
    .q      (reg2hw.repcnts_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (repcnts_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.repcnts_thresholds.bypass_thresh.qe = repcnts_thresholds_qe;


  // R[adaptp_hi_thresholds]: V(True)
  logic adaptp_hi_thresholds_qe;
  logic [1:0] adaptp_hi_thresholds_flds_we;
  assign adaptp_hi_thresholds_qe = &adaptp_hi_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic adaptp_hi_thresholds_gated_we;
  assign adaptp_hi_thresholds_gated_we = adaptp_hi_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_hi_thresholds_fips_thresh (
    .re     (adaptp_hi_thresholds_re),
    .we     (adaptp_hi_thresholds_gated_we),
    .wd     (adaptp_hi_thresholds_fips_thresh_wd),
    .d      (hw2reg.adaptp_hi_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (adaptp_hi_thresholds_flds_we[0]),
    .q      (reg2hw.adaptp_hi_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (adaptp_hi_thresholds_fips_thresh_qs)
  );
  assign reg2hw.adaptp_hi_thresholds.fips_thresh.qe = adaptp_hi_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_hi_thresholds_bypass_thresh (
    .re     (adaptp_hi_thresholds_re),
    .we     (adaptp_hi_thresholds_gated_we),
    .wd     (adaptp_hi_thresholds_bypass_thresh_wd),
    .d      (hw2reg.adaptp_hi_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (adaptp_hi_thresholds_flds_we[1]),
    .q      (reg2hw.adaptp_hi_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (adaptp_hi_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.adaptp_hi_thresholds.bypass_thresh.qe = adaptp_hi_thresholds_qe;


  // R[adaptp_lo_thresholds]: V(True)
  logic adaptp_lo_thresholds_qe;
  logic [1:0] adaptp_lo_thresholds_flds_we;
  assign adaptp_lo_thresholds_qe = &adaptp_lo_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic adaptp_lo_thresholds_gated_we;
  assign adaptp_lo_thresholds_gated_we = adaptp_lo_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_lo_thresholds_fips_thresh (
    .re     (adaptp_lo_thresholds_re),
    .we     (adaptp_lo_thresholds_gated_we),
    .wd     (adaptp_lo_thresholds_fips_thresh_wd),
    .d      (hw2reg.adaptp_lo_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (adaptp_lo_thresholds_flds_we[0]),
    .q      (reg2hw.adaptp_lo_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (adaptp_lo_thresholds_fips_thresh_qs)
  );
  assign reg2hw.adaptp_lo_thresholds.fips_thresh.qe = adaptp_lo_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_lo_thresholds_bypass_thresh (
    .re     (adaptp_lo_thresholds_re),
    .we     (adaptp_lo_thresholds_gated_we),
    .wd     (adaptp_lo_thresholds_bypass_thresh_wd),
    .d      (hw2reg.adaptp_lo_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (adaptp_lo_thresholds_flds_we[1]),
    .q      (reg2hw.adaptp_lo_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (adaptp_lo_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.adaptp_lo_thresholds.bypass_thresh.qe = adaptp_lo_thresholds_qe;


  // R[bucket_thresholds]: V(True)
  logic bucket_thresholds_qe;
  logic [1:0] bucket_thresholds_flds_we;
  assign bucket_thresholds_qe = &bucket_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic bucket_thresholds_gated_we;
  assign bucket_thresholds_gated_we = bucket_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_bucket_thresholds_fips_thresh (
    .re     (bucket_thresholds_re),
    .we     (bucket_thresholds_gated_we),
    .wd     (bucket_thresholds_fips_thresh_wd),
    .d      (hw2reg.bucket_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (bucket_thresholds_flds_we[0]),
    .q      (reg2hw.bucket_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (bucket_thresholds_fips_thresh_qs)
  );
  assign reg2hw.bucket_thresholds.fips_thresh.qe = bucket_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_bucket_thresholds_bypass_thresh (
    .re     (bucket_thresholds_re),
    .we     (bucket_thresholds_gated_we),
    .wd     (bucket_thresholds_bypass_thresh_wd),
    .d      (hw2reg.bucket_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (bucket_thresholds_flds_we[1]),
    .q      (reg2hw.bucket_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (bucket_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.bucket_thresholds.bypass_thresh.qe = bucket_thresholds_qe;


  // R[markov_hi_thresholds]: V(True)
  logic markov_hi_thresholds_qe;
  logic [1:0] markov_hi_thresholds_flds_we;
  assign markov_hi_thresholds_qe = &markov_hi_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic markov_hi_thresholds_gated_we;
  assign markov_hi_thresholds_gated_we = markov_hi_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_hi_thresholds_fips_thresh (
    .re     (markov_hi_thresholds_re),
    .we     (markov_hi_thresholds_gated_we),
    .wd     (markov_hi_thresholds_fips_thresh_wd),
    .d      (hw2reg.markov_hi_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (markov_hi_thresholds_flds_we[0]),
    .q      (reg2hw.markov_hi_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (markov_hi_thresholds_fips_thresh_qs)
  );
  assign reg2hw.markov_hi_thresholds.fips_thresh.qe = markov_hi_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_hi_thresholds_bypass_thresh (
    .re     (markov_hi_thresholds_re),
    .we     (markov_hi_thresholds_gated_we),
    .wd     (markov_hi_thresholds_bypass_thresh_wd),
    .d      (hw2reg.markov_hi_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (markov_hi_thresholds_flds_we[1]),
    .q      (reg2hw.markov_hi_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (markov_hi_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.markov_hi_thresholds.bypass_thresh.qe = markov_hi_thresholds_qe;


  // R[markov_lo_thresholds]: V(True)
  logic markov_lo_thresholds_qe;
  logic [1:0] markov_lo_thresholds_flds_we;
  assign markov_lo_thresholds_qe = &markov_lo_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic markov_lo_thresholds_gated_we;
  assign markov_lo_thresholds_gated_we = markov_lo_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_lo_thresholds_fips_thresh (
    .re     (markov_lo_thresholds_re),
    .we     (markov_lo_thresholds_gated_we),
    .wd     (markov_lo_thresholds_fips_thresh_wd),
    .d      (hw2reg.markov_lo_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (markov_lo_thresholds_flds_we[0]),
    .q      (reg2hw.markov_lo_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (markov_lo_thresholds_fips_thresh_qs)
  );
  assign reg2hw.markov_lo_thresholds.fips_thresh.qe = markov_lo_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_lo_thresholds_bypass_thresh (
    .re     (markov_lo_thresholds_re),
    .we     (markov_lo_thresholds_gated_we),
    .wd     (markov_lo_thresholds_bypass_thresh_wd),
    .d      (hw2reg.markov_lo_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (markov_lo_thresholds_flds_we[1]),
    .q      (reg2hw.markov_lo_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (markov_lo_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.markov_lo_thresholds.bypass_thresh.qe = markov_lo_thresholds_qe;


  // R[extht_hi_thresholds]: V(True)
  logic extht_hi_thresholds_qe;
  logic [1:0] extht_hi_thresholds_flds_we;
  assign extht_hi_thresholds_qe = &extht_hi_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic extht_hi_thresholds_gated_we;
  assign extht_hi_thresholds_gated_we = extht_hi_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_hi_thresholds_fips_thresh (
    .re     (extht_hi_thresholds_re),
    .we     (extht_hi_thresholds_gated_we),
    .wd     (extht_hi_thresholds_fips_thresh_wd),
    .d      (hw2reg.extht_hi_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (extht_hi_thresholds_flds_we[0]),
    .q      (reg2hw.extht_hi_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (extht_hi_thresholds_fips_thresh_qs)
  );
  assign reg2hw.extht_hi_thresholds.fips_thresh.qe = extht_hi_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_hi_thresholds_bypass_thresh (
    .re     (extht_hi_thresholds_re),
    .we     (extht_hi_thresholds_gated_we),
    .wd     (extht_hi_thresholds_bypass_thresh_wd),
    .d      (hw2reg.extht_hi_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (extht_hi_thresholds_flds_we[1]),
    .q      (reg2hw.extht_hi_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (extht_hi_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.extht_hi_thresholds.bypass_thresh.qe = extht_hi_thresholds_qe;


  // R[extht_lo_thresholds]: V(True)
  logic extht_lo_thresholds_qe;
  logic [1:0] extht_lo_thresholds_flds_we;
  assign extht_lo_thresholds_qe = &extht_lo_thresholds_flds_we;
  // Create REGWEN-gated WE signal
  logic extht_lo_thresholds_gated_we;
  assign extht_lo_thresholds_gated_we = extht_lo_thresholds_we & regwen_qs;
  //   F[fips_thresh]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_lo_thresholds_fips_thresh (
    .re     (extht_lo_thresholds_re),
    .we     (extht_lo_thresholds_gated_we),
    .wd     (extht_lo_thresholds_fips_thresh_wd),
    .d      (hw2reg.extht_lo_thresholds.fips_thresh.d),
    .qre    (),
    .qe     (extht_lo_thresholds_flds_we[0]),
    .q      (reg2hw.extht_lo_thresholds.fips_thresh.q),
    .ds     (),
    .qs     (extht_lo_thresholds_fips_thresh_qs)
  );
  assign reg2hw.extht_lo_thresholds.fips_thresh.qe = extht_lo_thresholds_qe;

  //   F[bypass_thresh]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_lo_thresholds_bypass_thresh (
    .re     (extht_lo_thresholds_re),
    .we     (extht_lo_thresholds_gated_we),
    .wd     (extht_lo_thresholds_bypass_thresh_wd),
    .d      (hw2reg.extht_lo_thresholds.bypass_thresh.d),
    .qre    (),
    .qe     (extht_lo_thresholds_flds_we[1]),
    .q      (reg2hw.extht_lo_thresholds.bypass_thresh.q),
    .ds     (),
    .qs     (extht_lo_thresholds_bypass_thresh_qs)
  );
  assign reg2hw.extht_lo_thresholds.bypass_thresh.qe = extht_lo_thresholds_qe;


  // R[repcnt_hi_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnt_hi_watermarks_fips_watermark (
    .re     (repcnt_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.repcnt_hi_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (repcnt_hi_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnt_hi_watermarks_bypass_watermark (
    .re     (repcnt_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.repcnt_hi_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (repcnt_hi_watermarks_bypass_watermark_qs)
  );


  // R[repcnts_hi_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnts_hi_watermarks_fips_watermark (
    .re     (repcnts_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.repcnts_hi_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (repcnts_hi_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_repcnts_hi_watermarks_bypass_watermark (
    .re     (repcnts_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.repcnts_hi_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (repcnts_hi_watermarks_bypass_watermark_qs)
  );


  // R[adaptp_hi_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_hi_watermarks_fips_watermark (
    .re     (adaptp_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.adaptp_hi_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (adaptp_hi_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_hi_watermarks_bypass_watermark (
    .re     (adaptp_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.adaptp_hi_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (adaptp_hi_watermarks_bypass_watermark_qs)
  );


  // R[adaptp_lo_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_lo_watermarks_fips_watermark (
    .re     (adaptp_lo_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.adaptp_lo_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (adaptp_lo_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_adaptp_lo_watermarks_bypass_watermark (
    .re     (adaptp_lo_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.adaptp_lo_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (adaptp_lo_watermarks_bypass_watermark_qs)
  );


  // R[extht_hi_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_hi_watermarks_fips_watermark (
    .re     (extht_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_hi_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_hi_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_hi_watermarks_bypass_watermark (
    .re     (extht_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_hi_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_hi_watermarks_bypass_watermark_qs)
  );


  // R[extht_lo_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_lo_watermarks_fips_watermark (
    .re     (extht_lo_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_lo_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_lo_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_extht_lo_watermarks_bypass_watermark (
    .re     (extht_lo_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_lo_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_lo_watermarks_bypass_watermark_qs)
  );


  // R[bucket_hi_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_bucket_hi_watermarks_fips_watermark (
    .re     (bucket_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.bucket_hi_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (bucket_hi_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_bucket_hi_watermarks_bypass_watermark (
    .re     (bucket_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.bucket_hi_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (bucket_hi_watermarks_bypass_watermark_qs)
  );


  // R[markov_hi_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_hi_watermarks_fips_watermark (
    .re     (markov_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.markov_hi_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (markov_hi_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_hi_watermarks_bypass_watermark (
    .re     (markov_hi_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.markov_hi_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (markov_hi_watermarks_bypass_watermark_qs)
  );


  // R[markov_lo_watermarks]: V(True)
  //   F[fips_watermark]: 15:0
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_lo_watermarks_fips_watermark (
    .re     (markov_lo_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.markov_lo_watermarks.fips_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (markov_lo_watermarks_fips_watermark_qs)
  );

  //   F[bypass_watermark]: 31:16
  prim_subreg_ext #(
    .DW    (16)
  ) u_markov_lo_watermarks_bypass_watermark (
    .re     (markov_lo_watermarks_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.markov_lo_watermarks.bypass_watermark.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (markov_lo_watermarks_bypass_watermark_qs)
  );


  // R[repcnt_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_repcnt_total_fails (
    .re     (repcnt_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.repcnt_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (repcnt_total_fails_qs)
  );


  // R[repcnts_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_repcnts_total_fails (
    .re     (repcnts_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.repcnts_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (repcnts_total_fails_qs)
  );


  // R[adaptp_hi_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_adaptp_hi_total_fails (
    .re     (adaptp_hi_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.adaptp_hi_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (adaptp_hi_total_fails_qs)
  );


  // R[adaptp_lo_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_adaptp_lo_total_fails (
    .re     (adaptp_lo_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.adaptp_lo_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (adaptp_lo_total_fails_qs)
  );


  // R[bucket_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_bucket_total_fails (
    .re     (bucket_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.bucket_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (bucket_total_fails_qs)
  );


  // R[markov_hi_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_markov_hi_total_fails (
    .re     (markov_hi_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.markov_hi_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (markov_hi_total_fails_qs)
  );


  // R[markov_lo_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_markov_lo_total_fails (
    .re     (markov_lo_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.markov_lo_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (markov_lo_total_fails_qs)
  );


  // R[extht_hi_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_extht_hi_total_fails (
    .re     (extht_hi_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_hi_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_hi_total_fails_qs)
  );


  // R[extht_lo_total_fails]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_extht_lo_total_fails (
    .re     (extht_lo_total_fails_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_lo_total_fails.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_lo_total_fails_qs)
  );


  // R[alert_threshold]: V(False)
  // Create REGWEN-gated WE signal
  logic alert_threshold_gated_we;
  assign alert_threshold_gated_we = alert_threshold_we & regwen_qs;
  //   F[alert_threshold]: 15:0
  prim_subreg #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h2)
  ) u_alert_threshold_alert_threshold (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (alert_threshold_gated_we),
    .wd     (alert_threshold_alert_threshold_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.alert_threshold.alert_threshold.q),
    .ds     (),

    // to register interface (read)
    .qs     (alert_threshold_alert_threshold_qs)
  );

  //   F[alert_threshold_inv]: 31:16
  prim_subreg #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'hfffd)
  ) u_alert_threshold_alert_threshold_inv (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (alert_threshold_gated_we),
    .wd     (alert_threshold_alert_threshold_inv_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.alert_threshold.alert_threshold_inv.q),
    .ds     (),

    // to register interface (read)
    .qs     (alert_threshold_alert_threshold_inv_qs)
  );


  // R[alert_summary_fail_counts]: V(True)
  prim_subreg_ext #(
    .DW    (16)
  ) u_alert_summary_fail_counts (
    .re     (alert_summary_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_summary_fail_counts.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_summary_fail_counts_qs)
  );


  // R[alert_fail_counts]: V(True)
  //   F[repcnt_fail_count]: 7:4
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_repcnt_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.repcnt_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_repcnt_fail_count_qs)
  );

  //   F[adaptp_hi_fail_count]: 11:8
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_adaptp_hi_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.adaptp_hi_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_adaptp_hi_fail_count_qs)
  );

  //   F[adaptp_lo_fail_count]: 15:12
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_adaptp_lo_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.adaptp_lo_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_adaptp_lo_fail_count_qs)
  );

  //   F[bucket_fail_count]: 19:16
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_bucket_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.bucket_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_bucket_fail_count_qs)
  );

  //   F[markov_hi_fail_count]: 23:20
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_markov_hi_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.markov_hi_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_markov_hi_fail_count_qs)
  );

  //   F[markov_lo_fail_count]: 27:24
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_markov_lo_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.markov_lo_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_markov_lo_fail_count_qs)
  );

  //   F[repcnts_fail_count]: 31:28
  prim_subreg_ext #(
    .DW    (4)
  ) u_alert_fail_counts_repcnts_fail_count (
    .re     (alert_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.alert_fail_counts.repcnts_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (alert_fail_counts_repcnts_fail_count_qs)
  );


  // R[extht_fail_counts]: V(True)
  //   F[extht_hi_fail_count]: 3:0
  prim_subreg_ext #(
    .DW    (4)
  ) u_extht_fail_counts_extht_hi_fail_count (
    .re     (extht_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_fail_counts.extht_hi_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_fail_counts_extht_hi_fail_count_qs)
  );

  //   F[extht_lo_fail_count]: 7:4
  prim_subreg_ext #(
    .DW    (4)
  ) u_extht_fail_counts_extht_lo_fail_count (
    .re     (extht_fail_counts_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.extht_fail_counts.extht_lo_fail_count.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (extht_fail_counts_extht_lo_fail_count_qs)
  );


  // R[fw_ov_control]: V(False)
  // Create REGWEN-gated WE signal
  logic fw_ov_control_gated_we;
  assign fw_ov_control_gated_we = fw_ov_control_we & regwen_qs;
  //   F[fw_ov_mode]: 3:0
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_fw_ov_control_fw_ov_mode (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (fw_ov_control_gated_we),
    .wd     (fw_ov_control_fw_ov_mode_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fw_ov_control.fw_ov_mode.q),
    .ds     (),

    // to register interface (read)
    .qs     (fw_ov_control_fw_ov_mode_qs)
  );

  //   F[fw_ov_entropy_insert]: 7:4
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_fw_ov_control_fw_ov_entropy_insert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (fw_ov_control_gated_we),
    .wd     (fw_ov_control_fw_ov_entropy_insert_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fw_ov_control.fw_ov_entropy_insert.q),
    .ds     (),

    // to register interface (read)
    .qs     (fw_ov_control_fw_ov_entropy_insert_qs)
  );


  // R[fw_ov_sha3_start]: V(False)
  prim_subreg #(
    .DW      (4),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (4'h9)
  ) u_fw_ov_sha3_start (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (fw_ov_sha3_start_we),
    .wd     (fw_ov_sha3_start_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fw_ov_sha3_start.q),
    .ds     (),

    // to register interface (read)
    .qs     (fw_ov_sha3_start_qs)
  );


  // R[fw_ov_wr_fifo_full]: V(True)
  prim_subreg_ext #(
    .DW    (1)
  ) u_fw_ov_wr_fifo_full (
    .re     (fw_ov_wr_fifo_full_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.fw_ov_wr_fifo_full.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (fw_ov_wr_fifo_full_qs)
  );


  // R[fw_ov_rd_fifo_overflow]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_fw_ov_rd_fifo_overflow (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (fw_ov_rd_fifo_overflow_we),
    .wd     (fw_ov_rd_fifo_overflow_wd),

    // from internal hardware
    .de     (hw2reg.fw_ov_rd_fifo_overflow.de),
    .d      (hw2reg.fw_ov_rd_fifo_overflow.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fw_ov_rd_fifo_overflow_qs)
  );


  // R[fw_ov_rd_data]: V(True)
  prim_subreg_ext #(
    .DW    (32)
  ) u_fw_ov_rd_data (
    .re     (fw_ov_rd_data_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.fw_ov_rd_data.d),
    .qre    (reg2hw.fw_ov_rd_data.re),
    .qe     (),
    .q      (reg2hw.fw_ov_rd_data.q),
    .ds     (),
    .qs     (fw_ov_rd_data_qs)
  );


  // R[fw_ov_wr_data]: V(True)
  logic fw_ov_wr_data_qe;
  logic [0:0] fw_ov_wr_data_flds_we;
  assign fw_ov_wr_data_qe = &fw_ov_wr_data_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_fw_ov_wr_data (
    .re     (1'b0),
    .we     (fw_ov_wr_data_we),
    .wd     (fw_ov_wr_data_wd),
    .d      ('0),
    .qre    (),
    .qe     (fw_ov_wr_data_flds_we[0]),
    .q      (reg2hw.fw_ov_wr_data.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.fw_ov_wr_data.qe = fw_ov_wr_data_qe;


  // R[observe_fifo_thresh]: V(False)
  // Create REGWEN-gated WE signal
  logic observe_fifo_thresh_gated_we;
  assign observe_fifo_thresh_gated_we = observe_fifo_thresh_we & regwen_qs;
  prim_subreg #(
    .DW      (7),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (7'h20)
  ) u_observe_fifo_thresh (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (observe_fifo_thresh_gated_we),
    .wd     (observe_fifo_thresh_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.observe_fifo_thresh.q),
    .ds     (),

    // to register interface (read)
    .qs     (observe_fifo_thresh_qs)
  );


  // R[observe_fifo_depth]: V(True)
  prim_subreg_ext #(
    .DW    (7)
  ) u_observe_fifo_depth (
    .re     (observe_fifo_depth_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.observe_fifo_depth.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (observe_fifo_depth_qs)
  );


  // R[debug_status]: V(True)
  //   F[entropy_fifo_depth]: 2:0
  prim_subreg_ext #(
    .DW    (3)
  ) u_debug_status_entropy_fifo_depth (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.entropy_fifo_depth.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_entropy_fifo_depth_qs)
  );

  //   F[sha3_fsm]: 5:3
  prim_subreg_ext #(
    .DW    (3)
  ) u_debug_status_sha3_fsm (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.sha3_fsm.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_sha3_fsm_qs)
  );

  //   F[sha3_block_pr]: 6:6
  prim_subreg_ext #(
    .DW    (1)
  ) u_debug_status_sha3_block_pr (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.sha3_block_pr.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_sha3_block_pr_qs)
  );

  //   F[sha3_squeezing]: 7:7
  prim_subreg_ext #(
    .DW    (1)
  ) u_debug_status_sha3_squeezing (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.sha3_squeezing.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_sha3_squeezing_qs)
  );

  //   F[sha3_absorbed]: 8:8
  prim_subreg_ext #(
    .DW    (1)
  ) u_debug_status_sha3_absorbed (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.sha3_absorbed.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_sha3_absorbed_qs)
  );

  //   F[sha3_err]: 9:9
  prim_subreg_ext #(
    .DW    (1)
  ) u_debug_status_sha3_err (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.sha3_err.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_sha3_err_qs)
  );

  //   F[main_sm_idle]: 16:16
  prim_subreg_ext #(
    .DW    (1)
  ) u_debug_status_main_sm_idle (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.main_sm_idle.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_main_sm_idle_qs)
  );

  //   F[main_sm_boot_done]: 17:17
  prim_subreg_ext #(
    .DW    (1)
  ) u_debug_status_main_sm_boot_done (
    .re     (debug_status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.debug_status.main_sm_boot_done.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (debug_status_main_sm_boot_done_qs)
  );


  // R[recov_alert_sts]: V(False)
  //   F[fips_enable_field_alert]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_fips_enable_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_fips_enable_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.fips_enable_field_alert.de),
    .d      (hw2reg.recov_alert_sts.fips_enable_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_fips_enable_field_alert_qs)
  );

  //   F[entropy_data_reg_en_field_alert]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_entropy_data_reg_en_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_entropy_data_reg_en_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.entropy_data_reg_en_field_alert.de),
    .d      (hw2reg.recov_alert_sts.entropy_data_reg_en_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_entropy_data_reg_en_field_alert_qs)
  );

  //   F[module_enable_field_alert]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_module_enable_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_module_enable_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.module_enable_field_alert.de),
    .d      (hw2reg.recov_alert_sts.module_enable_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_module_enable_field_alert_qs)
  );

  //   F[threshold_scope_field_alert]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_threshold_scope_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_threshold_scope_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.threshold_scope_field_alert.de),
    .d      (hw2reg.recov_alert_sts.threshold_scope_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_threshold_scope_field_alert_qs)
  );

  //   F[rng_bit_enable_field_alert]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_rng_bit_enable_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_rng_bit_enable_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.rng_bit_enable_field_alert.de),
    .d      (hw2reg.recov_alert_sts.rng_bit_enable_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_rng_bit_enable_field_alert_qs)
  );

  //   F[fw_ov_sha3_start_field_alert]: 7:7
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_fw_ov_sha3_start_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_fw_ov_sha3_start_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.fw_ov_sha3_start_field_alert.de),
    .d      (hw2reg.recov_alert_sts.fw_ov_sha3_start_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_fw_ov_sha3_start_field_alert_qs)
  );

  //   F[fw_ov_mode_field_alert]: 8:8
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_fw_ov_mode_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_fw_ov_mode_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.fw_ov_mode_field_alert.de),
    .d      (hw2reg.recov_alert_sts.fw_ov_mode_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_fw_ov_mode_field_alert_qs)
  );

  //   F[fw_ov_entropy_insert_field_alert]: 9:9
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_fw_ov_entropy_insert_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_fw_ov_entropy_insert_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.fw_ov_entropy_insert_field_alert.de),
    .d      (hw2reg.recov_alert_sts.fw_ov_entropy_insert_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_fw_ov_entropy_insert_field_alert_qs)
  );

  //   F[es_route_field_alert]: 10:10
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_route_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_route_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_route_field_alert.de),
    .d      (hw2reg.recov_alert_sts.es_route_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_route_field_alert_qs)
  );

  //   F[es_type_field_alert]: 11:11
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_type_field_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_type_field_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_type_field_alert.de),
    .d      (hw2reg.recov_alert_sts.es_type_field_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_type_field_alert_qs)
  );

  //   F[es_main_sm_alert]: 12:12
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_main_sm_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_main_sm_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_main_sm_alert.de),
    .d      (hw2reg.recov_alert_sts.es_main_sm_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_main_sm_alert_qs)
  );

  //   F[es_bus_cmp_alert]: 13:13
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_bus_cmp_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_bus_cmp_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_bus_cmp_alert.de),
    .d      (hw2reg.recov_alert_sts.es_bus_cmp_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_bus_cmp_alert_qs)
  );

  //   F[es_thresh_cfg_alert]: 14:14
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_thresh_cfg_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_thresh_cfg_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_thresh_cfg_alert.de),
    .d      (hw2reg.recov_alert_sts.es_thresh_cfg_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_thresh_cfg_alert_qs)
  );

  //   F[es_fw_ov_wr_alert]: 15:15
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_fw_ov_wr_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_fw_ov_wr_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_fw_ov_wr_alert.de),
    .d      (hw2reg.recov_alert_sts.es_fw_ov_wr_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_fw_ov_wr_alert_qs)
  );

  //   F[es_fw_ov_disable_alert]: 16:16
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_recov_alert_sts_es_fw_ov_disable_alert (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (recov_alert_sts_we),
    .wd     (recov_alert_sts_es_fw_ov_disable_alert_wd),

    // from internal hardware
    .de     (hw2reg.recov_alert_sts.es_fw_ov_disable_alert.de),
    .d      (hw2reg.recov_alert_sts.es_fw_ov_disable_alert.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (recov_alert_sts_es_fw_ov_disable_alert_qs)
  );


  // R[err_code]: V(False)
  //   F[sfifo_esrng_err]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_esrng_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_esrng_err.de),
    .d      (hw2reg.err_code.sfifo_esrng_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_esrng_err_qs)
  );

  //   F[sfifo_observe_err]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_observe_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_observe_err.de),
    .d      (hw2reg.err_code.sfifo_observe_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_observe_err_qs)
  );

  //   F[sfifo_esfinal_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sfifo_esfinal_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sfifo_esfinal_err.de),
    .d      (hw2reg.err_code.sfifo_esfinal_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sfifo_esfinal_err_qs)
  );

  //   F[es_ack_sm_err]: 20:20
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_es_ack_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.es_ack_sm_err.de),
    .d      (hw2reg.err_code.es_ack_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_es_ack_sm_err_qs)
  );

  //   F[es_main_sm_err]: 21:21
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_es_main_sm_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.es_main_sm_err.de),
    .d      (hw2reg.err_code.es_main_sm_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_es_main_sm_err_qs)
  );

  //   F[es_cntr_err]: 22:22
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_es_cntr_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.es_cntr_err.de),
    .d      (hw2reg.err_code.es_cntr_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_es_cntr_err_qs)
  );

  //   F[sha3_state_err]: 23:23
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sha3_state_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sha3_state_err.de),
    .d      (hw2reg.err_code.sha3_state_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sha3_state_err_qs)
  );

  //   F[sha3_rst_storage_err]: 24:24
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_sha3_rst_storage_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.sha3_rst_storage_err.de),
    .d      (hw2reg.err_code.sha3_rst_storage_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_sha3_rst_storage_err_qs)
  );

  //   F[fifo_write_err]: 28:28
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_write_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_write_err.de),
    .d      (hw2reg.err_code.fifo_write_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_write_err_qs)
  );

  //   F[fifo_read_err]: 29:29
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_read_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_read_err.de),
    .d      (hw2reg.err_code.fifo_read_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_read_err_qs)
  );

  //   F[fifo_state_err]: 30:30
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_err_code_fifo_state_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.fifo_state_err.de),
    .d      (hw2reg.err_code.fifo_state_err.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_fifo_state_err_qs)
  );


  // R[err_code_test]: V(False)
  logic err_code_test_qe;
  logic [0:0] err_code_test_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_err_code_test0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&err_code_test_flds_we),
    .q_o(err_code_test_qe)
  );
  prim_subreg #(
    .DW      (5),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (5'h0)
  ) u_err_code_test (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (err_code_test_we),
    .wd     (err_code_test_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (err_code_test_flds_we[0]),
    .q      (reg2hw.err_code_test.q),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_test_qs)
  );
  assign reg2hw.err_code_test.qe = err_code_test_qe;


  // R[main_sm_state]: V(False)
  prim_subreg #(
    .DW      (9),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (9'hf5)
  ) u_main_sm_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.main_sm_state.de),
    .d      (hw2reg.main_sm_state.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (main_sm_state_qs)
  );



  logic [56:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == ENTROPY_SRC_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == ENTROPY_SRC_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == ENTROPY_SRC_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == ENTROPY_SRC_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == ENTROPY_SRC_ME_REGWEN_OFFSET);
    addr_hit[ 5] = (reg_addr == ENTROPY_SRC_SW_REGUPD_OFFSET);
    addr_hit[ 6] = (reg_addr == ENTROPY_SRC_REGWEN_OFFSET);
    addr_hit[ 7] = (reg_addr == ENTROPY_SRC_REV_OFFSET);
    addr_hit[ 8] = (reg_addr == ENTROPY_SRC_MODULE_ENABLE_OFFSET);
    addr_hit[ 9] = (reg_addr == ENTROPY_SRC_CONF_OFFSET);
    addr_hit[10] = (reg_addr == ENTROPY_SRC_ENTROPY_CONTROL_OFFSET);
    addr_hit[11] = (reg_addr == ENTROPY_SRC_ENTROPY_DATA_OFFSET);
    addr_hit[12] = (reg_addr == ENTROPY_SRC_HEALTH_TEST_WINDOWS_OFFSET);
    addr_hit[13] = (reg_addr == ENTROPY_SRC_REPCNT_THRESHOLDS_OFFSET);
    addr_hit[14] = (reg_addr == ENTROPY_SRC_REPCNTS_THRESHOLDS_OFFSET);
    addr_hit[15] = (reg_addr == ENTROPY_SRC_ADAPTP_HI_THRESHOLDS_OFFSET);
    addr_hit[16] = (reg_addr == ENTROPY_SRC_ADAPTP_LO_THRESHOLDS_OFFSET);
    addr_hit[17] = (reg_addr == ENTROPY_SRC_BUCKET_THRESHOLDS_OFFSET);
    addr_hit[18] = (reg_addr == ENTROPY_SRC_MARKOV_HI_THRESHOLDS_OFFSET);
    addr_hit[19] = (reg_addr == ENTROPY_SRC_MARKOV_LO_THRESHOLDS_OFFSET);
    addr_hit[20] = (reg_addr == ENTROPY_SRC_EXTHT_HI_THRESHOLDS_OFFSET);
    addr_hit[21] = (reg_addr == ENTROPY_SRC_EXTHT_LO_THRESHOLDS_OFFSET);
    addr_hit[22] = (reg_addr == ENTROPY_SRC_REPCNT_HI_WATERMARKS_OFFSET);
    addr_hit[23] = (reg_addr == ENTROPY_SRC_REPCNTS_HI_WATERMARKS_OFFSET);
    addr_hit[24] = (reg_addr == ENTROPY_SRC_ADAPTP_HI_WATERMARKS_OFFSET);
    addr_hit[25] = (reg_addr == ENTROPY_SRC_ADAPTP_LO_WATERMARKS_OFFSET);
    addr_hit[26] = (reg_addr == ENTROPY_SRC_EXTHT_HI_WATERMARKS_OFFSET);
    addr_hit[27] = (reg_addr == ENTROPY_SRC_EXTHT_LO_WATERMARKS_OFFSET);
    addr_hit[28] = (reg_addr == ENTROPY_SRC_BUCKET_HI_WATERMARKS_OFFSET);
    addr_hit[29] = (reg_addr == ENTROPY_SRC_MARKOV_HI_WATERMARKS_OFFSET);
    addr_hit[30] = (reg_addr == ENTROPY_SRC_MARKOV_LO_WATERMARKS_OFFSET);
    addr_hit[31] = (reg_addr == ENTROPY_SRC_REPCNT_TOTAL_FAILS_OFFSET);
    addr_hit[32] = (reg_addr == ENTROPY_SRC_REPCNTS_TOTAL_FAILS_OFFSET);
    addr_hit[33] = (reg_addr == ENTROPY_SRC_ADAPTP_HI_TOTAL_FAILS_OFFSET);
    addr_hit[34] = (reg_addr == ENTROPY_SRC_ADAPTP_LO_TOTAL_FAILS_OFFSET);
    addr_hit[35] = (reg_addr == ENTROPY_SRC_BUCKET_TOTAL_FAILS_OFFSET);
    addr_hit[36] = (reg_addr == ENTROPY_SRC_MARKOV_HI_TOTAL_FAILS_OFFSET);
    addr_hit[37] = (reg_addr == ENTROPY_SRC_MARKOV_LO_TOTAL_FAILS_OFFSET);
    addr_hit[38] = (reg_addr == ENTROPY_SRC_EXTHT_HI_TOTAL_FAILS_OFFSET);
    addr_hit[39] = (reg_addr == ENTROPY_SRC_EXTHT_LO_TOTAL_FAILS_OFFSET);
    addr_hit[40] = (reg_addr == ENTROPY_SRC_ALERT_THRESHOLD_OFFSET);
    addr_hit[41] = (reg_addr == ENTROPY_SRC_ALERT_SUMMARY_FAIL_COUNTS_OFFSET);
    addr_hit[42] = (reg_addr == ENTROPY_SRC_ALERT_FAIL_COUNTS_OFFSET);
    addr_hit[43] = (reg_addr == ENTROPY_SRC_EXTHT_FAIL_COUNTS_OFFSET);
    addr_hit[44] = (reg_addr == ENTROPY_SRC_FW_OV_CONTROL_OFFSET);
    addr_hit[45] = (reg_addr == ENTROPY_SRC_FW_OV_SHA3_START_OFFSET);
    addr_hit[46] = (reg_addr == ENTROPY_SRC_FW_OV_WR_FIFO_FULL_OFFSET);
    addr_hit[47] = (reg_addr == ENTROPY_SRC_FW_OV_RD_FIFO_OVERFLOW_OFFSET);
    addr_hit[48] = (reg_addr == ENTROPY_SRC_FW_OV_RD_DATA_OFFSET);
    addr_hit[49] = (reg_addr == ENTROPY_SRC_FW_OV_WR_DATA_OFFSET);
    addr_hit[50] = (reg_addr == ENTROPY_SRC_OBSERVE_FIFO_THRESH_OFFSET);
    addr_hit[51] = (reg_addr == ENTROPY_SRC_OBSERVE_FIFO_DEPTH_OFFSET);
    addr_hit[52] = (reg_addr == ENTROPY_SRC_DEBUG_STATUS_OFFSET);
    addr_hit[53] = (reg_addr == ENTROPY_SRC_RECOV_ALERT_STS_OFFSET);
    addr_hit[54] = (reg_addr == ENTROPY_SRC_ERR_CODE_OFFSET);
    addr_hit[55] = (reg_addr == ENTROPY_SRC_ERR_CODE_TEST_OFFSET);
    addr_hit[56] = (reg_addr == ENTROPY_SRC_MAIN_SM_STATE_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(ENTROPY_SRC_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(ENTROPY_SRC_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(ENTROPY_SRC_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(ENTROPY_SRC_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(ENTROPY_SRC_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(ENTROPY_SRC_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(ENTROPY_SRC_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(ENTROPY_SRC_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(ENTROPY_SRC_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(ENTROPY_SRC_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(ENTROPY_SRC_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(ENTROPY_SRC_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(ENTROPY_SRC_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(ENTROPY_SRC_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(ENTROPY_SRC_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(ENTROPY_SRC_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(ENTROPY_SRC_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(ENTROPY_SRC_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(ENTROPY_SRC_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(ENTROPY_SRC_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(ENTROPY_SRC_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(ENTROPY_SRC_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(ENTROPY_SRC_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(ENTROPY_SRC_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(ENTROPY_SRC_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(ENTROPY_SRC_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(ENTROPY_SRC_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(ENTROPY_SRC_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(ENTROPY_SRC_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(ENTROPY_SRC_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(ENTROPY_SRC_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(ENTROPY_SRC_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(ENTROPY_SRC_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(ENTROPY_SRC_PERMIT[33] & ~reg_be))) |
               (addr_hit[34] & (|(ENTROPY_SRC_PERMIT[34] & ~reg_be))) |
               (addr_hit[35] & (|(ENTROPY_SRC_PERMIT[35] & ~reg_be))) |
               (addr_hit[36] & (|(ENTROPY_SRC_PERMIT[36] & ~reg_be))) |
               (addr_hit[37] & (|(ENTROPY_SRC_PERMIT[37] & ~reg_be))) |
               (addr_hit[38] & (|(ENTROPY_SRC_PERMIT[38] & ~reg_be))) |
               (addr_hit[39] & (|(ENTROPY_SRC_PERMIT[39] & ~reg_be))) |
               (addr_hit[40] & (|(ENTROPY_SRC_PERMIT[40] & ~reg_be))) |
               (addr_hit[41] & (|(ENTROPY_SRC_PERMIT[41] & ~reg_be))) |
               (addr_hit[42] & (|(ENTROPY_SRC_PERMIT[42] & ~reg_be))) |
               (addr_hit[43] & (|(ENTROPY_SRC_PERMIT[43] & ~reg_be))) |
               (addr_hit[44] & (|(ENTROPY_SRC_PERMIT[44] & ~reg_be))) |
               (addr_hit[45] & (|(ENTROPY_SRC_PERMIT[45] & ~reg_be))) |
               (addr_hit[46] & (|(ENTROPY_SRC_PERMIT[46] & ~reg_be))) |
               (addr_hit[47] & (|(ENTROPY_SRC_PERMIT[47] & ~reg_be))) |
               (addr_hit[48] & (|(ENTROPY_SRC_PERMIT[48] & ~reg_be))) |
               (addr_hit[49] & (|(ENTROPY_SRC_PERMIT[49] & ~reg_be))) |
               (addr_hit[50] & (|(ENTROPY_SRC_PERMIT[50] & ~reg_be))) |
               (addr_hit[51] & (|(ENTROPY_SRC_PERMIT[51] & ~reg_be))) |
               (addr_hit[52] & (|(ENTROPY_SRC_PERMIT[52] & ~reg_be))) |
               (addr_hit[53] & (|(ENTROPY_SRC_PERMIT[53] & ~reg_be))) |
               (addr_hit[54] & (|(ENTROPY_SRC_PERMIT[54] & ~reg_be))) |
               (addr_hit[55] & (|(ENTROPY_SRC_PERMIT[55] & ~reg_be))) |
               (addr_hit[56] & (|(ENTROPY_SRC_PERMIT[56] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_es_entropy_valid_wd = reg_wdata[0];

  assign intr_state_es_health_test_failed_wd = reg_wdata[1];

  assign intr_state_es_observe_fifo_ready_wd = reg_wdata[2];

  assign intr_state_es_fatal_err_wd = reg_wdata[3];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_es_entropy_valid_wd = reg_wdata[0];

  assign intr_enable_es_health_test_failed_wd = reg_wdata[1];

  assign intr_enable_es_observe_fifo_ready_wd = reg_wdata[2];

  assign intr_enable_es_fatal_err_wd = reg_wdata[3];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_es_entropy_valid_wd = reg_wdata[0];

  assign intr_test_es_health_test_failed_wd = reg_wdata[1];

  assign intr_test_es_observe_fifo_ready_wd = reg_wdata[2];

  assign intr_test_es_fatal_err_wd = reg_wdata[3];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_recov_alert_wd = reg_wdata[0];

  assign alert_test_fatal_alert_wd = reg_wdata[1];
  assign me_regwen_we = addr_hit[4] & reg_we & !reg_error;

  assign me_regwen_wd = reg_wdata[0];
  assign sw_regupd_we = addr_hit[5] & reg_we & !reg_error;

  assign sw_regupd_wd = reg_wdata[0];
  assign module_enable_we = addr_hit[8] & reg_we & !reg_error;

  assign module_enable_wd = reg_wdata[3:0];
  assign conf_we = addr_hit[9] & reg_we & !reg_error;

  assign conf_fips_enable_wd = reg_wdata[3:0];

  assign conf_entropy_data_reg_enable_wd = reg_wdata[7:4];

  assign conf_threshold_scope_wd = reg_wdata[15:12];

  assign conf_rng_bit_enable_wd = reg_wdata[23:20];

  assign conf_rng_bit_sel_wd = reg_wdata[25:24];
  assign entropy_control_we = addr_hit[10] & reg_we & !reg_error;

  assign entropy_control_es_route_wd = reg_wdata[3:0];

  assign entropy_control_es_type_wd = reg_wdata[7:4];
  assign entropy_data_re = addr_hit[11] & reg_re & !reg_error;
  assign health_test_windows_we = addr_hit[12] & reg_we & !reg_error;

  assign health_test_windows_fips_window_wd = reg_wdata[15:0];

  assign health_test_windows_bypass_window_wd = reg_wdata[31:16];
  assign repcnt_thresholds_re = addr_hit[13] & reg_re & !reg_error;
  assign repcnt_thresholds_we = addr_hit[13] & reg_we & !reg_error;

  assign repcnt_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign repcnt_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign repcnts_thresholds_re = addr_hit[14] & reg_re & !reg_error;
  assign repcnts_thresholds_we = addr_hit[14] & reg_we & !reg_error;

  assign repcnts_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign repcnts_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign adaptp_hi_thresholds_re = addr_hit[15] & reg_re & !reg_error;
  assign adaptp_hi_thresholds_we = addr_hit[15] & reg_we & !reg_error;

  assign adaptp_hi_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign adaptp_hi_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign adaptp_lo_thresholds_re = addr_hit[16] & reg_re & !reg_error;
  assign adaptp_lo_thresholds_we = addr_hit[16] & reg_we & !reg_error;

  assign adaptp_lo_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign adaptp_lo_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign bucket_thresholds_re = addr_hit[17] & reg_re & !reg_error;
  assign bucket_thresholds_we = addr_hit[17] & reg_we & !reg_error;

  assign bucket_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign bucket_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign markov_hi_thresholds_re = addr_hit[18] & reg_re & !reg_error;
  assign markov_hi_thresholds_we = addr_hit[18] & reg_we & !reg_error;

  assign markov_hi_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign markov_hi_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign markov_lo_thresholds_re = addr_hit[19] & reg_re & !reg_error;
  assign markov_lo_thresholds_we = addr_hit[19] & reg_we & !reg_error;

  assign markov_lo_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign markov_lo_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign extht_hi_thresholds_re = addr_hit[20] & reg_re & !reg_error;
  assign extht_hi_thresholds_we = addr_hit[20] & reg_we & !reg_error;

  assign extht_hi_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign extht_hi_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign extht_lo_thresholds_re = addr_hit[21] & reg_re & !reg_error;
  assign extht_lo_thresholds_we = addr_hit[21] & reg_we & !reg_error;

  assign extht_lo_thresholds_fips_thresh_wd = reg_wdata[15:0];

  assign extht_lo_thresholds_bypass_thresh_wd = reg_wdata[31:16];
  assign repcnt_hi_watermarks_re = addr_hit[22] & reg_re & !reg_error;
  assign repcnts_hi_watermarks_re = addr_hit[23] & reg_re & !reg_error;
  assign adaptp_hi_watermarks_re = addr_hit[24] & reg_re & !reg_error;
  assign adaptp_lo_watermarks_re = addr_hit[25] & reg_re & !reg_error;
  assign extht_hi_watermarks_re = addr_hit[26] & reg_re & !reg_error;
  assign extht_lo_watermarks_re = addr_hit[27] & reg_re & !reg_error;
  assign bucket_hi_watermarks_re = addr_hit[28] & reg_re & !reg_error;
  assign markov_hi_watermarks_re = addr_hit[29] & reg_re & !reg_error;
  assign markov_lo_watermarks_re = addr_hit[30] & reg_re & !reg_error;
  assign repcnt_total_fails_re = addr_hit[31] & reg_re & !reg_error;
  assign repcnts_total_fails_re = addr_hit[32] & reg_re & !reg_error;
  assign adaptp_hi_total_fails_re = addr_hit[33] & reg_re & !reg_error;
  assign adaptp_lo_total_fails_re = addr_hit[34] & reg_re & !reg_error;
  assign bucket_total_fails_re = addr_hit[35] & reg_re & !reg_error;
  assign markov_hi_total_fails_re = addr_hit[36] & reg_re & !reg_error;
  assign markov_lo_total_fails_re = addr_hit[37] & reg_re & !reg_error;
  assign extht_hi_total_fails_re = addr_hit[38] & reg_re & !reg_error;
  assign extht_lo_total_fails_re = addr_hit[39] & reg_re & !reg_error;
  assign alert_threshold_we = addr_hit[40] & reg_we & !reg_error;

  assign alert_threshold_alert_threshold_wd = reg_wdata[15:0];

  assign alert_threshold_alert_threshold_inv_wd = reg_wdata[31:16];
  assign alert_summary_fail_counts_re = addr_hit[41] & reg_re & !reg_error;
  assign alert_fail_counts_re = addr_hit[42] & reg_re & !reg_error;
  assign extht_fail_counts_re = addr_hit[43] & reg_re & !reg_error;
  assign fw_ov_control_we = addr_hit[44] & reg_we & !reg_error;

  assign fw_ov_control_fw_ov_mode_wd = reg_wdata[3:0];

  assign fw_ov_control_fw_ov_entropy_insert_wd = reg_wdata[7:4];
  assign fw_ov_sha3_start_we = addr_hit[45] & reg_we & !reg_error;

  assign fw_ov_sha3_start_wd = reg_wdata[3:0];
  assign fw_ov_wr_fifo_full_re = addr_hit[46] & reg_re & !reg_error;
  assign fw_ov_rd_fifo_overflow_we = addr_hit[47] & reg_we & !reg_error;

  assign fw_ov_rd_fifo_overflow_wd = reg_wdata[0];
  assign fw_ov_rd_data_re = addr_hit[48] & reg_re & !reg_error;
  assign fw_ov_wr_data_we = addr_hit[49] & reg_we & !reg_error;

  assign fw_ov_wr_data_wd = reg_wdata[31:0];
  assign observe_fifo_thresh_we = addr_hit[50] & reg_we & !reg_error;

  assign observe_fifo_thresh_wd = reg_wdata[6:0];
  assign observe_fifo_depth_re = addr_hit[51] & reg_re & !reg_error;
  assign debug_status_re = addr_hit[52] & reg_re & !reg_error;
  assign recov_alert_sts_we = addr_hit[53] & reg_we & !reg_error;

  assign recov_alert_sts_fips_enable_field_alert_wd = reg_wdata[0];

  assign recov_alert_sts_entropy_data_reg_en_field_alert_wd = reg_wdata[1];

  assign recov_alert_sts_module_enable_field_alert_wd = reg_wdata[2];

  assign recov_alert_sts_threshold_scope_field_alert_wd = reg_wdata[3];

  assign recov_alert_sts_rng_bit_enable_field_alert_wd = reg_wdata[5];

  assign recov_alert_sts_fw_ov_sha3_start_field_alert_wd = reg_wdata[7];

  assign recov_alert_sts_fw_ov_mode_field_alert_wd = reg_wdata[8];

  assign recov_alert_sts_fw_ov_entropy_insert_field_alert_wd = reg_wdata[9];

  assign recov_alert_sts_es_route_field_alert_wd = reg_wdata[10];

  assign recov_alert_sts_es_type_field_alert_wd = reg_wdata[11];

  assign recov_alert_sts_es_main_sm_alert_wd = reg_wdata[12];

  assign recov_alert_sts_es_bus_cmp_alert_wd = reg_wdata[13];

  assign recov_alert_sts_es_thresh_cfg_alert_wd = reg_wdata[14];

  assign recov_alert_sts_es_fw_ov_wr_alert_wd = reg_wdata[15];

  assign recov_alert_sts_es_fw_ov_disable_alert_wd = reg_wdata[16];
  assign err_code_test_we = addr_hit[55] & reg_we & !reg_error;

  assign err_code_test_wd = reg_wdata[4:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = me_regwen_we;
    reg_we_check[5] = sw_regupd_we;
    reg_we_check[6] = 1'b0;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = module_enable_gated_we;
    reg_we_check[9] = conf_gated_we;
    reg_we_check[10] = entropy_control_gated_we;
    reg_we_check[11] = 1'b0;
    reg_we_check[12] = health_test_windows_gated_we;
    reg_we_check[13] = repcnt_thresholds_gated_we;
    reg_we_check[14] = repcnts_thresholds_gated_we;
    reg_we_check[15] = adaptp_hi_thresholds_gated_we;
    reg_we_check[16] = adaptp_lo_thresholds_gated_we;
    reg_we_check[17] = bucket_thresholds_gated_we;
    reg_we_check[18] = markov_hi_thresholds_gated_we;
    reg_we_check[19] = markov_lo_thresholds_gated_we;
    reg_we_check[20] = extht_hi_thresholds_gated_we;
    reg_we_check[21] = extht_lo_thresholds_gated_we;
    reg_we_check[22] = 1'b0;
    reg_we_check[23] = 1'b0;
    reg_we_check[24] = 1'b0;
    reg_we_check[25] = 1'b0;
    reg_we_check[26] = 1'b0;
    reg_we_check[27] = 1'b0;
    reg_we_check[28] = 1'b0;
    reg_we_check[29] = 1'b0;
    reg_we_check[30] = 1'b0;
    reg_we_check[31] = 1'b0;
    reg_we_check[32] = 1'b0;
    reg_we_check[33] = 1'b0;
    reg_we_check[34] = 1'b0;
    reg_we_check[35] = 1'b0;
    reg_we_check[36] = 1'b0;
    reg_we_check[37] = 1'b0;
    reg_we_check[38] = 1'b0;
    reg_we_check[39] = 1'b0;
    reg_we_check[40] = alert_threshold_gated_we;
    reg_we_check[41] = 1'b0;
    reg_we_check[42] = 1'b0;
    reg_we_check[43] = 1'b0;
    reg_we_check[44] = fw_ov_control_gated_we;
    reg_we_check[45] = fw_ov_sha3_start_we;
    reg_we_check[46] = 1'b0;
    reg_we_check[47] = fw_ov_rd_fifo_overflow_we;
    reg_we_check[48] = 1'b0;
    reg_we_check[49] = fw_ov_wr_data_we;
    reg_we_check[50] = observe_fifo_thresh_gated_we;
    reg_we_check[51] = 1'b0;
    reg_we_check[52] = 1'b0;
    reg_we_check[53] = recov_alert_sts_we;
    reg_we_check[54] = 1'b0;
    reg_we_check[55] = err_code_test_we;
    reg_we_check[56] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_es_entropy_valid_qs;
        reg_rdata_next[1] = intr_state_es_health_test_failed_qs;
        reg_rdata_next[2] = intr_state_es_observe_fifo_ready_qs;
        reg_rdata_next[3] = intr_state_es_fatal_err_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_es_entropy_valid_qs;
        reg_rdata_next[1] = intr_enable_es_health_test_failed_qs;
        reg_rdata_next[2] = intr_enable_es_observe_fifo_ready_qs;
        reg_rdata_next[3] = intr_enable_es_fatal_err_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
        reg_rdata_next[2] = '0;
        reg_rdata_next[3] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[0] = me_regwen_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[0] = sw_regupd_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[0] = regwen_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[7:0] = rev_abi_revision_qs;
        reg_rdata_next[15:8] = rev_hw_revision_qs;
        reg_rdata_next[23:16] = rev_chip_type_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[3:0] = module_enable_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[3:0] = conf_fips_enable_qs;
        reg_rdata_next[7:4] = conf_entropy_data_reg_enable_qs;
        reg_rdata_next[15:12] = conf_threshold_scope_qs;
        reg_rdata_next[23:20] = conf_rng_bit_enable_qs;
        reg_rdata_next[25:24] = conf_rng_bit_sel_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[3:0] = entropy_control_es_route_qs;
        reg_rdata_next[7:4] = entropy_control_es_type_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = entropy_data_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[15:0] = health_test_windows_fips_window_qs;
        reg_rdata_next[31:16] = health_test_windows_bypass_window_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[15:0] = repcnt_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = repcnt_thresholds_bypass_thresh_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[15:0] = repcnts_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = repcnts_thresholds_bypass_thresh_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[15:0] = adaptp_hi_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = adaptp_hi_thresholds_bypass_thresh_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[15:0] = adaptp_lo_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = adaptp_lo_thresholds_bypass_thresh_qs;
      end

      addr_hit[17]: begin
        reg_rdata_next[15:0] = bucket_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = bucket_thresholds_bypass_thresh_qs;
      end

      addr_hit[18]: begin
        reg_rdata_next[15:0] = markov_hi_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = markov_hi_thresholds_bypass_thresh_qs;
      end

      addr_hit[19]: begin
        reg_rdata_next[15:0] = markov_lo_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = markov_lo_thresholds_bypass_thresh_qs;
      end

      addr_hit[20]: begin
        reg_rdata_next[15:0] = extht_hi_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = extht_hi_thresholds_bypass_thresh_qs;
      end

      addr_hit[21]: begin
        reg_rdata_next[15:0] = extht_lo_thresholds_fips_thresh_qs;
        reg_rdata_next[31:16] = extht_lo_thresholds_bypass_thresh_qs;
      end

      addr_hit[22]: begin
        reg_rdata_next[15:0] = repcnt_hi_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = repcnt_hi_watermarks_bypass_watermark_qs;
      end

      addr_hit[23]: begin
        reg_rdata_next[15:0] = repcnts_hi_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = repcnts_hi_watermarks_bypass_watermark_qs;
      end

      addr_hit[24]: begin
        reg_rdata_next[15:0] = adaptp_hi_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = adaptp_hi_watermarks_bypass_watermark_qs;
      end

      addr_hit[25]: begin
        reg_rdata_next[15:0] = adaptp_lo_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = adaptp_lo_watermarks_bypass_watermark_qs;
      end

      addr_hit[26]: begin
        reg_rdata_next[15:0] = extht_hi_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = extht_hi_watermarks_bypass_watermark_qs;
      end

      addr_hit[27]: begin
        reg_rdata_next[15:0] = extht_lo_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = extht_lo_watermarks_bypass_watermark_qs;
      end

      addr_hit[28]: begin
        reg_rdata_next[15:0] = bucket_hi_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = bucket_hi_watermarks_bypass_watermark_qs;
      end

      addr_hit[29]: begin
        reg_rdata_next[15:0] = markov_hi_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = markov_hi_watermarks_bypass_watermark_qs;
      end

      addr_hit[30]: begin
        reg_rdata_next[15:0] = markov_lo_watermarks_fips_watermark_qs;
        reg_rdata_next[31:16] = markov_lo_watermarks_bypass_watermark_qs;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = repcnt_total_fails_qs;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = repcnts_total_fails_qs;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = adaptp_hi_total_fails_qs;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = adaptp_lo_total_fails_qs;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = bucket_total_fails_qs;
      end

      addr_hit[36]: begin
        reg_rdata_next[31:0] = markov_hi_total_fails_qs;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = markov_lo_total_fails_qs;
      end

      addr_hit[38]: begin
        reg_rdata_next[31:0] = extht_hi_total_fails_qs;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = extht_lo_total_fails_qs;
      end

      addr_hit[40]: begin
        reg_rdata_next[15:0] = alert_threshold_alert_threshold_qs;
        reg_rdata_next[31:16] = alert_threshold_alert_threshold_inv_qs;
      end

      addr_hit[41]: begin
        reg_rdata_next[15:0] = alert_summary_fail_counts_qs;
      end

      addr_hit[42]: begin
        reg_rdata_next[7:4] = alert_fail_counts_repcnt_fail_count_qs;
        reg_rdata_next[11:8] = alert_fail_counts_adaptp_hi_fail_count_qs;
        reg_rdata_next[15:12] = alert_fail_counts_adaptp_lo_fail_count_qs;
        reg_rdata_next[19:16] = alert_fail_counts_bucket_fail_count_qs;
        reg_rdata_next[23:20] = alert_fail_counts_markov_hi_fail_count_qs;
        reg_rdata_next[27:24] = alert_fail_counts_markov_lo_fail_count_qs;
        reg_rdata_next[31:28] = alert_fail_counts_repcnts_fail_count_qs;
      end

      addr_hit[43]: begin
        reg_rdata_next[3:0] = extht_fail_counts_extht_hi_fail_count_qs;
        reg_rdata_next[7:4] = extht_fail_counts_extht_lo_fail_count_qs;
      end

      addr_hit[44]: begin
        reg_rdata_next[3:0] = fw_ov_control_fw_ov_mode_qs;
        reg_rdata_next[7:4] = fw_ov_control_fw_ov_entropy_insert_qs;
      end

      addr_hit[45]: begin
        reg_rdata_next[3:0] = fw_ov_sha3_start_qs;
      end

      addr_hit[46]: begin
        reg_rdata_next[0] = fw_ov_wr_fifo_full_qs;
      end

      addr_hit[47]: begin
        reg_rdata_next[0] = fw_ov_rd_fifo_overflow_qs;
      end

      addr_hit[48]: begin
        reg_rdata_next[31:0] = fw_ov_rd_data_qs;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[50]: begin
        reg_rdata_next[6:0] = observe_fifo_thresh_qs;
      end

      addr_hit[51]: begin
        reg_rdata_next[6:0] = observe_fifo_depth_qs;
      end

      addr_hit[52]: begin
        reg_rdata_next[2:0] = debug_status_entropy_fifo_depth_qs;
        reg_rdata_next[5:3] = debug_status_sha3_fsm_qs;
        reg_rdata_next[6] = debug_status_sha3_block_pr_qs;
        reg_rdata_next[7] = debug_status_sha3_squeezing_qs;
        reg_rdata_next[8] = debug_status_sha3_absorbed_qs;
        reg_rdata_next[9] = debug_status_sha3_err_qs;
        reg_rdata_next[16] = debug_status_main_sm_idle_qs;
        reg_rdata_next[17] = debug_status_main_sm_boot_done_qs;
      end

      addr_hit[53]: begin
        reg_rdata_next[0] = recov_alert_sts_fips_enable_field_alert_qs;
        reg_rdata_next[1] = recov_alert_sts_entropy_data_reg_en_field_alert_qs;
        reg_rdata_next[2] = recov_alert_sts_module_enable_field_alert_qs;
        reg_rdata_next[3] = recov_alert_sts_threshold_scope_field_alert_qs;
        reg_rdata_next[5] = recov_alert_sts_rng_bit_enable_field_alert_qs;
        reg_rdata_next[7] = recov_alert_sts_fw_ov_sha3_start_field_alert_qs;
        reg_rdata_next[8] = recov_alert_sts_fw_ov_mode_field_alert_qs;
        reg_rdata_next[9] = recov_alert_sts_fw_ov_entropy_insert_field_alert_qs;
        reg_rdata_next[10] = recov_alert_sts_es_route_field_alert_qs;
        reg_rdata_next[11] = recov_alert_sts_es_type_field_alert_qs;
        reg_rdata_next[12] = recov_alert_sts_es_main_sm_alert_qs;
        reg_rdata_next[13] = recov_alert_sts_es_bus_cmp_alert_qs;
        reg_rdata_next[14] = recov_alert_sts_es_thresh_cfg_alert_qs;
        reg_rdata_next[15] = recov_alert_sts_es_fw_ov_wr_alert_qs;
        reg_rdata_next[16] = recov_alert_sts_es_fw_ov_disable_alert_qs;
      end

      addr_hit[54]: begin
        reg_rdata_next[0] = err_code_sfifo_esrng_err_qs;
        reg_rdata_next[1] = err_code_sfifo_observe_err_qs;
        reg_rdata_next[2] = err_code_sfifo_esfinal_err_qs;
        reg_rdata_next[20] = err_code_es_ack_sm_err_qs;
        reg_rdata_next[21] = err_code_es_main_sm_err_qs;
        reg_rdata_next[22] = err_code_es_cntr_err_qs;
        reg_rdata_next[23] = err_code_sha3_state_err_qs;
        reg_rdata_next[24] = err_code_sha3_rst_storage_err_qs;
        reg_rdata_next[28] = err_code_fifo_write_err_qs;
        reg_rdata_next[29] = err_code_fifo_read_err_qs;
        reg_rdata_next[30] = err_code_fifo_state_err_qs;
      end

      addr_hit[55]: begin
        reg_rdata_next[4:0] = err_code_test_qs;
      end

      addr_hit[56]: begin
        reg_rdata_next[8:0] = main_sm_state_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src high or how watermark register module
//

module entropy_src_watermark_reg #(
  parameter int RegWidth = 16,
  parameter bit HighWatermark = 1
) (
  input logic                   clk_i,
  input logic                   rst_ni,

   // functional interface
  input logic                   clear_i,
  input logic                   event_i,
  input logic [RegWidth-1:0]    value_i,
  output logic [RegWidth-1:0]   value_o
);

  // signals
  logic [RegWidth-1:0] event_cntr_change;
  logic [RegWidth-1:0] reg_reset;

  // flops
  logic [RegWidth-1:0] event_cntr_q, event_cntr_d;

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      event_cntr_q       <= reg_reset;
    end else begin
      event_cntr_q       <= event_cntr_d;
    end

  assign event_cntr_d = clear_i ? reg_reset :
                        event_i ? event_cntr_change :
                        event_cntr_q;

  // Set mode of this counter to be either a high or low watermark
  if (HighWatermark) begin : gen_hi_wm

    assign reg_reset = {RegWidth{1'b0}};

    assign event_cntr_change = (value_i > event_cntr_q) ? (value_i) : event_cntr_q;

  end else begin : gen_lo_wm

    assign reg_reset = {RegWidth{1'b1}};

    assign event_cntr_change = (value_i < event_cntr_q) ? (value_i) : event_cntr_q;

  end

  // drive output
  assign value_o = event_cntr_q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Supports writing a field that enables
// a function within a module.
// Requirements are that the function will
// only be enabled when the field is written
// the it is the inverse of the current field
// setting. The can only toggle between the
// the on value and the off value.


module entropy_src_field_en #(
  parameter int FieldW  = 4,
  parameter int FieldEnVal = 'ha
) (
  input logic clk_i ,
  input logic rst_ni,
  input logic               wvalid_i,
  input logic [FieldW-1:0]  wdata_i,

  output logic              enable_o
);

  // signal
  logic  field_update;
  logic [FieldW-1:0] field_value;
  logic [FieldW-1:0] field_value_invert;

  // flops
  logic [FieldW-1:0] field_q, field_d;

  assign  field_value = FieldEnVal;
  assign  field_value_invert = ~field_value;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      field_q <= field_value_invert;
    end else begin
      field_q <= field_d;
    end
  end

  assign field_update = wvalid_i && (field_q == ~wdata_i) &&
                        ((wdata_i == field_value) ||
                         (wdata_i == field_value_invert));

  assign field_d = field_update ? wdata_i : field_q;

  assign enable_o = (field_q == field_value);


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src counter register module
//

module entropy_src_cntr_reg #(
  parameter int RegWidth = 16
) (
  input logic                   clk_i,
  input logic                   rst_ni,

   // functional interface
  input logic                   clear_i,
  input logic                   event_i,
  output logic [RegWidth-1:0]   value_o,
  output logic                  err_o
);

  // signals
  logic [RegWidth-1:0] counter_value;

  // counter will not wrap when full value is reached
  prim_count #(
    .Width(RegWidth)
  ) u_prim_count_cntr_reg (
    .clk_i,
    .rst_ni,
    .clr_i(clear_i),
    .set_i(1'b0),
    .set_cnt_i(RegWidth'(0)),
    .incr_en_i(event_i && (~counter_value != '0)),
    .decr_en_i(1'b0),
    .step_i(RegWidth'(1)),
    .cnt_o(counter_value),
    .cnt_next_o(),
    .err_o(err_o)
  );

  assign value_o = counter_value;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: interface between a req/ack interface and a fifo
//

module entropy_src_ack_sm (
  input logic                clk_i,
  input logic                rst_ni,

  input logic                enable_i,
  input logic                req_i,
  output logic               ack_o,
  input logic                fifo_not_empty_i,
  input logic                local_escalate_i,
  output logic               fifo_pop_o,
  output logic               ack_sm_err_o
);

  import entropy_src_ack_sm_pkg::*;

  state_e state_d, state_q;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, Idle)

  always_comb begin
    state_d = state_q;
    ack_o = 1'b0;
    fifo_pop_o = 1'b0;
    ack_sm_err_o = 1'b0;
    unique case (state_q)
      Idle: begin
        if (enable_i) begin
          if (req_i) begin
            state_d = Wait;
          end
        end
      end
      Wait: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          if (fifo_not_empty_i) begin
            ack_o = 1'b1;
            fifo_pop_o = 1'b1;
            state_d = Idle;
          end
        end
      end
      Error: begin
        ack_sm_err_o = 1'b1;
      end
      default: begin
        state_d = Error;
        ack_sm_err_o = 1'b1;
      end
    endcase
    if (local_escalate_i) begin
      state_d = Error;
    end
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src main state machine module
//
//   determines when new entropy is ready to be forwarded

module entropy_src_main_sm
  import entropy_src_main_sm_pkg::*;
(
  input logic                   clk_i,
  input logic                   rst_ni,

  input logic                   enable_i,
  input logic                   fw_ov_ent_insert_i,
  input logic                   fw_ov_sha3_start_i,
  input logic                   ht_done_pulse_i,
  input logic                   ht_fail_pulse_i,
  input logic                   alert_thresh_fail_i,
  output logic                  rst_alert_cntr_o,
  input logic                   bypass_mode_i,
  input logic                   main_stage_rdy_i,
  input logic                   bypass_stage_rdy_i,
  input logic                   sha3_state_vld_i,
  output logic                  main_stage_push_o,
  output logic                  bypass_stage_pop_o,
  output logic                  boot_phase_done_o,
  output logic                  sha3_start_o,
  output logic                  sha3_process_o,
  output prim_mubi_pkg::mubi4_t sha3_done_o,
  output logic                  cs_aes_halt_req_o,
  input logic                   cs_aes_halt_ack_i,
  input logic                   local_escalate_i,
  output logic                  main_sm_alert_o,
  output logic                  main_sm_idle_o,
  output logic [StateWidth-1:0] main_sm_state_o,
  output logic                  main_sm_err_o
);

  // The definition of state_e, the sparse FSM state enum, is in entropy_src_main_sm_pkg.sv
  state_e state_d, state_q;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, Idle)

  assign main_sm_state_o = state_q;

  always_comb begin
    state_d = state_q;
    rst_alert_cntr_o = 1'b0;
    main_stage_push_o = 1'b0;
    bypass_stage_pop_o = 1'b0;
    boot_phase_done_o = 1'b0;
    sha3_start_o = 1'b0;
    sha3_process_o = 1'b0;
    sha3_done_o = prim_mubi_pkg::MuBi4False;
    cs_aes_halt_req_o = 1'b0;
    main_sm_alert_o = 1'b0;
    main_sm_idle_o = 1'b0;
    main_sm_err_o = 1'b0;
    unique case (state_q)
      Idle: begin
        main_sm_idle_o = 1'b1;
        if (enable_i) begin
          // running fw override mode and in sha3 mode
          if (fw_ov_ent_insert_i && !bypass_mode_i) begin
            sha3_start_o = 1'b1;
            if (fw_ov_sha3_start_i) begin
              state_d = FWInsertMsg;
            end else begin
              state_d = FWInsertStart;
            end
          // running in bypass_mode and not fw override mode
          end else if (bypass_mode_i && !fw_ov_ent_insert_i) begin
            state_d = BootHTRunning;
          // running in bypass_mode and fw override mode
          end else if (bypass_mode_i && fw_ov_ent_insert_i) begin
            state_d = Idle;
          end else begin
            state_d = StartupHTStart;
          end
        end
      end
      BootHTRunning: begin
        if (!enable_i) begin
          state_d = Idle;
        end else if (ht_done_pulse_i) begin
          if (ht_fail_pulse_i) begin
            if (bypass_stage_rdy_i) begin
              // Remove failed data
              bypass_stage_pop_o = 1'b1;
            end
            if (alert_thresh_fail_i) begin
              state_d = AlertState;
            end else begin
              state_d = Idle;
            end
          end else begin
            // Window sizes other than 384 bits (the seed length) are currently not tested nor
            // supported in bypass or boot-time mode.
            state_d = BootPostHTChk;
            rst_alert_cntr_o = 1'b1;
          end
        end
      end
      BootPostHTChk: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          if (!bypass_stage_rdy_i) begin
          end else begin
            bypass_stage_pop_o = 1'b1;
            main_stage_push_o = 1'b1;
            state_d = BootPhaseDone;
          end
        end
      end
      BootPhaseDone: begin
        boot_phase_done_o = 1'b1;
        if (!enable_i) begin
          state_d = Idle;
        end
        // Even when stalled we keep monitoring for alerts and maintaining  alert statistics.
        // However, we don't signal alerts or clear HT stats in FW_OV mode.
        if(!fw_ov_ent_insert_i && ht_done_pulse_i) begin
          if (alert_thresh_fail_i) begin
            state_d = AlertState;
          end else if (!ht_fail_pulse_i) begin
            rst_alert_cntr_o = 1'b1;
          end
        end
      end
      StartupHTStart: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          sha3_start_o = 1'b1;
          state_d = StartupPhase1;
        end
      end
      StartupPhase1: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          if (ht_done_pulse_i) begin
            if (ht_fail_pulse_i) begin
              state_d = StartupFail1;
            end else begin
              state_d = StartupPass1;
              rst_alert_cntr_o = 1'b1;
            end
          end
        end
      end
      StartupPass1: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          if (ht_done_pulse_i) begin
            if (ht_fail_pulse_i) begin
              state_d = StartupFail1;
            end else begin
              // Passed two consecutive tests
              state_d = Sha3Prep;
              rst_alert_cntr_o = 1'b1;
            end
          end
        end
      end
      StartupFail1: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          if (ht_done_pulse_i) begin
            if (ht_fail_pulse_i) begin
              // Failed two consecutive tests
              state_d = AlertState;
            end else begin
              state_d = StartupPass1;
              rst_alert_cntr_o = 1'b1;
            end
          end
        end
      end
      ContHTStart: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          sha3_start_o = 1'b1;
          state_d = ContHTRunning;
        end
      end
      ContHTRunning: begin
        if (!enable_i) begin
          state_d = Idle;
        end else begin
          if (ht_done_pulse_i) begin
            if (alert_thresh_fail_i) begin
              state_d = AlertState;
            end else if (!ht_fail_pulse_i) begin
              state_d = Sha3Prep;
              rst_alert_cntr_o = 1'b1;
            end
          end
        end
      end
      FWInsertStart: begin
        if (!enable_i) begin
          state_d = Idle;
        end else if (fw_ov_sha3_start_i) begin
          state_d = FWInsertMsg;
        end
      end
      FWInsertMsg: begin
        if (!enable_i) begin
          state_d = Idle;
        end else if (!fw_ov_sha3_start_i) begin
          state_d = Sha3Prep;
        end
      end
      Sha3Prep: begin
        // for normal or halt cases, always prevent a power spike
        cs_aes_halt_req_o = 1'b1;
        if (cs_aes_halt_ack_i) begin
          state_d = Sha3Process;
        end
      end
      Sha3Process: begin
        cs_aes_halt_req_o = 1'b1;
        sha3_process_o = 1'b1;
        state_d = Sha3Valid;
      end
      Sha3Valid: begin
        cs_aes_halt_req_o = 1'b1;
        if (sha3_state_vld_i) begin
          state_d = Sha3Done;
        end
      end
      Sha3Done: begin
        if (!enable_i) begin
          sha3_done_o = prim_mubi_pkg::MuBi4True;
          state_d = Sha3MsgDone;
        end else begin
          if (main_stage_rdy_i) begin
            sha3_done_o = prim_mubi_pkg::MuBi4True;
            main_stage_push_o = 1'b1;
            state_d = Sha3MsgDone;
          end
        end
      end
      Sha3MsgDone: begin
        if (!cs_aes_halt_ack_i) begin
          state_d = Sha3Quiesce;
        end
      end
      Sha3Quiesce: begin
        if (!enable_i || fw_ov_ent_insert_i) begin
          state_d = Idle;
        end else begin
          state_d = ContHTStart;
        end
      end
      AlertState: begin
        main_sm_alert_o = 1'b1;
        state_d = AlertHang;
      end
      AlertHang: begin
        if (!enable_i) begin
          state_d = Idle;
        end
      end
      Error: begin
        main_sm_err_o = 1'b1;
      end
      default: begin
        state_d = Error;
        main_sm_err_o = 1'b1;
      end
    endcase
    if (local_escalate_i) begin
      state_d = Error;
    end
  end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src repetitive count health test module
//

module entropy_src_repcnt_ht #(
  parameter int RegWidth = 16,
  parameter int RngBusWidth = 4
) (
  input logic                   clk_i,
  input logic                   rst_ni,

   // ins req interface
  input logic [RngBusWidth-1:0] entropy_bit_i,
  input logic                   entropy_bit_vld_i,
  input logic                   clear_i,
  input logic                   active_i,
  input logic [RegWidth-1:0]    thresh_i,
  output logic [RegWidth-1:0]   test_cnt_o,
  output logic                  test_fail_pulse_o,
  output logic                  count_err_o
);

  // signals
  logic [RngBusWidth-1:0]               samples_match_pulse;
  logic [RngBusWidth-1:0]               samples_no_match_pulse;
  logic [RngBusWidth-1:0]               rep_cnt_fail;
  logic [RngBusWidth-1:0][RegWidth-1:0] rep_cntr;
  logic [RngBusWidth-1:0]               rep_cntr_err;
  logic [RegWidth-1:0]                  cntr_max;
  logic                                 fail_sampled;

  // flops
  logic [RngBusWidth-1:0] prev_sample_q, prev_sample_d;
  logic fail_sample_mask_d, fail_sample_mask_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      prev_sample_q       <= '0;
      fail_sample_mask_q  <= '0;
    end else begin
      prev_sample_q       <= prev_sample_d;
      fail_sample_mask_q  <= fail_sample_mask_d;
    end
  end

  // Repetitive Count Test
  //
  // Test operation
  //  This test will look for catastrophic stuck bit failures. The rep_cntr
  //  uses one as the starting value, just as the NIST algorithm does.


  for (genvar sh = 0; sh < RngBusWidth; sh = sh+1) begin : gen_cntrs


    // NIST A sample
    assign prev_sample_d[sh] = (!active_i || clear_i) ? '0 :
                               entropy_bit_vld_i ? entropy_bit_i[sh] :
                               prev_sample_q[sh];

    assign samples_match_pulse[sh] = entropy_bit_vld_i &&
           (prev_sample_q[sh] == entropy_bit_i[sh]);
    assign samples_no_match_pulse[sh] = entropy_bit_vld_i &&
           (prev_sample_q[sh] != entropy_bit_i[sh]);

    // NIST B counter
    // SEC_CM: CTR.REDUN
    prim_count #(
      .Width(RegWidth)
    ) u_prim_count_rep_cntr (
      .clk_i,
      .rst_ni,
      .clr_i(1'b0),
      .set_i(!active_i || clear_i || samples_no_match_pulse[sh]),
      .set_cnt_i(RegWidth'(1)),
      .incr_en_i(samples_match_pulse[sh]),
      .decr_en_i(1'b0),
      .step_i(RegWidth'(1)),
      .cnt_o(rep_cntr[sh]),
      .cnt_next_o(),
      .err_o(rep_cntr_err[sh])
    );

    assign rep_cnt_fail[sh] = (rep_cntr[sh] >= thresh_i);

  end : gen_cntrs

  prim_max_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_prim_max_tree_rep_cntr_max (
    .clk_i,
    .rst_ni,
    .values_i   (rep_cntr),
    .valid_i    ({RngBusWidth{1'b1}}),
    .max_value_o(cntr_max),
    .max_idx_o  (),
    .max_valid_o()
  );

  // For the purposes of failure pulse generation, we want to sample
  // the test output for only one cycle and do it immediately after
  // the counter has been updated.
  assign fail_sample_mask_d = entropy_bit_vld_i;
  assign fail_sampled       = |rep_cnt_fail & fail_sample_mask_q;

  assign test_fail_pulse_o = active_i & fail_sampled;

  assign test_cnt_o = cntr_max;
  assign count_err_o = (|rep_cntr_err);


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src repetitive count symbol based health test module
//

module entropy_src_repcnts_ht #(
  parameter int RegWidth = 16,
  parameter int RngBusWidth = 4
) (
  input logic clk_i,
  input logic rst_ni,

   // ins req interface
  input logic [RngBusWidth-1:0] entropy_bit_i,
  input logic                   entropy_bit_vld_i,
  input logic                   clear_i,
  input logic                   active_i,
  input logic [RegWidth-1:0]    thresh_i,
  output logic [RegWidth-1:0]   test_cnt_o,
  output logic                  test_fail_pulse_o,
  output logic                  count_err_o
);

  // signals
  logic  samples_match_pulse;
  logic  samples_no_match_pulse;
  logic  rep_cnt_fail;
  logic [RegWidth-1:0]    rep_cntr;
  logic                   rep_cntr_err;
  logic                   fail_sampled;

  // flops
  logic [RngBusWidth-1:0] prev_sample_q, prev_sample_d;
  logic fail_sample_mask_d, fail_sample_mask_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      prev_sample_q      <= '0;
      fail_sample_mask_q <= '0;
    end else begin
      prev_sample_q      <= prev_sample_d;
      fail_sample_mask_q <= fail_sample_mask_d;
    end
  end

  // Repetitive Count Test for symbols
  //
  // Test operation
  //  This test will look for catastrophic stuck bit failures. The rep_cntr
  //  uses one as the starting value, just as the NIST algorithm does.


  // NIST A sample
  assign prev_sample_d = (!active_i || clear_i) ? '0 :
                         entropy_bit_vld_i ? entropy_bit_i :
                         prev_sample_q;

  assign samples_match_pulse = entropy_bit_vld_i &&
         (prev_sample_q == entropy_bit_i);
  assign samples_no_match_pulse = entropy_bit_vld_i &&
         (prev_sample_q != entropy_bit_i);

  // NIST B counter
  // SEC_CM: CTR.REDUN
  prim_count #(
    .Width(RegWidth)
  ) u_prim_count_rep_cntr (
    .clk_i,
    .rst_ni,
    .clr_i(1'b0),
    .set_i(!active_i || clear_i || samples_no_match_pulse),
    .set_cnt_i(RegWidth'(1)),
    .incr_en_i(samples_match_pulse),
    .decr_en_i(1'b0),
    .step_i(RegWidth'(1)),
    .cnt_o(rep_cntr),
    .cnt_next_o(),
    .err_o(rep_cntr_err)
  );

  assign rep_cnt_fail = (rep_cntr >= thresh_i);

  // For the purposes of failure pulse generation, we want to sample
  // the test output for only one cycle and do it immediately after
  // the counter has been updated.
  assign fail_sample_mask_d = entropy_bit_vld_i;
  assign fail_sampled       = rep_cnt_fail & fail_sample_mask_q;

  assign test_fail_pulse_o = active_i & fail_sampled;

  assign test_cnt_o = rep_cntr;
  assign count_err_o = (|rep_cntr_err);


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src adaptive proportion health test module
//

module entropy_src_adaptp_ht #(
  parameter int RegWidth = 16,
  parameter int RngBusWidth = 4
) (
  input logic clk_i,
  input logic rst_ni,

   // ins req interface
  input logic [RngBusWidth-1:0] entropy_bit_i,
  input logic                   entropy_bit_vld_i,
  input logic                   clear_i,
  input logic                   active_i,
  input logic [RegWidth-1:0]    thresh_hi_i,
  input logic [RegWidth-1:0]    thresh_lo_i,
  input logic                   window_wrap_pulse_i,
  input logic                   threshold_scope_i,
  output logic [RegWidth-1:0]   test_cnt_hi_o,
  output logic [RegWidth-1:0]   test_cnt_lo_o,
  output logic                  test_fail_hi_pulse_o,
  output logic                  test_fail_lo_pulse_o,
  output logic                  count_err_o
);

  // signals
  logic [RegWidth-1:0]                  test_cnt_max;
  logic [RegWidth-1:0]                  test_cnt_min, test_cnt_min_tmp;
  logic [RegWidth-1:0]                  test_cnt_sum;
  logic [RngBusWidth-1:0][RegWidth-1:0] test_cnt;
  logic [RngBusWidth-1:0]               test_cnt_err;

  // Adaptive Proportion Test
  //
  // Test operation
  //  This is an approved modification of the NIST Adaptive Proportion test in that
  //  instead of counting the first sampled value (1'b1 or 1'b0), it will count
  //  only the 1's on all four bit streams and accumulate for the during of the
  //  window size (W) of the test.

  for (genvar sh = 0; sh < RngBusWidth; sh = sh+1) begin : gen_cntrs

    // cumulative ones counter
    // SEC_CM: CTR.REDUN
    prim_count #(
      .Width(RegWidth)
    ) u_prim_count_test_cnt (
      .clk_i,
      .rst_ni,
      .clr_i(window_wrap_pulse_i),
      .set_i(!active_i || clear_i),
      .set_cnt_i(RegWidth'(0)),
      .incr_en_i(entropy_bit_vld_i),
      .decr_en_i(1'b0),
      .step_i(RegWidth'(entropy_bit_i[sh])),
      .cnt_o(test_cnt[sh]),
      .cnt_next_o(),
      .err_o(test_cnt_err[sh])
    );
  end : gen_cntrs

  // determine the highest counter counter value
  prim_max_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_max (
    .clk_i       (clk_i),
    .rst_ni      (rst_ni),
    .values_i    (test_cnt),
    .valid_i     ({RngBusWidth{1'b1}}),
    .max_value_o (test_cnt_max),
    .max_idx_o   (),
    .max_valid_o ()
  );

  // determine the lowest counter value
  // Negate the inputs and outputs of prim_max_tree to find the minimum
  // For this unsigned application, one's complement negation (i.e. logical inversion) is fine.
  prim_max_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_min (
    .clk_i       (clk_i),
    .rst_ni      (rst_ni),
    .values_i    (~test_cnt),
    .valid_i     ({RngBusWidth{1'b1}}),
    .max_value_o (test_cnt_min_tmp),
    .max_idx_o   (),
    .max_valid_o ()
  );

  assign test_cnt_min = ~test_cnt_min_tmp;

  prim_sum_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_sum (
    .clk_i       (clk_i),
    .rst_ni      (rst_ni),
    .values_i    (test_cnt),
    .valid_i     ({RngBusWidth{1'b1}}),
    .sum_value_o (test_cnt_sum),
    .sum_valid_o ()
  );

  assign test_cnt_hi_o = threshold_scope_i ? test_cnt_sum : test_cnt_max;
  assign test_cnt_lo_o = threshold_scope_i ? test_cnt_sum : test_cnt_min;

  // the pulses will be only one clock in length
  assign test_fail_hi_pulse_o = active_i && window_wrap_pulse_i && (test_cnt_hi_o > thresh_hi_i);
  assign test_fail_lo_pulse_o = active_i && window_wrap_pulse_i && (test_cnt_lo_o < thresh_lo_i);
  assign count_err_o = |test_cnt_err;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src bucket health test module
//

module entropy_src_bucket_ht #(
  parameter int RegWidth = 16,
  parameter int RngBusWidth = 4
) (
  input logic clk_i,
  input logic rst_ni,

   // ins req interface
  input logic [RngBusWidth-1:0] entropy_bit_i,
  input logic                   entropy_bit_vld_i,
  input logic                   clear_i,
  input logic                   active_i,
  input logic [RegWidth-1:0]    thresh_i,
  input logic                   window_wrap_pulse_i,
  output logic [RegWidth-1:0]   test_cnt_o,
  output logic                  test_fail_pulse_o,
  output logic                  count_err_o
);

  localparam int NUM_BINS = 2**RngBusWidth;

  // signals
  logic [NUM_BINS-1:0] bin_incr;
  logic [NUM_BINS-1:0] bin_cnt_exceeds_thresh;
  logic [NUM_BINS - 1:0][RegWidth - 1:0] bin_cntr;
  logic [NUM_BINS-1:0] bin_cntr_err;
  logic [RegWidth-1:0] bin_max;

  // Bucket Test
  //
  // Test operation
  //  This test will look at 4 bit symbols and increment one of sixteen
  //  counters, or buckets, to show a histogram of the data stream.
  //  An error will occur if one of the counters reaches the thresh
  //  value.


  // Analyze the incoming symbols

  for (genvar i = 0; i < NUM_BINS; i = i + 1) begin : gen_symbol_match
    // set the bin incrementer if the symbol matches that bin
    assign bin_incr[i] = entropy_bit_vld_i && (entropy_bit_i == i);
    // use the bin incrementer to increase the bin total count
    // SEC_CM: CTR.REDUN
    prim_count #(
      .Width(RegWidth)
    ) u_prim_count_bin_cntr (
      .clk_i,
      .rst_ni,
      .clr_i(window_wrap_pulse_i),
      .set_i(!active_i || clear_i),
      .set_cnt_i(RegWidth'(0)),
      .incr_en_i(bin_incr[i]),
      .decr_en_i(1'b0),
      .step_i(RegWidth'(1)),
      .cnt_o(bin_cntr[i]),
      .cnt_next_o(),
      .err_o(bin_cntr_err[i])
    );
    assign bin_cnt_exceeds_thresh[i] = (bin_cntr[i] > thresh_i);
  end : gen_symbol_match

  prim_max_tree #(
    .NumSrc(NUM_BINS),
    .Width(RegWidth)
  ) u_prim_max_tree_bin_cntr_max (
    .clk_i,
    .rst_ni,
    .values_i   (bin_cntr),
    .valid_i    ({RegWidth{1'b1}}),
    .max_value_o(bin_max),
    .max_idx_o  (),
    .max_valid_o()
  );

  // the pulses will be only one clock in length
  assign test_fail_pulse_o = active_i && window_wrap_pulse_i && (|bin_cnt_exceeds_thresh);
  assign test_cnt_o = bin_max;
  assign count_err_o = |bin_cntr_err;


endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src Markov health test module
//

module entropy_src_markov_ht #(
  parameter int RegWidth = 16,
  parameter int RngBusWidth = 4
) (
  input logic clk_i,
  input logic rst_ni,

   // ins req interface
  input logic [RngBusWidth-1:0] entropy_bit_i,
  input logic                   entropy_bit_vld_i,
  input logic                   clear_i,
  input logic                   active_i,
  input logic [RegWidth-1:0]    thresh_hi_i,
  input logic [RegWidth-1:0]    thresh_lo_i,
  input logic                   window_wrap_pulse_i,
  input logic                   threshold_scope_i,
  output logic [RegWidth-1:0]   test_cnt_hi_o,
  output logic [RegWidth-1:0]   test_cnt_lo_o,
  output logic                  test_fail_hi_pulse_o,
  output logic                  test_fail_lo_pulse_o,
  output logic                  count_err_o
);

  // signals
  logic [RngBusWidth-1:0] samples_no_match_pulse;
  logic [RegWidth-1:0]                  pair_cntr_max;
  logic [RegWidth-1:0]                  pair_cntr_min, pair_cntr_min_tmp;
  logic [RegWidth-1:0]                  pair_cntr_sum;
  logic [RngBusWidth-1:0][RegWidth-1:0] pair_cntr;
  logic [RngBusWidth-1:0]               pair_cntr_err;

  // flops
  logic                toggle_q, toggle_d;
  logic [RngBusWidth-1:0] prev_sample_q, prev_sample_d;

  always_ff @(posedge clk_i or negedge rst_ni)
    if (!rst_ni) begin
      toggle_q         <= '0;
      prev_sample_q    <= '0;
    end else begin
      toggle_q         <= toggle_d;
      prev_sample_q    <= prev_sample_d;
    end


  // Markov Test
  //
  // Test operation
  //  This test will look at pairs of bit levels per bitstream. A counter for
  //  stream will only count when the pair equals 0b01 or 0b10.


  for (genvar sh = 0; sh < RngBusWidth; sh = sh+1) begin : gen_cntrs

    // bit sampler
    assign prev_sample_d[sh] = (!active_i || clear_i) ? '0 :
                               window_wrap_pulse_i ? '0  :
                               entropy_bit_vld_i ? entropy_bit_i[sh] :
                               prev_sample_q[sh];

    // pair check
    assign samples_no_match_pulse[sh] = entropy_bit_vld_i && toggle_q &&
           (prev_sample_q[sh] == !entropy_bit_i[sh]);

    // pair counter
    prim_count #(
      .Width(RegWidth)
    ) u_prim_count_pair_cntr (
      .clk_i,
      .rst_ni,
      .clr_i(window_wrap_pulse_i),
      .set_i(!active_i || clear_i),
      .set_cnt_i(RegWidth'(0)),
      .incr_en_i(samples_no_match_pulse[sh]),
      .decr_en_i(1'b0),
      .step_i(RegWidth'(1)),
      .cnt_o(pair_cntr[sh]),
      .cnt_next_o(),
      .err_o(pair_cntr_err[sh])
    );
  end : gen_cntrs

  // create a toggle signal to sample pairs with
  assign toggle_d = (!active_i || clear_i) ? '0 :
                    window_wrap_pulse_i ? '0  :
                    entropy_bit_vld_i ? (!toggle_q) :
                    toggle_q;

  // determine the highest counter pair counter value
  prim_max_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_max (
    .clk_i       (clk_i),
    .rst_ni      (rst_ni),
    .values_i    (pair_cntr),
    .valid_i     ({RngBusWidth{1'b1}}),
    .max_value_o (pair_cntr_max),
    .max_idx_o   (),
    .max_valid_o ()
  );

  // determine the lowest counter pair counter value
  // Negate the inputs and outputs of prim_max_tree to find the minimum
  // For this unsigned application, one's complement negation (i.e. logical inversion) is fine.
  prim_max_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_min (
    .clk_i       (clk_i),
    .rst_ni      (rst_ni),
    .values_i    (~pair_cntr),
    .valid_i     ({RngBusWidth{1'b1}}),
    .max_value_o (pair_cntr_min_tmp),
    .max_idx_o   (),
    .max_valid_o ()
  );

  // Invert the output back.
  assign pair_cntr_min = ~pair_cntr_min_tmp;

  prim_sum_tree #(
    .NumSrc(RngBusWidth),
    .Width(RegWidth)
  ) u_sum (
    .clk_i       (clk_i),
    .rst_ni      (rst_ni),
    .values_i    (pair_cntr),
    .valid_i     ({RngBusWidth{1'b1}}),
    .sum_value_o (pair_cntr_sum),
    .sum_valid_o ()
  );

  assign test_cnt_hi_o = threshold_scope_i ? pair_cntr_sum : pair_cntr_max;
  assign test_cnt_lo_o = threshold_scope_i ? pair_cntr_sum : pair_cntr_min;

  // the pulses will be only one clock in length
  assign test_fail_hi_pulse_o = active_i && window_wrap_pulse_i && (test_cnt_hi_o > thresh_hi_i);
  assign test_fail_lo_pulse_o = active_i && window_wrap_pulse_i && (test_cnt_lo_o < thresh_lo_i);
  assign count_err_o = (|pair_cntr_err);

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: Logic module indicate ongoing activity of after disablement of entropy_src_core
//
// The entropy_src has a great deal of internal state, and when shutting down most of this internal
// state should be cleared.  (The two notable exceptions are the health test statistics, which are
// only cleared at the next enable, and the SHA3 conditioning sponge which accumulates unused
// entropy until a seed is generated).  There are delays as incoming RNG data is processed, and for
// ease of verification we insist all elements of the data pipeline are cleared consistently.  This
// means that once an RNG sample enters the pipeline, that sample should be reflected in the health
// tests. The SHA3 conditioner is also assumed to successfully absorb every 64-bits that enters the
// module.
//
// To acheive this consistency goal the entropy_src delays the clearing of internal data buffers
// and the state machine until:
// 1. Any unprocessed data has been counted at the health checks (regardless of the mode)
// 2. Any RNG data bound for the SHA conditioner has been received at the conditioner.
// 3. Any ongoing SHA processing operations have completed, and the main FSM has been forced
//    back to idle.
//
// This block creates a modified version of the enable pulse which:
// 1. Postpones the disable event until any flowing data has passed through the RNG, ESBIT and
//    POSTHT FIFOs.  If packpressure is encountered at the Precon FIFO, the stalled data can
//    be discarded, and so a has a maximum time limit of MaxFifoWait=3 clocks is given for this
//    check.
// 2. Once the disable signal is received, the rising edge does not occur until:
//    2a. One clock after the falling edge OR
//    2b. One clock after the SHA engine completes,
//    Whichever comes later.

module entropy_src_enable_delay import prim_mubi_pkg::*; (
  input logic  clk_i,
  input logic  rst_ni,

  input logic  enable_i,

  // Unconsumed FIFO inputs
  input logic esrng_fifo_not_empty_i,
  input logic esbit_fifo_not_empty_i,
  input logic postht_fifo_not_empty_i,

  // SHA3 conditioner inputs
  input logic   cs_aes_halt_req_i,
  input mubi4_t sha3_done_i,

  input logic bypass_mode_i,

  output logic enable_o
);

  // Maximum number of cycles to wait for FIFOs to clear out.
  // Set to 3 to allow one cycle for each FIFO in the pipeline.
  localparam int MaxFifoWait = 3;

  logic suppress_reenable;
  logic extend_enable;

  logic data_in_flight;
  logic [2:0] fifos_not_empty;

  // Flops
  logic [MaxFifoWait - 1:0] fifo_timer_d, fifo_timer_q;
  logic                     sha3_active_post_en_d, sha3_active_post_en_q;
  mubi4_t                   sha3_done_q;
  logic                     extend_enable_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      sha3_active_post_en_q   <= 1'b0;
      fifo_timer_q            <= '0;
      sha3_done_q             <= prim_mubi_pkg::MuBi4False;
      extend_enable_q         <= 1'b0;
    end else begin
      sha3_active_post_en_q   <= sha3_active_post_en_d;
      fifo_timer_q            <= fifo_timer_d;
      sha3_done_q             <= sha3_done_i;
      extend_enable_q         <= extend_enable;
    end
  end

  // Output definition
  assign enable_o = (enable_i & ~suppress_reenable) | extend_enable;

  // In flight data monitoring.
  // The `fifo_timer` is a small shift register to count out the maximum number of cycles to wait
  // for the FIFOs to drain. Since this timer is very small (3 cycles), it is implemented as a shift
  // register.
  assign fifo_timer_d = enable_i ? {MaxFifoWait{1'b1}} : {fifo_timer_q[MaxFifoWait-2:0], 1'b0};
  assign fifos_not_empty = {esrng_fifo_not_empty_i, esbit_fifo_not_empty_i,
                            !bypass_mode_i & postht_fifo_not_empty_i};
  assign data_in_flight = |fifo_timer_q && |fifos_not_empty;

  // Extend the enable by at least one clock to give the FSM time to receive any last
  // Health checks.
  assign extend_enable = ((fifo_timer_q[0] | data_in_flight) & ~enable_i);

  // Pulse to extend from the falling edge of the incoming enable pulse
  // until one cycle after the SHA is done.
  assign sha3_active_post_en_d = cs_aes_halt_req_i && !enable_i ? 1'b1 :
                                 mubi4_test_true_strict(sha3_done_q) ? 1'b0 :
                                 sha3_active_post_en_q;

  // Force the output to be low until sha3_active_post_en_q falls or
  // for one more cycle after the falling each of extend_enable
  assign suppress_reenable = sha3_active_post_en_q | extend_enable_q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src core module
//

module entropy_src_core import entropy_src_pkg::*; #(
  parameter int EsFifoDepth = 4
) (
  input logic clk_i,
  input logic rst_ni,

  input  entropy_src_reg_pkg::entropy_src_reg2hw_t reg2hw,
  output entropy_src_reg_pkg::entropy_src_hw2reg_t hw2reg,

  // Efuse Interface
  input prim_mubi_pkg::mubi8_t otp_en_entropy_src_fw_read_i,
  input prim_mubi_pkg::mubi8_t otp_en_entropy_src_fw_over_i,

  // RNG Interface
  output logic rng_fips_o,

  // Entropy Interface
  input  entropy_src_hw_if_req_t entropy_src_hw_if_i,
  output entropy_src_hw_if_rsp_t entropy_src_hw_if_o,

  // RNG Interface
  output entropy_src_rng_req_t entropy_src_rng_o,
  input  entropy_src_rng_rsp_t entropy_src_rng_i,

  // CSRNG Interface
  output cs_aes_halt_req_t cs_aes_halt_o,
  input  cs_aes_halt_rsp_t cs_aes_halt_i,

  // External Health Test Interface
  output entropy_src_xht_req_t entropy_src_xht_o,
  input  entropy_src_xht_rsp_t entropy_src_xht_i,

  output logic           recov_alert_test_o,
  output logic           fatal_alert_test_o,
  output logic           recov_alert_o,
  output logic           fatal_alert_o,

  output logic           intr_es_entropy_valid_o,
  output logic           intr_es_health_test_failed_o,
  output logic           intr_es_observe_fifo_ready_o,
  output logic           intr_es_fatal_err_o
);

  import entropy_src_reg_pkg::*;
  import prim_mubi_pkg::mubi4_t;
  import prim_mubi_pkg::mubi4_test_true_strict;
  import prim_mubi_pkg::mubi4_and_hi;
  import prim_mubi_pkg::mubi4_test_false_loose;
  import prim_mubi_pkg::mubi4_test_invalid;

  localparam int Clog2EsFifoDepth = $clog2(EsFifoDepth);
  localparam int PostHTWidth = 32;
  localparam int RngBusWidth = 4;
  localparam int HalfRegWidth = 16;
  localparam int FullRegWidth = 32;
  localparam int EighthRegWidth = 4;
  localparam int SeedLen = 384;
  localparam int ObserveFifoWidth = 32;
  localparam int PreCondWidth = 64;
  localparam int Clog2ObserveFifoDepth = $clog2(ObserveFifoDepth);
  localparam int EsEnableCopies = 20;
  localparam int EsEnPulseCopies = 1;

  //-----------------------
  // SHA3parameters
  //-----------------------
  // Do not enable masking
  localparam bit Sha3EnMasking = 0;
  // derived parameter
  localparam int Sha3Share = (Sha3EnMasking) ? 2 : 1;

  // signals
  logic       fw_ov_mode;
  logic       fw_ov_mode_pfe;
  logic       fw_ov_mode_pfa;
  logic       fw_ov_wr_fifo_full;
  logic       fw_ov_mode_entropy_insert;
  logic       fw_ov_entropy_insert_pfe;
  logic       fw_ov_entropy_insert_pfa;
  logic       fw_ov_sha3_start_pfe;
  logic       fw_ov_sha3_start_pfe_q;
  logic       fw_ov_sha3_start_pfa;
  logic       fw_ov_sha3_disable_pulse;
  logic [ObserveFifoWidth-1:0] fw_ov_wr_data;
  logic       fw_ov_fifo_rd_pulse;
  logic       fw_ov_fifo_wr_pulse;
  logic       es_enable_pfa;

  logic       fips_enable_pfe;
  logic       fips_enable_pfa;

  logic       rng_bit_en;
  logic       rng_bit_enable_pfe;
  logic       rng_bit_enable_pfa;
  logic [1:0] rng_bit_sel;
  logic       rng_enable_q, rng_enable_d;
  logic       entropy_data_reg_en_pfe;
  logic       entropy_data_reg_en_pfa;
  logic       es_data_reg_rd_en;
  logic       sw_es_rd_pulse;
  logic       event_es_entropy_valid;
  logic       event_es_health_test_failed;
  logic       event_es_observe_fifo_ready;
  logic       event_es_fatal_err;
  logic       es_rng_src_valid;
  logic [RngBusWidth-1:0] es_rng_bus;

  logic [RngBusWidth-1:0] sfifo_esrng_wdata;
  logic [RngBusWidth-1:0] sfifo_esrng_rdata;
  logic                   sfifo_esrng_push;
  logic                   sfifo_esrng_pop;
  logic                   sfifo_esrng_clr;
  logic                   sfifo_esrng_full;
  logic                   sfifo_esrng_not_empty;
  logic                   sfifo_esrng_not_full;
  logic [2:0]             sfifo_esrng_err;

  logic [ObserveFifoWidth-1:0] sfifo_observe_wdata;
  logic [ObserveFifoWidth-1:0] sfifo_observe_rdata;
  logic                    sfifo_observe_push;
  logic                    sfifo_observe_pop;
  logic                    sfifo_observe_full;
  logic                    sfifo_observe_clr;
  logic                    sfifo_observe_not_empty;
  logic [Clog2ObserveFifoDepth:0] sfifo_observe_depth;
  logic [2:0]                     sfifo_observe_err;

  logic [Clog2EsFifoDepth:0] sfifo_esfinal_depth;
  logic [(1+SeedLen)-1:0] sfifo_esfinal_wdata;
  logic [(1+SeedLen)-1:0] sfifo_esfinal_rdata;
  logic                   sfifo_esfinal_push_enable;
  logic                   sfifo_esfinal_push;
  logic                   sfifo_esfinal_pop;
  logic                   sfifo_esfinal_clr;
  logic                   sfifo_esfinal_not_full;
  logic                   sfifo_esfinal_full;
  logic                   sfifo_esfinal_not_empty;
  logic [2:0]             sfifo_esfinal_err;
  logic [SeedLen-1:0]     esfinal_data;
  logic                   esfinal_fips_flag;

  logic                   any_fail_pulse;
  logic                   main_stage_push;
  logic                   main_stage_push_raw;
  logic                   bypass_stage_pop;
  logic                   boot_phase_done;
  logic [HalfRegWidth-1:0] any_fail_count;
  logic                    any_fails_cntr_err;
  logic                    alert_threshold_fail;
  logic [HalfRegWidth-1:0] alert_threshold;
  logic [HalfRegWidth-1:0] alert_threshold_inv;
  logic [Clog2ObserveFifoDepth:0] observe_fifo_thresh;
  logic                     observe_fifo_thresh_met;
  logic                     repcnt_active;
  logic                     repcnts_active;
  logic                     adaptp_active;
  logic                     bucket_active;
  logic                     markov_active;
  logic                     extht_active;
  logic                     alert_cntrs_clr;
  logic                     health_test_clr;
  logic                     health_test_done_pulse;
  logic [RngBusWidth-1:0]   health_test_esbus;
  logic                     health_test_esbus_vld;
  logic                     es_route_pfe;
  logic                     es_route_pfa;
  logic                     es_type_pfe;
  logic                     es_type_pfa;
  logic                     es_route_to_sw;
  logic                     es_bypass_to_sw;
  logic                     es_bypass_mode;
  logic                     rst_alert_cntr;
  logic                     threshold_scope;
  logic                     threshold_scope_pfe;
  logic                     threshold_scope_pfa;
  logic                     fips_compliance;

  logic [HalfRegWidth-1:0] health_test_fips_window;
  logic [HalfRegWidth-1:0] health_test_bypass_window;
  logic [HalfRegWidth-1:0] health_test_window;

  logic [HalfRegWidth-1:0] repcnt_fips_threshold;
  logic [HalfRegWidth-1:0] repcnt_fips_threshold_oneway;
  logic                    repcnt_fips_threshold_wr;
  logic [HalfRegWidth-1:0] repcnt_bypass_threshold;
  logic [HalfRegWidth-1:0] repcnt_bypass_threshold_oneway;
  logic                    repcnt_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] repcnt_threshold;
  logic [HalfRegWidth-1:0] repcnt_event_cnt;
  logic [HalfRegWidth-1:0] repcnt_event_hwm_fips;
  logic [HalfRegWidth-1:0] repcnt_event_hwm_bypass;
  logic [FullRegWidth-1:0] repcnt_total_fails;
  logic [EighthRegWidth-1:0] repcnt_fail_count;
  logic                     repcnt_fail_pulse;
  logic                     repcnt_fails_cntr_err;
  logic                     repcnt_alert_cntr_err;

  logic [HalfRegWidth-1:0] repcnts_fips_threshold;
  logic [HalfRegWidth-1:0] repcnts_fips_threshold_oneway;
  logic                    repcnts_fips_threshold_wr;
  logic [HalfRegWidth-1:0] repcnts_bypass_threshold;
  logic [HalfRegWidth-1:0] repcnts_bypass_threshold_oneway;
  logic                    repcnts_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] repcnts_threshold;
  logic [HalfRegWidth-1:0] repcnts_event_cnt;
  logic [HalfRegWidth-1:0] repcnts_event_hwm_fips;
  logic [HalfRegWidth-1:0] repcnts_event_hwm_bypass;
  logic [FullRegWidth-1:0] repcnts_total_fails;
  logic [EighthRegWidth-1:0] repcnts_fail_count;
  logic                     repcnts_fail_pulse;
  logic                     repcnts_fails_cntr_err;
  logic                     repcnts_alert_cntr_err;

  logic [HalfRegWidth-1:0] adaptp_hi_fips_threshold;
  logic [HalfRegWidth-1:0] adaptp_hi_fips_threshold_oneway;
  logic                    adaptp_hi_fips_threshold_wr;
  logic [HalfRegWidth-1:0] adaptp_hi_bypass_threshold;
  logic [HalfRegWidth-1:0] adaptp_hi_bypass_threshold_oneway;
  logic                    adaptp_hi_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] adaptp_hi_threshold;
  logic [HalfRegWidth-1:0] adaptp_lo_fips_threshold;
  logic [HalfRegWidth-1:0] adaptp_lo_fips_threshold_oneway;
  logic                    adaptp_lo_fips_threshold_wr;
  logic [HalfRegWidth-1:0] adaptp_lo_bypass_threshold;
  logic [HalfRegWidth-1:0] adaptp_lo_bypass_threshold_oneway;
  logic                    adaptp_lo_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] adaptp_lo_threshold;
  logic [HalfRegWidth-1:0] adaptp_hi_event_cnt;
  logic [HalfRegWidth-1:0] adaptp_lo_event_cnt;
  logic [HalfRegWidth-1:0] adaptp_hi_event_hwm_fips;
  logic [HalfRegWidth-1:0] adaptp_hi_event_hwm_bypass;
  logic [HalfRegWidth-1:0] adaptp_lo_event_hwm_fips;
  logic [HalfRegWidth-1:0] adaptp_lo_event_hwm_bypass;
  logic [FullRegWidth-1:0] adaptp_hi_total_fails;
  logic [FullRegWidth-1:0] adaptp_lo_total_fails;
  logic [EighthRegWidth-1:0] adaptp_hi_fail_count;
  logic [EighthRegWidth-1:0] adaptp_lo_fail_count;
  logic                     adaptp_hi_fail_pulse;
  logic                     adaptp_lo_fail_pulse;
  logic                     adaptp_hi_fails_cntr_err;
  logic                     adaptp_lo_fails_cntr_err;
  logic                     adaptp_hi_alert_cntr_err;
  logic                     adaptp_lo_alert_cntr_err;

  logic [HalfRegWidth-1:0] bucket_fips_threshold;
  logic [HalfRegWidth-1:0] bucket_fips_threshold_oneway;
  logic                    bucket_fips_threshold_wr;
  logic [HalfRegWidth-1:0] bucket_bypass_threshold;
  logic [HalfRegWidth-1:0] bucket_bypass_threshold_oneway;
  logic                    bucket_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] bucket_threshold;
  logic [HalfRegWidth-1:0] bucket_event_cnt;
  logic [HalfRegWidth-1:0] bucket_event_hwm_fips;
  logic [HalfRegWidth-1:0] bucket_event_hwm_bypass;
  logic [FullRegWidth-1:0] bucket_total_fails;
  logic [EighthRegWidth-1:0] bucket_fail_count;
  logic                     bucket_fail_pulse;
  logic                     bucket_fails_cntr_err;
  logic                     bucket_alert_cntr_err;

  logic [HalfRegWidth-1:0] markov_hi_fips_threshold;
  logic [HalfRegWidth-1:0] markov_hi_fips_threshold_oneway;
  logic                    markov_hi_fips_threshold_wr;
  logic [HalfRegWidth-1:0] markov_hi_bypass_threshold;
  logic [HalfRegWidth-1:0] markov_hi_bypass_threshold_oneway;
  logic                    markov_hi_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] markov_hi_threshold;
  logic [HalfRegWidth-1:0] markov_lo_fips_threshold;
  logic [HalfRegWidth-1:0] markov_lo_fips_threshold_oneway;
  logic                    markov_lo_fips_threshold_wr;
  logic [HalfRegWidth-1:0] markov_lo_bypass_threshold;
  logic [HalfRegWidth-1:0] markov_lo_bypass_threshold_oneway;
  logic                    markov_lo_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] markov_lo_threshold;
  logic [HalfRegWidth-1:0] markov_hi_event_cnt;
  logic [HalfRegWidth-1:0] markov_lo_event_cnt;
  logic [HalfRegWidth-1:0] markov_hi_event_hwm_fips;
  logic [HalfRegWidth-1:0] markov_hi_event_hwm_bypass;
  logic [HalfRegWidth-1:0] markov_lo_event_hwm_fips;
  logic [HalfRegWidth-1:0] markov_lo_event_hwm_bypass;
  logic [FullRegWidth-1:0] markov_hi_total_fails;
  logic [FullRegWidth-1:0] markov_lo_total_fails;
  logic [EighthRegWidth-1:0] markov_hi_fail_count;
  logic [EighthRegWidth-1:0] markov_lo_fail_count;
  logic                     markov_hi_fail_pulse;
  logic                     markov_lo_fail_pulse;
  logic                     markov_hi_fails_cntr_err;
  logic                     markov_lo_fails_cntr_err;
  logic                     markov_hi_alert_cntr_err;
  logic                     markov_lo_alert_cntr_err;

  logic [HalfRegWidth-1:0] extht_hi_fips_threshold;
  logic [HalfRegWidth-1:0] extht_hi_fips_threshold_oneway;
  logic                    extht_hi_fips_threshold_wr;
  logic [HalfRegWidth-1:0] extht_hi_bypass_threshold;
  logic [HalfRegWidth-1:0] extht_hi_bypass_threshold_oneway;
  logic                    extht_hi_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] extht_hi_threshold;
  logic [HalfRegWidth-1:0] extht_lo_fips_threshold;
  logic [HalfRegWidth-1:0] extht_lo_fips_threshold_oneway;
  logic                    extht_lo_fips_threshold_wr;
  logic [HalfRegWidth-1:0] extht_lo_bypass_threshold;
  logic [HalfRegWidth-1:0] extht_lo_bypass_threshold_oneway;
  logic                    extht_lo_bypass_threshold_wr;
  logic [HalfRegWidth-1:0] extht_lo_threshold;
  logic [HalfRegWidth-1:0] extht_event_cnt_hi;
  logic [HalfRegWidth-1:0] extht_event_cnt_lo;
  logic [HalfRegWidth-1:0] extht_hi_event_hwm_fips;
  logic [HalfRegWidth-1:0] extht_hi_event_hwm_bypass;
  logic [HalfRegWidth-1:0] extht_lo_event_hwm_fips;
  logic [HalfRegWidth-1:0] extht_lo_event_hwm_bypass;
  logic [FullRegWidth-1:0] extht_hi_total_fails;
  logic [FullRegWidth-1:0] extht_lo_total_fails;
  logic [EighthRegWidth-1:0] extht_hi_fail_count;
  logic [EighthRegWidth-1:0] extht_lo_fail_count;
  logic                     extht_hi_fail_pulse;
  logic                     extht_lo_fail_pulse;
  logic                     extht_cont_test;
  logic                     extht_hi_fails_cntr_err;
  logic                     extht_lo_fails_cntr_err;
  logic                     extht_hi_alert_cntr_err;
  logic                     extht_lo_alert_cntr_err;


  logic                     pfifo_esbit_wdata;
  logic [RngBusWidth-1:0]   pfifo_esbit_rdata;
  logic                     pfifo_esbit_not_empty;
  logic                     pfifo_esbit_not_full;
  logic                     pfifo_esbit_push;
  logic                     pfifo_esbit_clr;
  logic                     pfifo_esbit_pop;

  logic [RngBusWidth-1:0]   pfifo_postht_wdata;
  logic [PostHTWidth-1:0]   pfifo_postht_rdata;
  logic                     pfifo_postht_not_empty;
  logic                     pfifo_postht_not_full;
  logic                     pfifo_postht_push;
  logic                     pfifo_postht_clr;
  logic                     pfifo_postht_pop;

  logic [PreCondWidth-1:0]  pfifo_cond_wdata;
  logic [SeedLen-1:0]       pfifo_cond_rdata;
  logic                     pfifo_cond_not_empty;
  logic                     pfifo_cond_push;

  logic [ObserveFifoWidth-1:0] pfifo_precon_wdata;
  logic [PreCondWidth-1:0]     pfifo_precon_rdata;
  logic                        pfifo_precon_not_empty;
  logic                        pfifo_precon_not_full;
  logic                        pfifo_precon_push;
  logic                        pfifo_precon_clr;
  logic                        pfifo_precon_pop;

  logic [PostHTWidth-1:0]   pfifo_bypass_wdata;
  logic [SeedLen-1:0]       pfifo_bypass_rdata;
  logic                     pfifo_bypass_not_empty;
  logic                     pfifo_bypass_not_full;
  logic                     pfifo_bypass_push;
  logic                     pfifo_bypass_clr;
  logic                     pfifo_bypass_pop;

  logic [SeedLen-1:0]       pfifo_swread_wdata;
  logic                     pfifo_swread_not_full;
  logic [FullRegWidth-1:0]  pfifo_swread_rdata;
  logic                     pfifo_swread_not_empty;
  logic                     pfifo_swread_push;
  logic                     pfifo_swread_clr;
  logic                     pfifo_swread_pop;

  logic [SeedLen-1:0]       final_es_data;
  logic                     es_hw_if_req;
  logic                     es_hw_if_ack;
  logic                     es_hw_if_fifo_pop;
  logic                     sfifo_esrng_err_sum;
  logic                     sfifo_observe_err_sum;
  logic                     sfifo_esfinal_err_sum;
  // For fifo errors that are generated through the
  // ERR_CODE_TEST register, but are not associated
  // with any errors:
  logic                     sfifo_test_err_sum;
  logic                     es_ack_sm_err_sum;
  logic                     es_ack_sm_err;
  logic                     es_main_sm_err_sum;
  logic                     es_main_sm_err;
  logic                     es_main_sm_alert;
  logic                     es_bus_cmp_alert;
  logic                     es_thresh_cfg_alert;
  logic                     es_main_sm_idle;
  logic [8:0]               es_main_sm_state;
  logic                     fifo_write_err_sum;
  logic                     fifo_read_err_sum;
  logic                     fifo_status_err_sum;
  logic [30:0]              err_code_test_bit;
  logic                     sha3_msgfifo_ready;
  logic                     sha3_state_vld;
  logic                     sha3_start_raw;
  logic                     sha3_start;
  logic                     sha3_process;
  logic                     sha3_msg_end;
  logic                     sha3_msg_rdy_mask;
  logic                     sha3_block_processed;
  prim_mubi_pkg::mubi4_t    sha3_done;
  prim_mubi_pkg::mubi4_t    sha3_absorbed;
  logic                     sha3_squeezing;
  logic [2:0]               sha3_fsm;
  logic [32:0]              sha3_err;
  logic                     cs_aes_halt_req;
  logic                     sha3_msg_rdy;
  logic [HalfRegWidth-1:0]  window_cntr;

  logic [sha3_pkg::StateW-1:0] sha3_state[Sha3Share];
  logic [PreCondWidth-1:0] msg_data[Sha3Share];
  logic                    es_rdata_capt_vld;
  logic                    window_cntr_err;
  logic                    repcnt_cntr_err;
  logic                    repcnts_cntr_err;
  logic                    adaptp_cntr_err;
  logic                    bucket_cntr_err;
  logic                    markov_cntr_err;
  logic                    es_cntr_err;
  logic                    es_cntr_err_sum;
  logic                    sha3_state_error_sum;
  logic                    sha3_rst_storage_err_sum;
  logic                    efuse_es_sw_reg_en;
  logic                    efuse_es_sw_ov_en;

  logic                    sha3_state_error;
  logic                    sha3_count_error;
  logic                    sha3_rst_storage_err;
  logic                    es_hw_regwen;
  logic                    recov_alert_state;
  logic                    es_fw_ov_wr_alert;
  logic                    es_fw_ov_disable_alert;
  logic                    fw_ov_corrupted;

  logic                    stale_seed_processing;
  logic                    main_sm_enable;

  logic                    unused_err_code_test_bit;
  logic                    unused_sha3_state;
  logic                    unused_entropy_data;
  logic                    unused_fw_ov_rd_data;

  prim_mubi_pkg::mubi8_t en_entropy_src_fw_read;
  prim_mubi_pkg::mubi8_t en_entropy_src_fw_over;

  mubi4_t mubi_es_enable;
  mubi4_t mubi_module_en_pulse;

  mubi4_t       mubi_module_en_raw;
  mubi4_t [2:0] mubi_module_en_raw_fanout;

  mubi4_t [EsEnableCopies-1:0] mubi_es_enable_fanout;
  logic   [EsEnableCopies-1:0] es_enable_fo;

  mubi4_t [EsEnPulseCopies-1:0] mubi_module_en_pulse_fanout;
  logic   [EsEnPulseCopies-1:0] module_en_pulse_fo;

  // A delayed copy of the enable signal, and enable pulse which are needed to cleanly handle any
  // long-duration operations from the previous run.
  logic                        es_delayed_enable;

  mubi4_t [1:0] mubi_rng_bit_en_fanout;
  mubi4_t mubi_rng_bit_en;

  // flops
  logic        ht_failed_q, ht_failed_d;
  logic        ht_done_pulse_q, ht_done_pulse_d;
  logic        sha3_err_q, sha3_err_d;
  logic        cs_aes_halt_q, cs_aes_halt_d;
  logic [63:0] es_rdata_capt_q, es_rdata_capt_d;
  logic        es_rdata_capt_vld_q, es_rdata_capt_vld_d;
  logic        sha3_msg_rdy_mask_q, sha3_msg_rdy_mask_d;
  mubi4_t      mubi_mod_en_dly_d, mubi_mod_en_dly_q;


  logic        sha3_start_mask_q, sha3_start_mask_d;
  logic        sha3_flush_q, sha3_flush_d;
  logic [1:0]  fw_ov_corrupted_q, fw_ov_corrupted_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      ht_failed_q            <= '0;
      ht_done_pulse_q        <= '0;
      sha3_err_q             <= '0;
      cs_aes_halt_q          <= '0;
      es_rdata_capt_q        <= '0;
      es_rdata_capt_vld_q    <= '0;
      fw_ov_sha3_start_pfe_q <= '0;
      sha3_msg_rdy_mask_q    <= '0;
      mubi_mod_en_dly_q      <= prim_mubi_pkg::MuBi4False;
      sha3_flush_q           <= '0;
      sha3_start_mask_q      <= '0;
      fw_ov_corrupted_q      <= 2'b00;
      rng_enable_q           <= 1'b 0;
    end else begin
      ht_failed_q            <= ht_failed_d;
      ht_done_pulse_q        <= ht_done_pulse_d;
      sha3_err_q             <= sha3_err_d;
      cs_aes_halt_q          <= cs_aes_halt_d;
      es_rdata_capt_q        <= es_rdata_capt_d;
      es_rdata_capt_vld_q    <= es_rdata_capt_vld_d;
      fw_ov_sha3_start_pfe_q <= fw_ov_sha3_start_pfe;
      sha3_msg_rdy_mask_q    <= sha3_msg_rdy_mask_d;
      sha3_flush_q           <= sha3_flush_d;
      sha3_start_mask_q      <= sha3_start_mask_d;
      mubi_mod_en_dly_q      <= mubi_mod_en_dly_d;
      fw_ov_corrupted_q      <= fw_ov_corrupted_d;
      rng_enable_q           <= rng_enable_d;
    end
  end

  assign fw_ov_sha3_disable_pulse = fw_ov_sha3_start_pfe_q & ~fw_ov_sha3_start_pfe;

  //--------------------------------------------
  // register lock gating
  //--------------------------------------------

  // Allow writes only if
  // 1. SW_REGUPD is true,
  // 2. The DUT is disabled
  //   Block writes if enabled or if internal activities are still in progress (as indicated by
  //   es_delayed_enable).
  assign es_hw_regwen = reg2hw.sw_regupd.q &&
                        mubi4_test_false_loose(mubi_module_en_raw_fanout[0]) &&
                        !es_delayed_enable;
  assign hw2reg.regwen.de = 1'b1;
  assign hw2reg.regwen.d = es_hw_regwen;

  //--------------------------------------------
  // set up secure enable bits
  //--------------------------------------------

  // check for illegal enable field states, and set alert if detected

  // SEC_CM: CONFIG.MUBI
  assign mubi_module_en_raw = mubi4_t'(reg2hw.module_enable.q);
  assign es_enable_pfa      = mubi4_test_invalid(mubi_module_en_raw_fanout[1]);
  assign hw2reg.recov_alert_sts.module_enable_field_alert.de = es_enable_pfa;
  assign hw2reg.recov_alert_sts.module_enable_field_alert.d  = es_enable_pfa;

  prim_mubi4_sync #(
    .NumCopies(3),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_entropy_module_en (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_module_en_raw),
    .mubi_o(mubi_module_en_raw_fanout)
  );

  // Generation of enable pulse, and main enable signals.
  //
  // This module creates a single mubi_encoded module_enable_pulse, as well as
  // a general mubi_es_enable signal.
  //
  // The module enable pulse is MuBi4True for a single clock after the
  // module_enable register is asserted MuBi4True. However in this first clock cycle
  // most of the module is not enabled.  (The enable pulse is for clearing the
  // residual internal state.)
  //
  // The rest of the module is enabled in the second clock cycle after seting the
  // module_enable register to MuBi4True.
  //
  // When module_enable is set to MuBi4False the module is disabled.  No further
  // RNG input is accepted and the state machines transition to Idle as soon as
  // possible. Some delay may occur if the SHA3 conditioning block is busy, though
  // otherwise the main_sm transitions to Idle without delay.

  assign mubi_mod_en_dly_d = mubi_module_en_raw_fanout[2];
  assign mubi_module_en_pulse = mubi4_and_hi(mubi_mod_en_dly_d, mubi4_t'(~mubi_mod_en_dly_q));
  assign mubi_es_enable = mubi4_and_hi(mubi_mod_en_dly_d, mubi_mod_en_dly_q);

  for (genvar i = 0; i < EsEnableCopies; i = i+1) begin : gen_mubi_en_copies
    assign es_enable_fo[i] = mubi4_test_true_strict(mubi_es_enable_fanout[i]);
  end : gen_mubi_en_copies

  prim_mubi4_sync #(
    .NumCopies(EsEnableCopies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_es_enable (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_es_enable),
    .mubi_o(mubi_es_enable_fanout)
  );

  for (genvar i = 0; i < EsEnPulseCopies; i = i+1) begin : gen_mubi_en_pulse_copies
    assign module_en_pulse_fo[i] = mubi4_test_true_strict(mubi_module_en_pulse_fanout[i]);
  end : gen_mubi_en_pulse_copies

  prim_mubi4_sync #(
    .NumCopies(EsEnPulseCopies),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_es_enable_pulse (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_module_en_pulse),
    .mubi_o(mubi_module_en_pulse_fanout)
  );

  entropy_src_enable_delay u_enable_delay (
    .clk_i,
    .rst_ni,
    .enable_i(es_enable_fo[0]),
    .esrng_fifo_not_empty_i(sfifo_esrng_not_empty),
    .esbit_fifo_not_empty_i(pfifo_esbit_not_empty),
    .postht_fifo_not_empty_i(pfifo_postht_not_empty),
    .cs_aes_halt_req_i(cs_aes_halt_req),
    .sha3_done_i(sha3_done),
    .bypass_mode_i(es_bypass_mode),
    .enable_o(es_delayed_enable)
  );

  mubi4_t mubi_fips_en;
  mubi4_t [1:0] mubi_fips_en_fanout;
  assign mubi_fips_en  = mubi4_t'(reg2hw.conf.fips_enable.q);
  assign fips_enable_pfe = mubi4_test_true_strict(mubi_fips_en_fanout[0]);
  assign fips_enable_pfa = mubi4_test_invalid(mubi_fips_en_fanout[1]);
  assign hw2reg.recov_alert_sts.fips_enable_field_alert.de = fips_enable_pfa;
  assign hw2reg.recov_alert_sts.fips_enable_field_alert.d  = fips_enable_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_entropy_fips_en (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_fips_en),
    .mubi_o(mubi_fips_en_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_entropy_reg_en;
  mubi4_t [1:0] mubi_entropy_reg_en_fanout;
  assign mubi_entropy_reg_en = mubi4_t'(reg2hw.conf.entropy_data_reg_enable.q);
  assign entropy_data_reg_en_pfe = mubi4_test_true_strict(mubi_entropy_reg_en_fanout[0]);
  assign entropy_data_reg_en_pfa = mubi4_test_invalid(mubi_entropy_reg_en_fanout[1]);
  assign hw2reg.recov_alert_sts.entropy_data_reg_en_field_alert.de = entropy_data_reg_en_pfa;
  assign hw2reg.recov_alert_sts.entropy_data_reg_en_field_alert.d =  entropy_data_reg_en_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_entropy_data_reg_en (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_entropy_reg_en),
    .mubi_o(mubi_entropy_reg_en_fanout)
  );

  assign observe_fifo_thresh = reg2hw.observe_fifo_thresh.q;

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_fw_ov_mode;
  mubi4_t [1:0] mubi_fw_ov_mode_fanout;
  assign mubi_fw_ov_mode = mubi4_t'(reg2hw.fw_ov_control.fw_ov_mode.q);
  assign fw_ov_mode_pfe = mubi4_test_true_strict(mubi_fw_ov_mode_fanout[0]);
  assign fw_ov_mode_pfa = mubi4_test_invalid(mubi_fw_ov_mode_fanout[1]);
  assign hw2reg.recov_alert_sts.fw_ov_mode_field_alert.de = fw_ov_mode_pfa;
  assign hw2reg.recov_alert_sts.fw_ov_mode_field_alert.d  = fw_ov_mode_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_fw_ov_mode (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_fw_ov_mode),
    .mubi_o(mubi_fw_ov_mode_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_fw_ov_entropy_insert;
  mubi4_t [1:0] mubi_fw_ov_entropy_insert_fanout;
  assign mubi_fw_ov_entropy_insert = mubi4_t'(reg2hw.fw_ov_control.fw_ov_entropy_insert.q);
  assign fw_ov_entropy_insert_pfe = mubi4_test_true_strict(mubi_fw_ov_entropy_insert_fanout[0]);
  assign fw_ov_entropy_insert_pfa = mubi4_test_invalid(mubi_fw_ov_entropy_insert_fanout[1]);
  assign hw2reg.recov_alert_sts.fw_ov_entropy_insert_field_alert.de = fw_ov_entropy_insert_pfa;
  assign hw2reg.recov_alert_sts.fw_ov_entropy_insert_field_alert.d  = fw_ov_entropy_insert_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_fw_ov_entropy_insert (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_fw_ov_entropy_insert),
    .mubi_o(mubi_fw_ov_entropy_insert_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_fw_ov_sha3_start;
  mubi4_t [1:0] mubi_fw_ov_sha3_start_fanout;
  assign mubi_fw_ov_sha3_start = mubi4_t'(reg2hw.fw_ov_sha3_start.q);
  assign fw_ov_sha3_start_pfe = mubi4_test_true_strict(mubi_fw_ov_sha3_start_fanout[0]);
  assign fw_ov_sha3_start_pfa = mubi4_test_invalid(mubi_fw_ov_sha3_start_fanout[1]);
  assign hw2reg.recov_alert_sts.fw_ov_sha3_start_field_alert.de = fw_ov_sha3_start_pfa;
  assign hw2reg.recov_alert_sts.fw_ov_sha3_start_field_alert.d  = fw_ov_sha3_start_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_fw_ov_sha3_start (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_fw_ov_sha3_start),
    .mubi_o(mubi_fw_ov_sha3_start_fanout)
  );

  // firmware override controls
  assign fw_ov_mode = efuse_es_sw_ov_en && fw_ov_mode_pfe;
  assign fw_ov_mode_entropy_insert = fw_ov_mode && fw_ov_entropy_insert_pfe;
  assign fw_ov_fifo_rd_pulse = reg2hw.fw_ov_rd_data.re;
  assign hw2reg.fw_ov_rd_data.d = sfifo_observe_rdata;
  assign fw_ov_fifo_wr_pulse = reg2hw.fw_ov_wr_data.qe;
  assign fw_ov_wr_data = reg2hw.fw_ov_wr_data.q;

  assign efuse_es_sw_ov_en = prim_mubi_pkg::mubi8_test_true_strict(en_entropy_src_fw_over);

  prim_mubi8_sync #(
    .NumCopies(1),
    .AsyncOn(1) // must be set to one, see note below
  ) u_prim_mubi8_sync_es_fw_over (
    .clk_i,
    .rst_ni,
    .mubi_i(otp_en_entropy_src_fw_over_i),
    .mubi_o({en_entropy_src_fw_over})
  );

  // note: the input to the above sync module is from the OTP block.
  //       It is assumed that the source is in a different time domain,
  //       and requires the AsyncOn parameter to be set.

  // rng_enable is being used in other clock domains. Need to latch the
  // signal.
  assign rng_enable_d = es_enable_fo[1] &&
                        es_delayed_enable &&
                        sfifo_esrng_not_full;

  assign entropy_src_rng_o.rng_enable = rng_enable_q;

  assign es_rng_src_valid = entropy_src_rng_i.rng_valid;
  assign es_rng_bus = entropy_src_rng_i.rng_b;


  //--------------------------------------------
  // instantiate interrupt hardware primitives
  //--------------------------------------------

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_es_entropy_valid (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_es_entropy_valid),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.es_entropy_valid.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.es_entropy_valid.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.es_entropy_valid.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.es_entropy_valid.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.es_entropy_valid.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.es_entropy_valid.d),
    .intr_o                 (intr_es_entropy_valid_o)
  );

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_es_health_test_failed (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_es_health_test_failed),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.es_health_test_failed.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.es_health_test_failed.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.es_health_test_failed.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.es_health_test_failed.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.es_health_test_failed.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.es_health_test_failed.d),
    .intr_o                 (intr_es_health_test_failed_o)
  );


  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_es_observe_fifo_ready (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_es_observe_fifo_ready),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.es_observe_fifo_ready.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.es_observe_fifo_ready.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.es_observe_fifo_ready.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.es_observe_fifo_ready.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.es_observe_fifo_ready.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.es_observe_fifo_ready.d),
    .intr_o                 (intr_es_observe_fifo_ready_o)
  );

  prim_intr_hw #(
    .Width(1)
  ) u_intr_hw_es_fatal_err (
    .clk_i                  (clk_i),
    .rst_ni                 (rst_ni),
    .event_intr_i           (event_es_fatal_err),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.es_fatal_err.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.es_fatal_err.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.es_fatal_err.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.es_fatal_err.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.es_fatal_err.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.es_fatal_err.d),
    .intr_o                 (intr_es_fatal_err_o)
  );

  //--------------------------------------------
  // tlul register settings
  //--------------------------------------------


  // set the interrupt event when enabled
  assign event_es_entropy_valid = pfifo_swread_not_empty && es_enable_fo[2];


  // set the interrupt sources
  assign event_es_fatal_err = (es_enable_fo[3] &&
                                 (sfifo_esrng_err_sum   ||
                                  sfifo_observe_err_sum ||
                                  sfifo_esfinal_err_sum ||
                                  sfifo_test_err_sum) ) ||
                              es_ack_sm_err_sum ||
                              es_main_sm_err_sum ||
                              es_cntr_err_sum || // prim_count err is always active
                              sha3_rst_storage_err_sum ||
                              sha3_state_error_sum;

  // set fifo errors that are single instances of source
  assign sfifo_esrng_err_sum = (|sfifo_esrng_err) ||
         err_code_test_bit[0];
  assign sfifo_observe_err_sum = (|sfifo_observe_err) ||
         err_code_test_bit[1];
  assign sfifo_esfinal_err_sum = (|sfifo_esfinal_err) ||
         err_code_test_bit[2];

  // The following test bits help normally diagnose the _type_ of
  // error when they are triggred by the fifo. However when
  // they are triggered by softwre they are not linked to a
  // particular sfifo and do not trigger an alert, unless
  // we capture them here.
  assign sfifo_test_err_sum = err_code_test_bit[28] ||
                              err_code_test_bit[29] ||
                              err_code_test_bit[30];

  assign es_ack_sm_err_sum = es_ack_sm_err ||
         err_code_test_bit[20];
  assign es_main_sm_err_sum = es_main_sm_err ||
         err_code_test_bit[21];
  assign es_cntr_err_sum = es_cntr_err ||
         err_code_test_bit[22];
  assign sha3_state_error_sum = sha3_state_error ||
         err_code_test_bit[23];
  assign sha3_rst_storage_err_sum = sha3_rst_storage_err ||
         err_code_test_bit[24];
  assign fifo_write_err_sum =
         sfifo_esrng_err[2] ||
         sfifo_observe_err[2] ||
         sfifo_esfinal_err[2] ||
         err_code_test_bit[28];
  assign fifo_read_err_sum =
         sfifo_esrng_err[1] ||
         sfifo_observe_err[1] ||
         sfifo_esfinal_err[1] ||
         err_code_test_bit[29];
  assign fifo_status_err_sum =
         sfifo_esrng_err[0] ||
         sfifo_observe_err[0] ||
         sfifo_esfinal_err[0] ||
         err_code_test_bit[30];

  // set the err code source bits
  assign hw2reg.err_code.sfifo_esrng_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_esrng_err.de = sfifo_esrng_err_sum;

  assign hw2reg.err_code.sfifo_observe_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_observe_err.de = sfifo_observe_err_sum;

  assign hw2reg.err_code.sfifo_esfinal_err.d = 1'b1;
  assign hw2reg.err_code.sfifo_esfinal_err.de = sfifo_esfinal_err_sum;

  assign hw2reg.err_code.es_ack_sm_err.d = 1'b1;
  assign hw2reg.err_code.es_ack_sm_err.de = es_ack_sm_err_sum;

  assign hw2reg.err_code.es_main_sm_err.d = 1'b1;
  assign hw2reg.err_code.es_main_sm_err.de = es_main_sm_err_sum;

  assign hw2reg.err_code.es_cntr_err.d = 1'b1;
  assign hw2reg.err_code.es_cntr_err.de = es_cntr_err_sum;

  assign hw2reg.err_code.sha3_state_err.d = 1'b1;
  assign hw2reg.err_code.sha3_state_err.de = sha3_state_error_sum;

  assign hw2reg.err_code.sha3_rst_storage_err.d = 1'b1;
  assign hw2reg.err_code.sha3_rst_storage_err.de = sha3_rst_storage_err_sum;


 // set the err code type bits
  assign hw2reg.err_code.fifo_write_err.d = 1'b1;
  assign hw2reg.err_code.fifo_write_err.de = fifo_write_err_sum;

  assign hw2reg.err_code.fifo_read_err.d = 1'b1;
  assign hw2reg.err_code.fifo_read_err.de = fifo_read_err_sum;

  assign hw2reg.err_code.fifo_state_err.d = 1'b1;
  assign hw2reg.err_code.fifo_state_err.de = fifo_status_err_sum;

  // Error forcing
  for (genvar i = 0; i < 31; i = i+1) begin : gen_err_code_test_bit
    assign err_code_test_bit[i] = (reg2hw.err_code_test.q == i) && reg2hw.err_code_test.qe;
  end : gen_err_code_test_bit

  // alert - send all interrupt sources to the alert for the fatal case
  assign fatal_alert_o = event_es_fatal_err;

  // alert test
  assign recov_alert_test_o = {
    reg2hw.alert_test.recov_alert.q &&
    reg2hw.alert_test.recov_alert.qe
  };
  assign fatal_alert_test_o = {
    reg2hw.alert_test.fatal_alert.q &&
    reg2hw.alert_test.fatal_alert.qe
  };


  // set the debug status reg
  assign hw2reg.debug_status.entropy_fifo_depth.d = sfifo_esfinal_depth;
  assign hw2reg.debug_status.sha3_fsm.d = sha3_fsm;
  assign hw2reg.debug_status.sha3_block_pr.d = sha3_block_processed;
  assign hw2reg.debug_status.sha3_squeezing.d = sha3_squeezing;
  assign hw2reg.debug_status.sha3_absorbed.d =
    prim_mubi_pkg::mubi4_test_true_strict(sha3_absorbed) ? 1'b 1 : 1'b 0;
  assign hw2reg.debug_status.sha3_err.d = sha3_err_q;

  assign sha3_err_d =
         es_enable_fo[4] ? 1'b0 :
         {|sha3_err} ? 1'b1 :
         sha3_err_q;

  // state machine status
  assign hw2reg.debug_status.main_sm_idle.d = es_main_sm_idle;
  assign hw2reg.debug_status.main_sm_boot_done.d = boot_phase_done;
  assign hw2reg.main_sm_state.de = 1'b1;
  assign hw2reg.main_sm_state.d = es_main_sm_state;

  // fw override wr data status indication
  assign fw_ov_wr_fifo_full = fw_ov_mode_entropy_insert &&
                              (es_bypass_mode ? !pfifo_bypass_not_full : !pfifo_precon_not_full);

  assign hw2reg.fw_ov_wr_fifo_full.d = fw_ov_wr_fifo_full;


  //--------------------------------------------
  // receive in RNG bus input
  //--------------------------------------------


  prim_fifo_sync #(
    .Width(RngBusWidth),
    .Pass(0),
    .Depth(2),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_esrng (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (sfifo_esrng_clr),
    .wvalid_i   (sfifo_esrng_push),
    .wdata_i    (sfifo_esrng_wdata),
    .wready_o   (sfifo_esrng_not_full),
    .rvalid_o   (sfifo_esrng_not_empty),
    .rdata_o    (sfifo_esrng_rdata),
    .rready_i   (sfifo_esrng_pop),
    .full_o     (sfifo_esrng_full),
    .depth_o    (),
    .err_o      ()
  );

  // fifo controls
  assign sfifo_esrng_push = es_enable_fo[5] && es_delayed_enable && es_rng_src_valid &&
                            rng_enable_q;

  assign sfifo_esrng_clr   = ~es_delayed_enable;
  assign sfifo_esrng_wdata = es_rng_bus;
  assign sfifo_esrng_pop   = sfifo_esrng_not_empty & (rng_bit_en ? pfifo_esbit_not_full :
                                                                   pfifo_postht_not_full );

  // fifo err
  // Note: for prim_fifo_sync is not an error to push to a fifo that is full.  In fact, the
  // backpressure mechanism applied to the RNG inputs counts on this.
  assign sfifo_esrng_err =
         {1'b0,
          (sfifo_esrng_pop && !sfifo_esrng_not_empty),
          (sfifo_esrng_full && !sfifo_esrng_not_empty)};


  // pack esrng bus into signal bit packer

  // SEC_CM: CONFIG.MUBI
  assign mubi_rng_bit_en = mubi4_t'(reg2hw.conf.rng_bit_enable.q);
  assign rng_bit_enable_pfe = mubi4_test_true_strict(mubi_rng_bit_en_fanout[0]);
  assign rng_bit_enable_pfa = mubi4_test_invalid(mubi_rng_bit_en_fanout[1]);
  assign hw2reg.recov_alert_sts.rng_bit_enable_field_alert.de = rng_bit_enable_pfa;
  assign hw2reg.recov_alert_sts.rng_bit_enable_field_alert.d  = rng_bit_enable_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_rng_bit_en (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_rng_bit_en),
    .mubi_o(mubi_rng_bit_en_fanout)
  );


  assign rng_bit_en = rng_bit_enable_pfe;
  assign rng_bit_sel = reg2hw.conf.rng_bit_sel.q;

  prim_packer_fifo #(
    .InW(1),
    .OutW(RngBusWidth),
    .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_esbit (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (pfifo_esbit_clr),
    .wvalid_i   (pfifo_esbit_push),
    .wdata_i    (pfifo_esbit_wdata),
    .wready_o   (pfifo_esbit_not_full),
    .rvalid_o   (pfifo_esbit_not_empty),
    .rdata_o    (pfifo_esbit_rdata),
    .rready_i   (pfifo_esbit_pop),
    .depth_o    ()
  );

  assign pfifo_esbit_push = rng_bit_en && sfifo_esrng_not_empty;
  assign pfifo_esbit_clr = ~es_delayed_enable;
  assign pfifo_esbit_pop = rng_bit_en && pfifo_esbit_not_empty && pfifo_postht_not_full;
  assign pfifo_esbit_wdata =
         (rng_bit_sel == 2'h0) ? sfifo_esrng_rdata[0] :
         (rng_bit_sel == 2'h1) ? sfifo_esrng_rdata[1] :
         (rng_bit_sel == 2'h2) ? sfifo_esrng_rdata[2] :
         sfifo_esrng_rdata[3];


  // select source for health testing

  assign health_test_esbus     = pfifo_postht_wdata;
  assign health_test_esbus_vld = pfifo_postht_push & pfifo_postht_not_full & ~pfifo_postht_clr;

  // Health test any data that comes in on the RNG interface.
  assign repcnt_active = 1'b1;
  assign repcnts_active = 1'b1;
  assign adaptp_active = 1'b1;
  assign bucket_active = 1'b1;
  assign markov_active = 1'b1;
  assign extht_active = 1'b1;

  // Only reset health tests on re-enable
  assign health_test_clr = module_en_pulse_fo[0];

  assign health_test_fips_window = reg2hw.health_test_windows.fips_window.q;
  assign health_test_bypass_window = reg2hw.health_test_windows.bypass_window.q;

  assign repcnt_fips_threshold = reg2hw.repcnt_thresholds.fips_thresh.q;
  assign repcnt_fips_threshold_wr = reg2hw.repcnt_thresholds.fips_thresh.qe;
  assign hw2reg.repcnt_thresholds.fips_thresh.d = repcnt_fips_threshold_oneway;
  assign repcnt_bypass_threshold = reg2hw.repcnt_thresholds.bypass_thresh.q;
  assign repcnt_bypass_threshold_wr = reg2hw.repcnt_thresholds.bypass_thresh.qe;
  assign hw2reg.repcnt_thresholds.bypass_thresh.d = repcnt_bypass_threshold_oneway;

  assign repcnts_fips_threshold = reg2hw.repcnts_thresholds.fips_thresh.q;
  assign repcnts_fips_threshold_wr = reg2hw.repcnts_thresholds.fips_thresh.qe;
  assign hw2reg.repcnts_thresholds.fips_thresh.d = repcnts_fips_threshold_oneway;
  assign repcnts_bypass_threshold = reg2hw.repcnts_thresholds.bypass_thresh.q;
  assign repcnts_bypass_threshold_wr = reg2hw.repcnts_thresholds.bypass_thresh.qe;
  assign hw2reg.repcnts_thresholds.bypass_thresh.d = repcnts_bypass_threshold_oneway;


  assign adaptp_hi_fips_threshold = reg2hw.adaptp_hi_thresholds.fips_thresh.q;
  assign adaptp_hi_fips_threshold_wr = reg2hw.adaptp_hi_thresholds.fips_thresh.qe;
  assign hw2reg.adaptp_hi_thresholds.fips_thresh.d = adaptp_hi_fips_threshold_oneway;
  assign adaptp_hi_bypass_threshold = reg2hw.adaptp_hi_thresholds.bypass_thresh.q;
  assign adaptp_hi_bypass_threshold_wr = reg2hw.adaptp_hi_thresholds.bypass_thresh.qe;
  assign hw2reg.adaptp_hi_thresholds.bypass_thresh.d = adaptp_hi_bypass_threshold_oneway;

  assign adaptp_lo_fips_threshold = reg2hw.adaptp_lo_thresholds.fips_thresh.q;
  assign adaptp_lo_fips_threshold_wr = reg2hw.adaptp_lo_thresholds.fips_thresh.qe;
  assign hw2reg.adaptp_lo_thresholds.fips_thresh.d = adaptp_lo_fips_threshold_oneway;
  assign adaptp_lo_bypass_threshold = reg2hw.adaptp_lo_thresholds.bypass_thresh.q;
  assign adaptp_lo_bypass_threshold_wr = reg2hw.adaptp_lo_thresholds.bypass_thresh.qe;
  assign hw2reg.adaptp_lo_thresholds.bypass_thresh.d = adaptp_lo_bypass_threshold_oneway;


  assign bucket_fips_threshold = reg2hw.bucket_thresholds.fips_thresh.q;
  assign bucket_fips_threshold_wr = reg2hw.bucket_thresholds.fips_thresh.qe;
  assign hw2reg.bucket_thresholds.fips_thresh.d = bucket_fips_threshold_oneway;
  assign bucket_bypass_threshold = reg2hw.bucket_thresholds.bypass_thresh.q;
  assign bucket_bypass_threshold_wr = reg2hw.bucket_thresholds.bypass_thresh.qe;
  assign hw2reg.bucket_thresholds.bypass_thresh.d = bucket_bypass_threshold_oneway;


  assign markov_hi_fips_threshold = reg2hw.markov_hi_thresholds.fips_thresh.q;
  assign markov_hi_fips_threshold_wr = reg2hw.markov_hi_thresholds.fips_thresh.qe;
  assign hw2reg.markov_hi_thresholds.fips_thresh.d = markov_hi_fips_threshold_oneway;
  assign markov_hi_bypass_threshold = reg2hw.markov_hi_thresholds.bypass_thresh.q;
  assign markov_hi_bypass_threshold_wr = reg2hw.markov_hi_thresholds.bypass_thresh.qe;
  assign hw2reg.markov_hi_thresholds.bypass_thresh.d = markov_hi_bypass_threshold_oneway;

  assign markov_lo_fips_threshold = reg2hw.markov_lo_thresholds.fips_thresh.q;
  assign markov_lo_fips_threshold_wr = reg2hw.markov_lo_thresholds.fips_thresh.qe;
  assign hw2reg.markov_lo_thresholds.fips_thresh.d = markov_lo_fips_threshold_oneway;
  assign markov_lo_bypass_threshold = reg2hw.markov_lo_thresholds.bypass_thresh.q;
  assign markov_lo_bypass_threshold_wr = reg2hw.markov_lo_thresholds.bypass_thresh.qe;
  assign hw2reg.markov_lo_thresholds.bypass_thresh.d = markov_lo_bypass_threshold_oneway;


  assign extht_hi_fips_threshold = reg2hw.extht_hi_thresholds.fips_thresh.q;
  assign extht_hi_fips_threshold_wr = reg2hw.extht_hi_thresholds.fips_thresh.qe;
  assign hw2reg.extht_hi_thresholds.fips_thresh.d = extht_hi_fips_threshold_oneway;
  assign extht_hi_bypass_threshold = reg2hw.extht_hi_thresholds.bypass_thresh.q;
  assign extht_hi_bypass_threshold_wr = reg2hw.extht_hi_thresholds.bypass_thresh.qe;
  assign hw2reg.extht_hi_thresholds.bypass_thresh.d = extht_hi_bypass_threshold_oneway;

  assign extht_lo_fips_threshold = reg2hw.extht_lo_thresholds.fips_thresh.q;
  assign extht_lo_fips_threshold_wr = reg2hw.extht_lo_thresholds.fips_thresh.qe;
  assign hw2reg.extht_lo_thresholds.fips_thresh.d = extht_lo_fips_threshold_oneway;
  assign extht_lo_bypass_threshold = reg2hw.extht_lo_thresholds.bypass_thresh.q;
  assign extht_lo_bypass_threshold_wr = reg2hw.extht_lo_thresholds.bypass_thresh.qe;
  assign hw2reg.extht_lo_thresholds.bypass_thresh.d = extht_lo_bypass_threshold_oneway;



  assign health_test_window = es_bypass_mode ? health_test_bypass_window : health_test_fips_window;

  // Window sizes other than 384 bits (the seed length) are currently not tested nor supported in
  // bypass or boot-time mode.
  `ASSERT(EsBootTimeHtWindowSizeSupported_A,
      main_sm_enable && es_bypass_mode && !fw_ov_mode_entropy_insert
      |-> health_test_bypass_window == HalfRegWidth'(SeedLen/4))

  //------------------------------
  // repcnt one-way thresholds
  //------------------------------
  assign repcnt_threshold = es_bypass_mode ? repcnt_bypass_threshold_oneway :
         repcnt_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_repcnt_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (repcnt_fips_threshold_wr),
    .value_i             (repcnt_fips_threshold),
    .value_o             (repcnt_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_repcnt_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (repcnt_bypass_threshold_wr),
    .value_i             (repcnt_bypass_threshold),
    .value_o             (repcnt_bypass_threshold_oneway)
  );

  //------------------------------
  // repcnts one-way thresholds
  //------------------------------
  assign repcnts_threshold = es_bypass_mode ? repcnts_bypass_threshold_oneway :
         repcnts_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_repcnts_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (repcnts_fips_threshold_wr),
    .value_i             (repcnts_fips_threshold),
    .value_o             (repcnts_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_repcnts_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (repcnts_bypass_threshold_wr),
    .value_i             (repcnts_bypass_threshold),
    .value_o             (repcnts_bypass_threshold_oneway)
  );


  //------------------------------
  // adaptp one-way thresholds
  //------------------------------
  assign adaptp_hi_threshold = es_bypass_mode ? adaptp_hi_bypass_threshold_oneway :
         adaptp_hi_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_adaptp_hi_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (adaptp_hi_fips_threshold_wr),
    .value_i             (adaptp_hi_fips_threshold),
    .value_o             (adaptp_hi_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_adaptp_hi_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (adaptp_hi_bypass_threshold_wr),
    .value_i             (adaptp_hi_bypass_threshold),
    .value_o             (adaptp_hi_bypass_threshold_oneway)
  );

  assign adaptp_lo_threshold = es_bypass_mode ? adaptp_lo_bypass_threshold_oneway :
         adaptp_lo_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_adaptp_lo_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (adaptp_lo_fips_threshold_wr),
    .value_i             (adaptp_lo_fips_threshold),
    .value_o             (adaptp_lo_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_adaptp_lo_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (adaptp_lo_bypass_threshold_wr),
    .value_i             (adaptp_lo_bypass_threshold),
    .value_o             (adaptp_lo_bypass_threshold_oneway)
  );


  //------------------------------
  // bucket one-way thresholds
  //------------------------------
  assign bucket_threshold = es_bypass_mode ? bucket_bypass_threshold_oneway :
         bucket_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_bucket_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (bucket_fips_threshold_wr),
    .value_i             (bucket_fips_threshold),
    .value_o             (bucket_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_bucket_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (bucket_bypass_threshold_wr),
    .value_i             (bucket_bypass_threshold),
    .value_o             (bucket_bypass_threshold_oneway)
  );


  //------------------------------
  // markov one-way thresholds
  //------------------------------
  assign markov_hi_threshold = es_bypass_mode ? markov_hi_bypass_threshold_oneway :
         markov_hi_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_markov_hi_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (markov_hi_fips_threshold_wr),
    .value_i             (markov_hi_fips_threshold),
    .value_o             (markov_hi_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_markov_hi_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (markov_hi_bypass_threshold_wr),
    .value_i             (markov_hi_bypass_threshold),
    .value_o             (markov_hi_bypass_threshold_oneway)
  );

  assign markov_lo_threshold = es_bypass_mode ? markov_lo_bypass_threshold_oneway :
         markov_lo_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_markov_lo_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (markov_lo_fips_threshold_wr),
    .value_i             (markov_lo_fips_threshold),
    .value_o             (markov_lo_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_markov_lo_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (markov_lo_bypass_threshold_wr),
    .value_i             (markov_lo_bypass_threshold),
    .value_o             (markov_lo_bypass_threshold_oneway)
  );


  //------------------------------
  // extht one-way thresholds
  //------------------------------
  assign extht_hi_threshold = es_bypass_mode ? extht_hi_bypass_threshold_oneway :
         extht_hi_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_extht_hi_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (extht_hi_fips_threshold_wr),
    .value_i             (extht_hi_fips_threshold),
    .value_o             (extht_hi_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_extht_hi_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (extht_hi_bypass_threshold_wr),
    .value_i             (extht_hi_bypass_threshold),
    .value_o             (extht_hi_bypass_threshold_oneway)
  );


  assign extht_lo_threshold = es_bypass_mode ? extht_lo_bypass_threshold_oneway :
         extht_lo_fips_threshold_oneway;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_extht_lo_thresh_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (extht_lo_fips_threshold_wr),
    .value_i             (extht_lo_fips_threshold),
    .value_o             (extht_lo_fips_threshold_oneway)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_extht_lo_thresh_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (1'b0),
    .event_i             (extht_lo_bypass_threshold_wr),
    .value_i             (extht_lo_bypass_threshold),
    .value_o             (extht_lo_bypass_threshold_oneway)
  );



  //------------------------------
  // misc control settings
  //------------------------------

  assign event_es_health_test_failed = es_main_sm_alert;

  assign event_es_observe_fifo_ready = observe_fifo_thresh_met;

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_es_route;
  mubi4_t [1:0] mubi_es_route_fanout;
  assign mubi_es_route = mubi4_t'(reg2hw.entropy_control.es_route.q);
  assign es_route_pfe = mubi4_test_true_strict(mubi_es_route_fanout[0]);
  assign es_route_pfa = mubi4_test_invalid(mubi_es_route_fanout[1]);
  assign hw2reg.recov_alert_sts.es_route_field_alert.de = es_route_pfa;
  assign hw2reg.recov_alert_sts.es_route_field_alert.d  = es_route_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_es_route (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_es_route),
    .mubi_o(mubi_es_route_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_es_type;
  mubi4_t [1:0] mubi_es_type_fanout;
  assign mubi_es_type = mubi4_t'(reg2hw.entropy_control.es_type.q);
  assign es_type_pfe = mubi4_test_true_strict(mubi_es_type_fanout[0]);
  assign es_type_pfa = mubi4_test_invalid(mubi_es_type_fanout[1]);
  assign hw2reg.recov_alert_sts.es_type_field_alert.de = es_type_pfa;
  assign hw2reg.recov_alert_sts.es_type_field_alert.d  = es_type_pfa;

  prim_mubi4_sync #(
    .NumCopies(2),
    .AsyncOn(0)
  ) u_prim_mubi4_sync_es_type (
    .clk_i,
    .rst_ni,
    .mubi_i(mubi_es_type),
    .mubi_o(mubi_es_type_fanout)
  );

  // SEC_CM: CONFIG.MUBI
  mubi4_t mubi_thresh_scope;
  assign mubi_thresh_scope = mubi4_t'(reg2hw.conf.threshold_scope.q);
  assign threshold_scope_pfe = mubi4_test_true_strict(mubi_thresh_scope);
  assign threshold_scope_pfa = mubi4_test_invalid(mubi_thresh_scope);
  assign hw2reg.recov_alert_sts.threshold_scope_field_alert.de = threshold_scope_pfa;
  assign hw2reg.recov_alert_sts.threshold_scope_field_alert.d  = threshold_scope_pfa;

  assign es_route_to_sw = es_route_pfe;
  assign es_bypass_to_sw = es_type_pfe;
  assign threshold_scope = threshold_scope_pfe;

  assign es_bypass_mode = (!fips_enable_pfe) || (es_bypass_to_sw && es_route_to_sw);

  // send off to AST RNG for possibly faster entropy generation
  assign rng_fips_o = !es_bypass_mode;

  //--------------------------------------------
  // common health test window counter
  //--------------------------------------------

  // Window counter
  // SEC_CM: CTR.REDUN
  prim_count #(
    .Width(HalfRegWidth)
  ) u_prim_count_window_cntr (
    .clk_i,
    .rst_ni,
    .clr_i(!es_delayed_enable),
    .set_i(health_test_done_pulse),
    .set_cnt_i(HalfRegWidth'(0)),
    .incr_en_i(health_test_esbus_vld),
    .decr_en_i(1'b0),
    .step_i(HalfRegWidth'(1)),
    .cnt_o(window_cntr),
    .cnt_next_o(),
    .err_o(window_cntr_err)
  );

  // Window wrap condition
  assign health_test_done_pulse = (window_cntr >= health_test_window);

  // Summary of counter errors
  assign es_cntr_err =
         (window_cntr_err ||
          repcnt_cntr_err ||
          repcnts_cntr_err ||
          adaptp_cntr_err ||
          bucket_cntr_err ||
          markov_cntr_err ||
          repcnt_fails_cntr_err ||
          repcnt_alert_cntr_err ||
          repcnts_fails_cntr_err ||
          repcnts_alert_cntr_err ||
          adaptp_hi_fails_cntr_err ||
          adaptp_lo_fails_cntr_err ||
          adaptp_hi_alert_cntr_err ||
          adaptp_lo_alert_cntr_err ||
          bucket_fails_cntr_err ||
          bucket_alert_cntr_err ||
          markov_hi_fails_cntr_err ||
          markov_lo_fails_cntr_err ||
          markov_hi_alert_cntr_err ||
          markov_lo_alert_cntr_err ||
          extht_hi_fails_cntr_err ||
          extht_lo_fails_cntr_err ||
          extht_hi_alert_cntr_err ||
          extht_lo_alert_cntr_err ||
          any_fails_cntr_err ||
          sha3_count_error);

  //--------------------------------------------
  // repetitive count test
  //--------------------------------------------

  // SEC_CM: RNG.BKGN_CHK
  entropy_src_repcnt_ht #(
    .RegWidth(HalfRegWidth),
    .RngBusWidth(RngBusWidth)
  ) u_entropy_src_repcnt_ht (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .entropy_bit_i       (health_test_esbus),
    .entropy_bit_vld_i   (health_test_esbus_vld),
    .clear_i             (health_test_clr),
    .active_i            (repcnt_active),
    .thresh_i            (repcnt_threshold),
    .test_cnt_o          (repcnt_event_cnt),
    .test_fail_pulse_o   (repcnt_fail_pulse),
    .count_err_o         (repcnt_cntr_err)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_repcnt_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (!es_bypass_mode),
    .value_i             (repcnt_event_cnt),
    .value_o             (repcnt_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_repcnt_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (es_bypass_mode),
    .value_i             (repcnt_event_cnt),
    .value_o             (repcnt_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_repcnt (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (repcnt_fail_pulse),
    .value_o             (repcnt_total_fails),
    .err_o               (repcnt_fails_cntr_err)
  );

  assign hw2reg.repcnt_hi_watermarks.fips_watermark.d = repcnt_event_hwm_fips;
  assign hw2reg.repcnt_hi_watermarks.bypass_watermark.d = repcnt_event_hwm_bypass;
  assign hw2reg.repcnt_total_fails.d = repcnt_total_fails;

  //--------------------------------------------
  // repetitive count symbol test
  //--------------------------------------------

  // SEC_CM: RNG.BKGN_CHK
  entropy_src_repcnts_ht #(
    .RegWidth(HalfRegWidth),
    .RngBusWidth(RngBusWidth)
  ) u_entropy_src_repcnts_ht (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .entropy_bit_i       (health_test_esbus),
    .entropy_bit_vld_i   (health_test_esbus_vld),
    .clear_i             (health_test_clr),
    .active_i            (repcnts_active),
    .thresh_i            (repcnts_threshold),
    .test_cnt_o          (repcnts_event_cnt),
    .test_fail_pulse_o   (repcnts_fail_pulse),
    .count_err_o         (repcnts_cntr_err)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_repcnts_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (!es_bypass_mode),
    .value_i             (repcnts_event_cnt),
    .value_o             (repcnts_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_repcnts_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (es_bypass_mode),
    .value_i             (repcnts_event_cnt),
    .value_o             (repcnts_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_repcnts (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (repcnts_fail_pulse),
    .value_o             (repcnts_total_fails),
    .err_o               (repcnts_fails_cntr_err)
  );

  assign hw2reg.repcnts_hi_watermarks.fips_watermark.d = repcnts_event_hwm_fips;
  assign hw2reg.repcnts_hi_watermarks.bypass_watermark.d = repcnts_event_hwm_bypass;
  assign hw2reg.repcnts_total_fails.d = repcnts_total_fails;

  //--------------------------------------------
  // adaptive proportion test
  //--------------------------------------------

  // SEC_CM: RNG.BKGN_CHK
  entropy_src_adaptp_ht #(
    .RegWidth(HalfRegWidth),
    .RngBusWidth(RngBusWidth)
  ) u_entropy_src_adaptp_ht (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .entropy_bit_i       (health_test_esbus),
    .entropy_bit_vld_i   (health_test_esbus_vld),
    .clear_i             (health_test_clr),
    .active_i            (adaptp_active),
    .thresh_hi_i         (adaptp_hi_threshold),
    .thresh_lo_i         (adaptp_lo_threshold),
    .window_wrap_pulse_i (health_test_done_pulse),
    .threshold_scope_i   (threshold_scope),
    .test_cnt_hi_o       (adaptp_hi_event_cnt),
    .test_cnt_lo_o       (adaptp_lo_event_cnt),
    .test_fail_hi_pulse_o(adaptp_hi_fail_pulse),
    .test_fail_lo_pulse_o(adaptp_lo_fail_pulse),
    .count_err_o         (adaptp_cntr_err)
  );


  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_adaptp_hi_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && !es_bypass_mode),
    .value_i             (adaptp_hi_event_cnt),
    .value_o             (adaptp_hi_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_adaptp_hi_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && es_bypass_mode),
    .value_i             (adaptp_hi_event_cnt),
    .value_o             (adaptp_hi_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_adaptp_hi (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (adaptp_hi_fail_pulse),
    .value_o             (adaptp_hi_total_fails),
    .err_o               (adaptp_hi_fails_cntr_err)
  );


  assign hw2reg.adaptp_hi_watermarks.fips_watermark.d = adaptp_hi_event_hwm_fips;
  assign hw2reg.adaptp_hi_watermarks.bypass_watermark.d = adaptp_hi_event_hwm_bypass;
  assign hw2reg.adaptp_hi_total_fails.d = adaptp_hi_total_fails;


  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_adaptp_lo_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && !es_bypass_mode),
    .value_i             (adaptp_lo_event_cnt),
    .value_o             (adaptp_lo_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_adaptp_lo_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && es_bypass_mode),
    .value_i             (adaptp_lo_event_cnt),
    .value_o             (adaptp_lo_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_adaptp_lo (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (adaptp_lo_fail_pulse),
    .value_o             (adaptp_lo_total_fails),
    .err_o               (adaptp_lo_fails_cntr_err)
  );

  assign hw2reg.adaptp_lo_watermarks.fips_watermark.d = adaptp_lo_event_hwm_fips;
  assign hw2reg.adaptp_lo_watermarks.bypass_watermark.d = adaptp_lo_event_hwm_bypass;
  assign hw2reg.adaptp_lo_total_fails.d = adaptp_lo_total_fails;


  //--------------------------------------------
  // bucket test
  //--------------------------------------------

  // SEC_CM: RNG.BKGN_CHK
  entropy_src_bucket_ht #(
    .RegWidth(HalfRegWidth),
    .RngBusWidth(RngBusWidth)
  ) u_entropy_src_bucket_ht (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .entropy_bit_i       (health_test_esbus),
    .entropy_bit_vld_i   (health_test_esbus_vld),
    .clear_i             (health_test_clr),
    .active_i            (bucket_active),
    .thresh_i            (bucket_threshold),
    .window_wrap_pulse_i (health_test_done_pulse),
    .test_cnt_o          (bucket_event_cnt),
    .test_fail_pulse_o   (bucket_fail_pulse),
    .count_err_o         (bucket_cntr_err)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_bucket_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && !es_bypass_mode),
    .value_i             (bucket_event_cnt),
    .value_o             (bucket_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_bucket_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && es_bypass_mode),
    .value_i             (bucket_event_cnt),
    .value_o             (bucket_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_bucket (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (bucket_fail_pulse),
    .value_o             (bucket_total_fails),
    .err_o               (bucket_fails_cntr_err)
  );

  assign hw2reg.bucket_hi_watermarks.fips_watermark.d = bucket_event_hwm_fips;
  assign hw2reg.bucket_hi_watermarks.bypass_watermark.d = bucket_event_hwm_bypass;
  assign hw2reg.bucket_total_fails.d = bucket_total_fails;


  //--------------------------------------------
  // Markov test
  //--------------------------------------------

  // SEC_CM: RNG.BKGN_CHK
  entropy_src_markov_ht #(
    .RegWidth(HalfRegWidth),
    .RngBusWidth(RngBusWidth)
  ) u_entropy_src_markov_ht (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .entropy_bit_i       (health_test_esbus),
    .entropy_bit_vld_i   (health_test_esbus_vld),
    .clear_i             (health_test_clr),
    .active_i            (markov_active),
    .thresh_hi_i         (markov_hi_threshold),
    .thresh_lo_i         (markov_lo_threshold),
    .window_wrap_pulse_i (health_test_done_pulse),
    .threshold_scope_i   (threshold_scope),
    .test_cnt_hi_o       (markov_hi_event_cnt),
    .test_cnt_lo_o       (markov_lo_event_cnt),
    .test_fail_hi_pulse_o (markov_hi_fail_pulse),
    .test_fail_lo_pulse_o (markov_lo_fail_pulse),
    .count_err_o         (markov_cntr_err)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_markov_hi_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && !es_bypass_mode),
    .value_i             (markov_hi_event_cnt),
    .value_o             (markov_hi_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_markov_hi_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && es_bypass_mode),
    .value_i             (markov_hi_event_cnt),
    .value_o             (markov_hi_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_markov_hi (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (markov_hi_fail_pulse),
    .value_o             (markov_hi_total_fails),
    .err_o               (markov_hi_fails_cntr_err)
  );

  assign hw2reg.markov_hi_watermarks.fips_watermark.d = markov_hi_event_hwm_fips;
  assign hw2reg.markov_hi_watermarks.bypass_watermark.d = markov_hi_event_hwm_bypass;
  assign hw2reg.markov_hi_total_fails.d = markov_hi_total_fails;


  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_markov_lo_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && !es_bypass_mode),
    .value_i             (markov_lo_event_cnt),
    .value_o             (markov_lo_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_markov_lo_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (health_test_done_pulse && es_bypass_mode),
    .value_i             (markov_lo_event_cnt),
    .value_o             (markov_lo_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_markov_lo (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (markov_lo_fail_pulse),
    .value_o             (markov_lo_total_fails),
    .err_o               (markov_lo_fails_cntr_err)
  );

  assign hw2reg.markov_lo_watermarks.fips_watermark.d = markov_lo_event_hwm_fips;
  assign hw2reg.markov_lo_watermarks.bypass_watermark.d = markov_lo_event_hwm_bypass;
  assign hw2reg.markov_lo_total_fails.d = markov_lo_total_fails;


  //--------------------------------------------
  // External health test
  //--------------------------------------------

  // set outputs to external health test
  assign entropy_src_xht_o.entropy_bit = health_test_esbus;
  assign entropy_src_xht_o.entropy_bit_valid = health_test_esbus_vld;
  assign entropy_src_xht_o.clear = health_test_clr;
  assign entropy_src_xht_o.active = extht_active;
  assign entropy_src_xht_o.thresh_hi = extht_hi_threshold;
  assign entropy_src_xht_o.thresh_lo = extht_lo_threshold;
  assign entropy_src_xht_o.window_wrap_pulse = health_test_done_pulse;
  assign entropy_src_xht_o.health_test_window = health_test_window;
  assign entropy_src_xht_o.threshold_scope = threshold_scope;
  // get inputs from external health test
  assign extht_event_cnt_hi = entropy_src_xht_i.test_cnt_hi;
  assign extht_event_cnt_lo = entropy_src_xht_i.test_cnt_lo;
  assign extht_hi_fail_pulse = entropy_src_xht_i.test_fail_hi_pulse;
  assign extht_lo_fail_pulse = entropy_src_xht_i.test_fail_lo_pulse;
  assign extht_cont_test = entropy_src_xht_i.continuous_test;

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_extht_hi_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             ((extht_cont_test || health_test_done_pulse) && !es_bypass_mode),
    .value_i             (extht_event_cnt_hi),
    .value_o             (extht_hi_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(1)
  ) u_entropy_src_watermark_reg_extht_hi_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             ((extht_cont_test || health_test_done_pulse) && es_bypass_mode),
    .value_i             (extht_event_cnt_hi),
    .value_o             (extht_hi_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_extht_hi (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (extht_hi_fail_pulse),
    .value_o             (extht_hi_total_fails),
    .err_o               (extht_hi_fails_cntr_err)
  );


  assign hw2reg.extht_hi_watermarks.fips_watermark.d = extht_hi_event_hwm_fips;
  assign hw2reg.extht_hi_watermarks.bypass_watermark.d = extht_hi_event_hwm_bypass;
  assign hw2reg.extht_hi_total_fails.d = extht_hi_total_fails;


  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_extht_lo_fips (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             ((extht_cont_test || health_test_done_pulse) && !es_bypass_mode),
    .value_i             (extht_event_cnt_lo),
    .value_o             (extht_lo_event_hwm_fips)
  );

  entropy_src_watermark_reg #(
    .RegWidth(HalfRegWidth),
    .HighWatermark(0)
  ) u_entropy_src_watermark_reg_extht_lo_bypass (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             ((extht_cont_test || health_test_done_pulse) && es_bypass_mode),
    .value_i             (extht_event_cnt_lo),
    .value_o             (extht_lo_event_hwm_bypass)
  );

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(FullRegWidth)
  ) u_entropy_src_cntr_reg_extht_lo (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (health_test_clr),
    .event_i             (extht_lo_fail_pulse),
    .value_o             (extht_lo_total_fails),
    .err_o               (extht_lo_fails_cntr_err)
  );

  assign hw2reg.extht_lo_watermarks.fips_watermark.d = extht_lo_event_hwm_fips;
  assign hw2reg.extht_lo_watermarks.bypass_watermark.d = extht_lo_event_hwm_bypass;
  assign hw2reg.extht_lo_total_fails.d = extht_lo_total_fails;


  //--------------------------------------------
  // summary and alert registers
  //--------------------------------------------

  assign alert_cntrs_clr = health_test_clr || rst_alert_cntr;

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(HalfRegWidth)
  ) u_entropy_src_cntr_reg_any_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (any_fail_pulse),
    .value_o             (any_fail_count),
    .err_o               (any_fails_cntr_err)
  );

  assign any_fail_pulse =
         repcnt_fail_pulse ||
         repcnts_fail_pulse ||
         adaptp_hi_fail_pulse || adaptp_lo_fail_pulse ||
         bucket_fail_pulse ||
         markov_hi_fail_pulse || markov_lo_fail_pulse ||
         extht_hi_fail_pulse || extht_lo_fail_pulse;

  assign ht_failed_d =
         (!es_enable_fo[6]) ? 1'b0 :
         ht_done_pulse_q ? 1'b0 :
         any_fail_pulse ? 1'b1 :
         ht_failed_q;


  // delay health pulse so that main_sm will
  // get the correct threshold value comparisons
  assign ht_done_pulse_d = health_test_done_pulse;

  assign hw2reg.alert_summary_fail_counts.d = any_fail_count;

  // signal an alert
  // SEC_CM: CONFIG.REDUN
  assign alert_threshold = reg2hw.alert_threshold.alert_threshold.q;
  assign alert_threshold_inv = reg2hw.alert_threshold.alert_threshold_inv.q;
  assign es_thresh_cfg_alert = (~alert_threshold_inv != alert_threshold);

  assign alert_threshold_fail =
         ((any_fail_count >= ~alert_threshold_inv) && (~alert_threshold_inv != '0)) ||
         (any_fail_count >= alert_threshold) && (alert_threshold != '0);


  prim_edge_detector #(
    .Width(1),
    .ResetValue(0),
    .EnSync(0)
  ) u_prim_edge_detector_recov_alert (
    .clk_i,
    .rst_ni,
    .d_i(recov_alert_state),
    .q_sync_o(),
    .q_posedge_pulse_o(recov_alert_o),
    .q_negedge_pulse_o()
  );

  assign recov_alert_state =
         es_enable_pfa ||
         fips_enable_pfa ||
         entropy_data_reg_en_pfa ||
         threshold_scope_pfa ||
         rng_bit_enable_pfa ||
         fw_ov_mode_pfa ||
         fw_ov_entropy_insert_pfa ||
         fw_ov_sha3_start_pfa ||
         es_route_pfa ||
         es_type_pfa ||
         es_main_sm_alert ||
         es_bus_cmp_alert ||
         es_thresh_cfg_alert ||
         es_fw_ov_wr_alert ||
         es_fw_ov_disable_alert;

  assign hw2reg.recov_alert_sts.es_main_sm_alert.de = es_main_sm_alert;
  assign hw2reg.recov_alert_sts.es_main_sm_alert.d  = es_main_sm_alert;

  assign hw2reg.recov_alert_sts.es_bus_cmp_alert.de = es_bus_cmp_alert;
  assign hw2reg.recov_alert_sts.es_bus_cmp_alert.d  = es_bus_cmp_alert;

  assign hw2reg.recov_alert_sts.es_thresh_cfg_alert.de = es_thresh_cfg_alert;
  assign hw2reg.recov_alert_sts.es_thresh_cfg_alert.d  = es_thresh_cfg_alert;

  assign hw2reg.recov_alert_sts.es_fw_ov_wr_alert.de = es_fw_ov_wr_alert;
  assign hw2reg.recov_alert_sts.es_fw_ov_wr_alert.d  = es_fw_ov_wr_alert;

  assign hw2reg.recov_alert_sts.es_fw_ov_disable_alert.de = es_fw_ov_disable_alert;
  assign hw2reg.recov_alert_sts.es_fw_ov_disable_alert.d  = es_fw_ov_disable_alert;

  // repcnt fail counter
  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_repcnt_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (repcnt_fail_pulse),
    .value_o             (repcnt_fail_count),
    .err_o               (repcnt_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.repcnt_fail_count.d = repcnt_fail_count;

  // repcnts fail counter
  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_repcnts_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (repcnts_fail_pulse),
    .value_o             (repcnts_fail_count),
    .err_o               (repcnts_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.repcnts_fail_count.d = repcnts_fail_count;

  // adaptp fail counter hi and lo
  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_adaptp_hi_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (adaptp_hi_fail_pulse),
    .value_o             (adaptp_hi_fail_count),
    .err_o               (adaptp_hi_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.adaptp_hi_fail_count.d = adaptp_hi_fail_count;

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_adaptp_lo_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (adaptp_lo_fail_pulse),
    .value_o             (adaptp_lo_fail_count),
    .err_o               (adaptp_lo_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.adaptp_lo_fail_count.d = adaptp_lo_fail_count;

  // bucket fail counter
  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_bucket_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (bucket_fail_pulse),
    .value_o             (bucket_fail_count),
    .err_o               (bucket_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.bucket_fail_count.d = bucket_fail_count;


  // markov fail counter hi and lo
  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_markov_hi_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (markov_hi_fail_pulse),
    .value_o             (markov_hi_fail_count),
    .err_o               (markov_hi_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.markov_hi_fail_count.d = markov_hi_fail_count;

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_markov_lo_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (markov_lo_fail_pulse),
    .value_o             (markov_lo_fail_count),
    .err_o               (markov_lo_alert_cntr_err)
  );

  assign hw2reg.alert_fail_counts.markov_lo_fail_count.d = markov_lo_fail_count;

  // extht fail counter hi and lo
  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_extht_hi_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (extht_hi_fail_pulse),
    .value_o             (extht_hi_fail_count),
    .err_o               (extht_hi_alert_cntr_err)
  );

  assign hw2reg.extht_fail_counts.extht_hi_fail_count.d = extht_hi_fail_count;

  // SEC_CM: CTR.REDUN
  entropy_src_cntr_reg #(
    .RegWidth(EighthRegWidth)
  ) u_entropy_src_cntr_reg_extht_lo_alert_fails (
    .clk_i               (clk_i),
    .rst_ni              (rst_ni),
    .clear_i             (alert_cntrs_clr),
    .event_i             (extht_lo_fail_pulse),
    .value_o             (extht_lo_fail_count),
    .err_o               (extht_lo_alert_cntr_err)
  );

  assign hw2reg.extht_fail_counts.extht_lo_fail_count.d = extht_lo_fail_count;


  //--------------------------------------------
  // pack tested entropy into 32 bit packer
  //--------------------------------------------

  prim_packer_fifo #(
    .InW(RngBusWidth),
    .OutW(PostHTWidth),
    .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_postht (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (pfifo_postht_clr),
    .wvalid_i   (pfifo_postht_push),
    .wdata_i    (pfifo_postht_wdata),
    .wready_o   (pfifo_postht_not_full),
    .rvalid_o   (pfifo_postht_not_empty),
    .rdata_o    (pfifo_postht_rdata),
    .rready_i   (pfifo_postht_pop),
    .depth_o    ()
  );

  assign pfifo_postht_push = rng_bit_en ? pfifo_esbit_not_empty :
                             sfifo_esrng_not_empty;

  assign pfifo_postht_wdata = rng_bit_en ? pfifo_esbit_rdata :
                              sfifo_esrng_rdata;

  // For verification purposes, let post-disable data continue through to the SHA engine if it has
  // made it past the health checks, when in standard (non-fw_ov) mode.  This allows scoreboards
  // to use the same data set for computing both the SHA engine outputs and the health-check stats.
  //
  // In fw_ov mode it is preferable (from a verification standpoint) to clear all FIFOs whenever
  // disabled. Given the lack of handshaking on the fw_ov register path, this is easier to predict.
  // Also, there is no association between SHA data and health test windows in FW_OV mode, so there
  // is no benefit in this mode to clearing the SHA FIFOs at the same time we clear the HT
  // statistics.

  assign pfifo_postht_clr = fw_ov_mode_entropy_insert ? !es_enable_fo[7] : !es_delayed_enable;

  // In firmware override mode with extract & insert enabled, post-health test entropy bits can
  // only move into the observe FIFO. Once the observe FIFO is full, post-health test entropy is
  // just discarded.
  assign pfifo_postht_pop = fw_ov_mode_entropy_insert ? pfifo_postht_not_empty :
                            // In firmware override mode (observe only) or during normal
                            // operation, post-health test entropy bits continue to flow
                            // through the hardware pipeline.
                            es_bypass_mode ? pfifo_bypass_push :
                            pfifo_precon_push & pfifo_precon_not_full;


  //--------------------------------------------
  // store entropy into a 64 entry deep FIFO
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(ObserveFifoWidth),
    .Pass(0),
    .Depth(ObserveFifoDepth)
  ) u_prim_fifo_sync_observe (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (sfifo_observe_clr),
    .wvalid_i   (sfifo_observe_push),
    .wdata_i    (sfifo_observe_wdata),
    .wready_o   (),
    .rvalid_o   (sfifo_observe_not_empty),
    .rdata_o    (sfifo_observe_rdata),
    .rready_i   (sfifo_observe_pop),
    .full_o     (sfifo_observe_full),
    .depth_o    (sfifo_observe_depth),
    .err_o      ()
  );

  // The Observe fifo is intended to hold kilobits of contiguous data, yet still gracefully
  // drop data when full.  This flop gates the observe fifo. If it ever overflows, no new data is
  // allowed until it is empty.  Thus if the rate of CSR uptake almost matches the RNG data rate
  // the FIFO avoids unnecessary segmentation, and guarantees that the remaining RNG data is as
  // contiguous as possible.
  logic sfifo_observe_gate_d, sfifo_observe_gate_q;

  assign sfifo_observe_gate_d = (sfifo_observe_push && sfifo_observe_full) ? 1'b0 :
                                !sfifo_observe_not_empty                   ? 1'b1 :
                                sfifo_observe_gate_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      sfifo_observe_gate_q <= 1'b1;
    end else begin
      sfifo_observe_gate_q <= sfifo_observe_gate_d;
    end
  end

  assign hw2reg.fw_ov_rd_fifo_overflow.d  = (pfifo_postht_pop && sfifo_observe_full);
  assign hw2reg.fw_ov_rd_fifo_overflow.de = 1'b1;

  assign observe_fifo_thresh_met = fw_ov_mode && (observe_fifo_thresh != '0) &&
         (observe_fifo_thresh <= sfifo_observe_depth) && es_enable_fo[8];

  assign hw2reg.observe_fifo_depth.d = sfifo_observe_depth;

  // fifo controls
  assign sfifo_observe_push = fw_ov_mode && pfifo_postht_pop && !sfifo_observe_full &&
                              (sfifo_observe_gate_q || !sfifo_observe_not_empty);

  assign sfifo_observe_clr  = ~es_enable_fo[9];

  assign sfifo_observe_wdata = pfifo_postht_rdata;

  assign sfifo_observe_pop =
         (fw_ov_mode && fw_ov_fifo_rd_pulse);

  // fifo err
  assign sfifo_observe_err =
         {(sfifo_observe_push && sfifo_observe_full),
         (sfifo_observe_pop && !sfifo_observe_not_empty),
         (sfifo_observe_full && !sfifo_observe_not_empty)};


  //--------------------------------------------
  // pack entropy into 64 bit packer
  //--------------------------------------------

  prim_packer_fifo #(
    .InW(ObserveFifoWidth),
    .OutW(PreCondWidth),
    .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_precon (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (pfifo_precon_clr),
    .wvalid_i   (pfifo_precon_push),
    .wdata_i    (pfifo_precon_wdata),
    .wready_o   (pfifo_precon_not_full),
    .rvalid_o   (pfifo_precon_not_empty),
    .rdata_o    (pfifo_precon_rdata),
    .rready_i   (pfifo_precon_pop),
    .depth_o    ()
  );

  // When bypassing the hardware conditioning - due to a) disabling FIPS mode or b) routing entropy
  // to the ENTROPY_DATA register (ES_ROUTE) and bypassing the conditioner (ES_TYPE) - nothing is
  // going into the conditioner.
  assign pfifo_precon_push = es_bypass_mode ? 1'b0 :
                             // In firmware override mode with extract & insert enabled, only bits
                             // inserted by firmware continue down the pipeline.
                             fw_ov_mode_entropy_insert ? fw_ov_fifo_wr_pulse :
                             // Otherwise post-health test entropy bits continue to flow
                             // downstream. This includes observe-only firmware override mode.
                             pfifo_postht_not_empty;

  assign pfifo_precon_wdata = fw_ov_mode_entropy_insert ? fw_ov_wr_data :
                              pfifo_postht_rdata;

  // For verification purposes, let post-disable data continue through to the SHA engine if it has
  // made it past the health checks, when in standard (non-fw_ov) mode.  This allows scoreboards
  // to use the same data set for computing both the SHA engine outputs and the health-check stats.
  //
  // In fw_ov mode it is preferable (from a verification standpoint) to clear all FIFOs whenever
  // disabled. Given the lack of handshaking on the fw_ov register path, this is easier to predict.
  // Also, there is no association between SHA data and health test windows in FW_OV mode, so there
  // is no benefit in this mode to clearing the SHA FIFOs at the same time we clear the HT
  // statistics.
  //
  // Corner case: Even in FW_OV mode, if a full SHA word is ready as the disable comes in,
  // let it stay in the FIFO until the SHA engine has picked it up, as verification has no way
  // of knowing if a word will get stalled by SHA backpressure.  This is not a problem however
  // as the reset is only important for clearing 32-bit half-SHA-words.
  assign pfifo_precon_clr = fw_ov_mode_entropy_insert ?
                            ~es_enable_fo[10] & ~pfifo_precon_not_empty :
                            ~es_delayed_enable & ~pfifo_precon_not_empty;

  assign pfifo_precon_pop = (pfifo_cond_push && sha3_msgfifo_ready);

  assign es_fw_ov_wr_alert = fw_ov_mode && fw_ov_mode_entropy_insert &&
         fw_ov_fifo_wr_pulse && fw_ov_wr_fifo_full;

  assign es_fw_ov_disable_alert = fw_ov_mode && fw_ov_mode_entropy_insert &&
         !es_bypass_mode && fw_ov_sha3_disable_pulse && fw_ov_wr_fifo_full;

  //--------------------------------------------
  // entropy conditioner
  //--------------------------------------------
  // This block will take in raw entropy from the noise source block
  // and compress it such that a perfect entropy source is created
  // This block will take in 2048 (by default setting) bits to create 384 bits.

  // Note on backpressure from the SHA block:
  // If we use the full sha3_msgfifo_ready signal, we create a combinational logic
  // loop.  However, the SHA3 seems to have a hiccup by which it some times
  // asserts ready even though it is processing data, so we mask our push
  // signal with our (flop-based) sha3_msg_rdy_mask
  assign pfifo_cond_push  = pfifo_precon_not_empty && !es_bypass_mode && sha3_msg_rdy_mask;

  assign pfifo_cond_wdata = pfifo_precon_rdata;

  assign msg_data[0] = pfifo_cond_wdata;

  // The SHA3 block cannot take messages except between the
  // start and cs_aes_req pulses
  assign sha3_msg_end        = cs_aes_halt_req;

  assign sha3_msg_rdy_mask_d = sha3_start ? 1'b1 :
                               sha3_msg_end ? 1'b0 :
                               sha3_msg_rdy_mask_q;

  assign sha3_msg_rdy_mask = sha3_msg_rdy_mask_q & ~sha3_msg_end &
                             ~cs_aes_halt_req;

  assign pfifo_cond_rdata = sha3_state[0][SeedLen-1:0];
  assign pfifo_cond_not_empty = sha3_state_vld;
  assign sha3_msgfifo_ready = sha3_msg_rdy & sha3_msg_rdy_mask;

  // SHA3 hashing engine
  sha3 #(
    .EnMasking (Sha3EnMasking)
  ) u_sha3 (
    .clk_i,
    .rst_ni,

    // MSG_FIFO interface
    .msg_valid_i (pfifo_cond_push),
    .msg_data_i  (msg_data),
    .msg_strb_i  ({8{pfifo_cond_push}}),
    .msg_ready_o (sha3_msg_rdy),

    // Entropy interface - not using
    .rand_valid_i    (1'b0),
    .rand_early_i    (1'b0),
    .rand_data_i     ('0),
    .rand_aux_i      ('0),
    .rand_consumed_o (),

    // N, S: Used in cSHAKE mode
    .ns_data_i       ('0), // ns_prefix),

    // Configurations
    .mode_i     (sha3_pkg::Sha3), // Use SHA3 mode
    .strength_i (sha3_pkg::L384), // Use keccak_strength_e of L384

    // Controls (CMD register)
    .start_i    (sha3_start       ),
    .process_i  (sha3_process     ),
    .run_i      (1'b0             ), // For software application
    .done_i     (sha3_done        ),

    // LC escalation
    .lc_escalate_en_i (lc_ctrl_pkg::Off),

    .absorbed_o (sha3_absorbed),
    .squeezing_o (sha3_squeezing),

    .block_processed_o (sha3_block_processed),

    .sha3_fsm_o (sha3_fsm),

    .state_valid_o (sha3_state_vld),
    .state_o       (sha3_state),

    .error_o (sha3_err),
    .sparse_fsm_error_o (sha3_state_error),
    .count_error_o  (sha3_count_error),
    .keccak_storage_rst_error_o (sha3_rst_storage_err)
  );

  //--------------------------------------------
  // bypass SHA conditioner path
  //--------------------------------------------

  prim_packer_fifo #(
     .InW(PostHTWidth),
     .OutW(SeedLen),
     .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_bypass (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (pfifo_bypass_clr),
    .wvalid_i   (pfifo_bypass_push),
    .wdata_i    (pfifo_bypass_wdata),
    .wready_o   (pfifo_bypass_not_full),
    .rvalid_o   (pfifo_bypass_not_empty),
    .rdata_o    (pfifo_bypass_rdata),
    .rready_i   (pfifo_bypass_pop),
    .depth_o    ()
  );

  // Unless the hardware conditioning is bypassed - due to a) disabling FIPS mode or b) routing
  // entropy to the ENTROPY_DATA register (ES_ROUTE) and bypassing the conditioner (ES_TYPE) -
  // nothing is going into the bypass FIFO.
  assign pfifo_bypass_push = !es_bypass_mode ? 1'b0 :
                             // In firmware override mode with extract & insert enabled, only bits
                             // inserted by firmware continue down the pipeline
                             fw_ov_mode_entropy_insert ? fw_ov_fifo_wr_pulse :
                             // Otherwise post-health test entropy bits continue to flow
                             // downstream. This includes observe-only firmware override mode.
                             pfifo_postht_not_empty;

  assign pfifo_bypass_wdata = fw_ov_mode_entropy_insert ? fw_ov_wr_data :
                              pfifo_postht_rdata;

  assign pfifo_bypass_clr = !es_enable_fo[11];

  // Corner case: If the main state machine encounters an alert, drain the
  // bypass fifo, to get rid of the seeds and let the HT stats continue.
  assign pfifo_bypass_pop =
         fw_ov_mode_entropy_insert ? pfifo_bypass_not_empty :
         bypass_stage_pop;

  // mux to select between fips and bypass mode
  assign final_es_data = es_bypass_mode ? pfifo_bypass_rdata : pfifo_cond_rdata;


  //--------------------------------------------
  // state machine to coordinate fifo flow
  //--------------------------------------------

  // SEC_CM: CTR.LOCAL_ESC
  // SEC_CM: MAIN_SM.FSM.SPARSE
  entropy_src_main_sm
    u_entropy_src_main_sm (
    .clk_i                (clk_i),
    .rst_ni               (rst_ni),
    .enable_i             (main_sm_enable),
    .fw_ov_ent_insert_i   (fw_ov_mode_entropy_insert),
    .fw_ov_sha3_start_i   (fw_ov_sha3_start_pfe),
    .ht_done_pulse_i      (ht_done_pulse_q),
    .ht_fail_pulse_i      (ht_failed_q),
    .alert_thresh_fail_i  (alert_threshold_fail),
    .rst_alert_cntr_o     (rst_alert_cntr),
    .bypass_mode_i        (es_bypass_mode),
    .main_stage_rdy_i     (pfifo_cond_not_empty),
    .bypass_stage_rdy_i   (pfifo_bypass_not_empty),
    .sha3_state_vld_i     (sha3_state_vld),
    .main_stage_push_o    (main_stage_push_raw),
    .bypass_stage_pop_o   (bypass_stage_pop),
    .boot_phase_done_o    (boot_phase_done),
    .sha3_start_o         (sha3_start_raw),
    .sha3_process_o       (sha3_process),
    .sha3_done_o          (sha3_done),
    .cs_aes_halt_req_o    (cs_aes_halt_req),
    .cs_aes_halt_ack_i    (cs_aes_halt_i.cs_aes_halt_ack),
    .local_escalate_i     (es_cntr_err_sum),
    .main_sm_alert_o      (es_main_sm_alert),
    .main_sm_idle_o       (es_main_sm_idle),
    .main_sm_state_o      (es_main_sm_state),
    .main_sm_err_o        (es_main_sm_err)
  );

  // es to cs halt request to reduce power spikes
  assign cs_aes_halt_d = cs_aes_halt_req;
  assign cs_aes_halt_o.cs_aes_halt_req = cs_aes_halt_q;

  //--------------------------------------------
  // Corner case masking of main_sm inputs/outputs
  //--------------------------------------------

  // When operating in RNG mode the state machine does not respond
  // immediately to disable requests if it processing the SHA output
  // (here indicated by the cs_aes_halt_req handshake).  The SHA engine
  // will continue to process even if the module is disabled.  These seeds
  // that continue to process after the disable signal are referred to as
  // stale.
  //
  // If the SHA processing were instantaneous, stale seeds would be discarded
  // when the esfinal fifo was cleard on diable.  Though since processing
  // can push through a disable pulse, stale seeds need to be identified,
  // and held back from the esfinal FIFO.
  //
  // There is at most one seed processing at a time so, we simply need to
  // detect when a stale seed has commenced processing, and mask the following
  // main_stage_push signal.

  assign stale_seed_processing = ~es_bypass_mode & ~fw_ov_mode_entropy_insert &
                                 cs_aes_halt_req & ~es_enable_fo[12];
  assign sha3_flush_d = stale_seed_processing ? 1'b1 :
                        main_stage_push_raw ? 1'b0 :
                        sha3_flush_q;

  // If the user incorrectly disables the fw_ov SHA3 processing while
  // data is in the pipeline, it can potentially scramble two outputs.
  // Thus in addition to triggering a recoverable alert, we mark the
  // following _two_ outputs as corrupted and to not let them in the
  // esfinal FIFO
  assign fw_ov_corrupted_d = es_fw_ov_disable_alert ? 2'b11 :
                             !es_bypass_mode && main_stage_push_raw ? {1'b0, fw_ov_corrupted_q[1]} :
                             fw_ov_corrupted_q;

  assign fw_ov_corrupted = (|fw_ov_corrupted_q) & !es_bypass_mode;


  assign main_stage_push = main_stage_push_raw & !sha3_flush_q & !fw_ov_corrupted;

  // Use the delayed enable signal to keep the Main SM enabled while Data is in flight, and
  // to make sure it receives a delayed disable pulse after finishing any final SHA processing
  // commands
  assign main_sm_enable = es_delayed_enable;

  // The main SM can also generate redundant start pulses. After data can be pushed into SHA,
  // the SM can be disabled leaving entropy in the SHA sponge.  This is fine, but the SM will
  // have no recollection of this previous start pulse.  We track redundant start pulses
  // outside the SM and suppress them as needed.
  assign sha3_start_mask_d = sha3_start_raw ? 1'b1 :
                             sha3_process   ? 1'b0 :
                             sha3_start_mask_q;
  assign sha3_start = sha3_start_raw & ~sha3_start_mask_q;

  //--------------------------------------------
  // send processed entropy to final fifo
  //--------------------------------------------

  prim_fifo_sync #(
    .Width(1+SeedLen),
    .Pass(0),
    .Depth(EsFifoDepth),
    .OutputZeroIfEmpty(1'b0)
  ) u_prim_fifo_sync_esfinal (
    .clk_i          (clk_i),
    .rst_ni         (rst_ni),
    .clr_i          (sfifo_esfinal_clr),
    .wvalid_i       (sfifo_esfinal_push),
    .wready_o       (sfifo_esfinal_not_full),
    .wdata_i        (sfifo_esfinal_wdata),
    .rvalid_o       (sfifo_esfinal_not_empty),
    .rready_i       (sfifo_esfinal_pop),
    .rdata_o        (sfifo_esfinal_rdata),
    .full_o         (sfifo_esfinal_full),
    .depth_o        (sfifo_esfinal_depth),
    .err_o          ()
  );

  assign fips_compliance = !es_bypass_mode && es_enable_fo[13] && !rng_bit_en;

  // fifo controls
  assign sfifo_esfinal_push_enable =
         fw_ov_mode_entropy_insert && es_bypass_mode ? pfifo_bypass_not_empty :
         main_stage_push;

  assign sfifo_esfinal_push = sfifo_esfinal_not_full && sfifo_esfinal_push_enable;
  assign sfifo_esfinal_clr  = !es_enable_fo[14];
  assign sfifo_esfinal_wdata = {fips_compliance,final_es_data};
  assign sfifo_esfinal_pop = es_route_to_sw ? pfifo_swread_push :
         es_hw_if_fifo_pop;
  assign {esfinal_fips_flag,esfinal_data} = sfifo_esfinal_rdata;

  // fifo err
  // Note: for prim_fifo_sync is not an error to push to a fifo that is full.  In fact, the
  // backpressure mechanism applied to the previous FIFO counts on this.
  assign sfifo_esfinal_err =
         {1'b0,
          (sfifo_esfinal_pop && !sfifo_esfinal_not_empty),
          (sfifo_esfinal_full && !sfifo_esfinal_not_empty)};

  // drive out hw interface
  assign es_hw_if_req = entropy_src_hw_if_i.es_req;
  assign entropy_src_hw_if_o.es_ack = es_hw_if_ack;
  assign entropy_src_hw_if_o.es_bits = esfinal_data;
  assign entropy_src_hw_if_o.es_fips = esfinal_fips_flag;

  // SEC_CM: ACK_SM.FSM.SPARSE
  entropy_src_ack_sm u_entropy_src_ack_sm (
    .clk_i            (clk_i),
    .rst_ni           (rst_ni),
    .enable_i         (es_enable_fo[15]),
    .req_i            (es_hw_if_req),
    .ack_o            (es_hw_if_ack),
    .fifo_not_empty_i (sfifo_esfinal_not_empty && !es_route_to_sw),
    .local_escalate_i (es_cntr_err),
    .fifo_pop_o       (es_hw_if_fifo_pop),
    .ack_sm_err_o     (es_ack_sm_err)
  );

  //--------------------------------------------
  // data path integrity check
  // - a countermeasure to detect entropy bus tampering attempts
  // - checks to make sure repeated data sets off
  //   an alert for sw to handle
  //--------------------------------------------

  // SEC_CM: ESFINAL_RDATA.BUS.CONSISTENCY

  // capture a copy of the entropy data
  assign es_rdata_capt_vld = (sfifo_esfinal_pop && sfifo_esfinal_not_empty);

  assign es_rdata_capt_d = es_rdata_capt_vld ? sfifo_esfinal_rdata[63:0] : es_rdata_capt_q;

  assign es_rdata_capt_vld_d =
         !es_enable_fo[16] ? 1'b0 :
         es_rdata_capt_vld ? 1'b1 :
         es_rdata_capt_vld_q;

  // continuous compare of the entropy data
  assign es_bus_cmp_alert = es_rdata_capt_vld && es_rdata_capt_vld_q &&
         (es_rdata_capt_q == sfifo_esfinal_rdata[63:0]);


  //--------------------------------------------
  // software es read path
  //--------------------------------------------

  prim_packer_fifo #(
    .InW(SeedLen),
    .OutW(FullRegWidth),
    .ClearOnRead(1'b0)
  ) u_prim_packer_fifo_swread (
    .clk_i      (clk_i),
    .rst_ni     (rst_ni),
    .clr_i      (pfifo_swread_clr),
    .wvalid_i   (pfifo_swread_push),
    .wdata_i    (pfifo_swread_wdata),
    .wready_o   (pfifo_swread_not_full),
    .rvalid_o   (pfifo_swread_not_empty),
    .rdata_o    (pfifo_swread_rdata),
    .rready_i   (pfifo_swread_pop),
    .depth_o    ()
  );

  assign pfifo_swread_push = es_route_to_sw && pfifo_swread_not_full && sfifo_esfinal_not_empty;
  assign pfifo_swread_wdata = esfinal_data;

  assign pfifo_swread_clr = !(es_enable_fo[17] && es_data_reg_rd_en);
  assign pfifo_swread_pop =  es_enable_fo[18] && sw_es_rd_pulse;

  // set the es entropy to the read reg
  assign es_data_reg_rd_en = es_enable_fo[19] && efuse_es_sw_reg_en && entropy_data_reg_en_pfe;
  assign hw2reg.entropy_data.d = es_data_reg_rd_en ? pfifo_swread_rdata : '0;
  assign sw_es_rd_pulse = es_data_reg_rd_en && reg2hw.entropy_data.re;

  assign efuse_es_sw_reg_en = prim_mubi_pkg::mubi8_test_true_strict(en_entropy_src_fw_read);

  prim_mubi8_sync #(
    .NumCopies(1),
    .AsyncOn(1) // must be set to one, see note below
  ) u_prim_mubi8_sync_es_fw_read (
    .clk_i,
    .rst_ni,
    .mubi_i(otp_en_entropy_src_fw_read_i),
    .mubi_o({en_entropy_src_fw_read})
  );

  // note: the input to the above sync module is from the OTP block.
  //       It is assumed that the source is in a different time domain,
  //       and requires the AsyncOn parameter to be set.


  //--------------------------------------------
  // unused signals
  //--------------------------------------------

  assign unused_err_code_test_bit = (|{err_code_test_bit[27:25],err_code_test_bit[19:3]});
  assign unused_sha3_state = (|sha3_state[0][sha3_pkg::StateW-1:SeedLen]);
  assign unused_entropy_data = (|reg2hw.entropy_data.q);
  assign unused_fw_ov_rd_data = (|reg2hw.fw_ov_rd_data.q);

  //--------------------------------------------
  // Assertions
  //--------------------------------------------

`ifdef INC_ASSERT
  // entropy_src is known to activate Keccak without AES Halt handshakes with CSRNG (#17941).
  // This code ensures that this does not happen too often (i.e., at most `KAWAH_THRESHOLD` out of
  // `KAWAH_WINDOW_SIZE` consecutive clock cycles) outside *Firmware Override - Extract & Insert*
  // mode.  When firmware inserts entropy, it is essentially in control of the SHA3 core
  // and the current HW implementation cannot make guarantees around AES Halt and Keccak activity.
  //
  // When issue #17941 gets resolved and there are assertions (or equivalent checks) in place to
  // ensure that Keccak is not activated without AES Halt handshakes, this code should be removed.

  // Track activity of Keccak.
  logic keccak_active;
  assign keccak_active = u_sha3.u_keccak.keccak_st != sha3_pkg::KeccakStIdle;
  `ASSERT_KNOWN(KeccakActiveKnown_A, keccak_active)

  // Track state of AES Halt req/ack with CSRNG.
  logic cs_aes_halt_active;
  assign cs_aes_halt_active = cs_aes_halt_o.cs_aes_halt_req && cs_aes_halt_i.cs_aes_halt_ack;
  `ASSERT_KNOWN(CsAesHaltActiveKnown_A, cs_aes_halt_active)

  // Track when Keccak is active without AES Halt ('KAWAH') outside FW entropy insertion mode.
  localparam int unsigned KAWAH_WINDOW_SIZE = 512;
  logic [KAWAH_WINDOW_SIZE-1:0] kawah_window_d, kawah_window_q;
  assign kawah_window_d[0] = keccak_active & ~cs_aes_halt_active & ~fw_ov_mode_entropy_insert;
  assign kawah_window_d[KAWAH_WINDOW_SIZE-1:1] = kawah_window_q[KAWAH_WINDOW_SIZE-2:0];

  // Count how many cycles Keccak was active without AES Halt in the current window.
  localparam int unsigned KAWAH_COUNTER_SIZE = $clog2(KAWAH_WINDOW_SIZE);
  logic [KAWAH_COUNTER_SIZE-1:0] kawah_counter_d, kawah_counter_q;
  always_comb begin
    kawah_counter_d = kawah_counter_q;
    // Increment counter if Keccak is active without AES Halt in the current cycle.
    if (kawah_window_d[0]) kawah_counter_d += 1;
    // Decrement counter if Keccak was active without AES Halt in the cycle that falls out of the
    // sliding window in this cycle.
    if (kawah_window_q[KAWAH_WINDOW_SIZE-1]) begin
      // If the counter would underflow, a testbench error has happened (only relevant if reset is
      // deasserted).
      `ASSERT_I(KawahCounterNoUnderflow_A, rst_ni !== 1'b1 || kawah_counter_d > 0)
      kawah_counter_d -= 1;
    end
  end
  // Ensure counter does not overflow.
  `ASSERT(KawahCounterNoOverflow_A, kawah_counter_d < KAWAH_WINDOW_SIZE - 1)

  // Assert that in the last KAWAH_WINDOW_SIZE clock cycles, Keccak was active without AES Halt for
  // at most KAWAH_THRESHOLD clock cycles.
  localparam int unsigned KAWAH_THRESHOLD = 24;
  `ASSERT(KeccakNotTooActiveWithoutAesHalt_A, kawah_counter_q <= KAWAH_THRESHOLD)
  `ASSERT_INIT(KawahParametersLegal_A, KAWAH_THRESHOLD < KAWAH_WINDOW_SIZE)

  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      kawah_counter_q <= '0;
      kawah_window_q  <= '0;
    end else begin
      kawah_counter_q <= kawah_counter_d;
      kawah_window_q  <= kawah_window_d;
    end
  end
`endif

  //--------------------------------------------
  // Assertions
  //--------------------------------------------
`ifdef INC_ASSERT
`include "prim_macros.svh"

  // Count number of disables since last reset.
  logic [63:0] disable_cnt_d, disable_cnt_q;
  always_comb begin
    disable_cnt_d = disable_cnt_q;
    if (!mubi4_test_true_strict(mubi_mod_en_dly_d) &&
        mubi4_test_true_strict(mubi_mod_en_dly_q)) begin
      disable_cnt_d += 1;
    end
  end

  // Assert that no entropy gets dropped during FIPS-compliant operation mode.
  //
  // The following code, which includes counters, small FSMs, and assertions, tracks entropy bits
  // from the noise source input through Entropy Source to the hardware interface output and checks
  // that in FIPS-compliant mode entropy does not get dropped unless it should get dropped.  The
  // code is arranged in the same order as entropy flows through Entropy Source, so having Entropy
  // Source's block diagram ready when reading this code is highly recommended.

  // Delay `es_delayed_enable` by one clock cycle to track when Entropy Source actually accepts RNG
  // inputs.
  logic es_delayed_enable_d, es_delayed_enable_q;
  assign es_delayed_enable_d = es_delayed_enable;

  // Count number of valid bits from RNG input (RNG_BUS_WIDTH wide) while Entropy Source is enabled.
  logic [63:0] rng_valid_bit_cnt_d, rng_valid_bit_cnt_q;
  assign rng_valid_bit_cnt_d = entropy_src_rng_i.rng_valid && es_delayed_enable_q ?
                               rng_valid_bit_cnt_q + RNG_BUS_WIDTH :
                               rng_valid_bit_cnt_q;

  // Count number of bits pushed into esrng FIFO (RngBusWidth wide).
  logic [63:0] esrng_push_bit_cnt_d, esrng_push_bit_cnt_q;
  assign esrng_push_bit_cnt_d = sfifo_esrng_push & sfifo_esrng_not_full ?
                                esrng_push_bit_cnt_q + RngBusWidth :
                                esrng_push_bit_cnt_q;

  // Assert that as many bits got pushed into the esrng FIFO (destination) as there were valid RNG
  // input bits (source).  RngBusWidth bits may get lost after every re-enable; add a margin to
  // account for that.
  `ASSERT_AT_RESET_AND_FINAL(ValidRngBitsPushedIntoEsrngFifo_A,
                             `WITHIN_MARGIN(esrng_push_bit_cnt_q,        // actual
                                            rng_valid_bit_cnt_q,         // expected
                                            disable_cnt_q * RngBusWidth, // allowed less
                                            0))                          // allowed more

  // Count number of bits pushed into esbit FIFO (1 wide input, RngBusWidth wide output).
  logic [63:0] esbit_push_bit_cnt_d, esbit_push_bit_cnt_q;
  assign esbit_push_bit_cnt_d = pfifo_esbit_push & pfifo_esbit_not_full ?
                                esbit_push_bit_cnt_q + 1 :
                                esbit_push_bit_cnt_q;

  // Count number of bits pushed into postht FIFO (RngBusWidth wide input, PostHTWidth wide output).
  logic [63:0] postht_push_bit_cnt_d, postht_push_bit_cnt_q;
  assign postht_push_bit_cnt_d = pfifo_postht_push & pfifo_postht_not_full ?
                                 postht_push_bit_cnt_q + RngBusWidth :
                                 postht_push_bit_cnt_q;

  // Count number of bits pushed into postht FIFO from esrng FIFO.
  logic [63:0] postht_from_esrng_push_bit_cnt_d, postht_from_esrng_push_bit_cnt_q;
  assign postht_from_esrng_push_bit_cnt_d =
      pfifo_postht_push & pfifo_postht_not_full & ~rng_bit_en ?
      postht_from_esrng_push_bit_cnt_q + RngBusWidth :
      postht_from_esrng_push_bit_cnt_q;

  // Assert that as many bits got pushed into the esbit FIFO or the postht FIFO (destinations) as
  // into the esrng FIFO (source).  The number of bits pushed into the esbit FIFO has to be
  // multiplied by the output width of the esrng FIFO (RngBusWidth) because only 1 bit gets pushed
  // into the esbit FIFO for every pop from the esrng FIFO.  Add a margin (allowed less) because:
  // - RngBusWidth bits may get lost after every re-enable
  // - one entry may just have been pushed into esrng FIFO when the assertion gets evaluated.
  `ASSERT_AT_RESET_AND_FINAL(EsrngFifoPushedIntoEsbitOrPosthtFifos_A,
                             `WITHIN_MARGIN((esbit_push_bit_cnt_q * RngBusWidth +
                                             postht_from_esrng_push_bit_cnt_q), // actual
                                            esrng_push_bit_cnt_q,               // expected
                                            (disable_cnt_q + 1) * RngBusWidth,  // allowed less
                                            0))                                 // allowed more

  // Count number of bits pushed into postht FIFO from esbit FIFO.
  logic [63:0] postht_from_esbit_push_bit_cnt_d, postht_from_esbit_push_bit_cnt_q;
  assign postht_from_esbit_push_bit_cnt_d =
      pfifo_postht_push & pfifo_postht_not_full & rng_bit_en ?
      postht_from_esbit_push_bit_cnt_q + RngBusWidth :
      postht_from_esbit_push_bit_cnt_q;

  // Assert that as many bits got pushed into the postht FIFO (destination) as into the esbit FIFO
  // (source) when the latter was selected as source.  Add a margin (allowed less) because:
  // - RngBusWidth bits may get lost after every re-enable
  // - esbit FIFO may be partially full when the assertion gets evaluated.
  `ASSERT_AT_RESET_AND_FINAL(EsbitFifoPushedIntoPosthtFifo_A,
                             `WITHIN_MARGIN(postht_from_esbit_push_bit_cnt_q,      // actual
                                            esbit_push_bit_cnt_q,                  // expected
                                            (disable_cnt_q + 1) * RngBusWidth - 1, // allowed less
                                            0))                                    // allowed more

  // Assert that as many bits got pushed into the postht FIFO as got counted from the esrng FIFO or
  // the esbit FIFO.  This assertion checks more the completeness of the other assertions than the
  // design itself.
  `ASSERT_AT_RESET_AND_FINAL(PosthtFifoPushedFromEsbitOrEsrngFifos_A,
                             postht_push_bit_cnt_q == (postht_from_esrng_push_bit_cnt_q +
                                                       postht_from_esbit_push_bit_cnt_q))

  // Count number of bits popped from postht FIFO (PostHTWidth wide output) when bypass mode was
  // disabled.
  logic [63:0] postht_non_bypass_pop_bit_cnt_d, postht_non_bypass_pop_bit_cnt_q;
  assign postht_non_bypass_pop_bit_cnt_d =
      pfifo_postht_pop & pfifo_postht_not_empty & ~es_bypass_mode ?
      postht_non_bypass_pop_bit_cnt_q + PostHTWidth :
      postht_non_bypass_pop_bit_cnt_q;

  // Count number of bits pushed into precon FIFO (ObserveFifoWidth wide input, PreCondWidth wide
  // output).
  logic [63:0] precon_push_bit_cnt_d, precon_push_bit_cnt_q;
  assign precon_push_bit_cnt_d = pfifo_precon_push & pfifo_precon_not_full ?
                                 precon_push_bit_cnt_q + ObserveFifoWidth :
                                 precon_push_bit_cnt_q;

  // Assert that as many bits got pushed into the precon FIFO (destination) as got popped from the
  // postht FIFO when bypass mode was disabled (source).
  `ASSERT_AT_RESET_AND_FINAL(PosthtFifoPushedIntoPreconFifo_A,
                             precon_push_bit_cnt_q == postht_non_bypass_pop_bit_cnt_q)

  // Track when boot and startup checks are completing.
  logic boot_startup_checks_completing;
  assign boot_startup_checks_completing =
      (u_entropy_src_main_sm.state_q == entropy_src_main_sm_pkg::StartupPass1 &
       u_entropy_src_main_sm.ht_done_pulse_i &
       ~u_entropy_src_main_sm.ht_fail_pulse_i);

  // Track state of boot and startup checks.
  typedef enum logic [1:0] {
    BscStIncomplete,  // checks incomplete
    BscStPassed,      // checks passed
    BscStPushed       // entropy from passed checks pushed
  } bsc_state_e;
  bsc_state_e bsc_state_d, bsc_state_q;
  always_comb begin
    bsc_state_d = bsc_state_q;
    unique case (bsc_state_q)
      BscStIncomplete: begin
        if (boot_startup_checks_completing) begin
          // Checks have just completed.
          bsc_state_d = BscStPassed;
        end
      end
      BscStPassed: begin
        if (main_stage_push) begin
          // Entropy from passed checks is being pushed.
          bsc_state_d = BscStPushed;
        end
      end
      BscStPushed: begin
        // Boot and startup checks remained passed and their entropy pushed until Entropy Source
        // gets disabled again (which is handled below).
        bsc_state_d = bsc_state_q;
      end
      default: bsc_state_d = BscStIncomplete;
    endcase
    // If not enabled, always clear to incomplete.
    if (!mubi4_test_true_strict(mubi_es_enable)) begin
      bsc_state_d = BscStIncomplete;
    end
  end

  // Count number of bits pushed into precon FIFO (ObserveFifoWidth wide input, PreCondWidth wide
  // output) after boot and startup checks.
  logic [63:0] precon_post_startup_push_bit_cnt_d, precon_post_startup_push_bit_cnt_q;
  assign precon_post_startup_push_bit_cnt_d =
      pfifo_precon_push & pfifo_precon_not_full & (bsc_state_q != BscStIncomplete) ?
      precon_post_startup_push_bit_cnt_q + ObserveFifoWidth :
      precon_post_startup_push_bit_cnt_q;

  // Track when esfinal FIFO gets pushed while bypass mode is disabled.
  logic esfinal_non_bypass_push;
  assign esfinal_non_bypass_push = sfifo_esfinal_push & sfifo_esfinal_not_full & ~es_bypass_mode;

  // Count number of bits pushed into esfinal FIFO (SeedLen bits per push) while bypass mode was
  // disabled.
  logic [63:0] esfinal_non_bypass_push_cnt_d, esfinal_non_bypass_push_cnt_q;
  assign esfinal_non_bypass_push_cnt_d = esfinal_non_bypass_push ?
                                         esfinal_non_bypass_push_cnt_q + SeedLen :
                                         esfinal_non_bypass_push_cnt_q;

  // Count number of bits pushed into esfinal FIFO (SeedLen bits per push) after startup checks have
  // passed and while bypass mode was disabled.
  logic [63:0] esfinal_post_startup_push_bit_cnt_d, esfinal_post_startup_push_bit_cnt_q;
  assign esfinal_post_startup_push_bit_cnt_d =
      esfinal_non_bypass_push & (bsc_state_q != BscStIncomplete) ?
      esfinal_post_startup_push_bit_cnt_q + SeedLen :
      esfinal_post_startup_push_bit_cnt_q;

  // Assert that all bits pushed into the esfinal FIFO came from or after passed startup checks.
  `ASSERT_AT_RESET_AND_FINAL(EsfinalFifoPushed_A,
                             esfinal_non_bypass_push_cnt_q == esfinal_post_startup_push_bit_cnt_q)

  // Track result of health tests after boot and startup tests.
  typedef enum logic [1:0] {
    HtStNoResult, // no health test result is currently available
    HtStPassed,   // last health test has passed and entropy has not propagated from conditioner yet
    HtStFailed    // last health test has failed
  } ht_state_e;
  ht_state_e ht_state_d, ht_state_q;
  always_comb begin
    ht_state_d = ht_state_q;
    if (bsc_state_q == BscStPushed) begin
      if (ht_state_q inside {HtStNoResult, HtStFailed}) begin
        if (health_test_done_pulse) begin
          if (!any_fail_pulse && !alert_threshold_fail) begin
            ht_state_d = HtStPassed;
          end else begin
            ht_state_d = HtStFailed;
          end
        end
      end else if (ht_state_q == HtStPassed) begin
        if (main_stage_push_raw) begin
          ht_state_d = HtStNoResult;
        end
      end else begin
        ht_state_d = HtStNoResult;
      end
      if (ht_state_q == HtStFailed) begin
        `ASSERT_I(NoPushAfterFailedHealthTest_A, rst_ni !== 1'b1 || !main_stage_push_raw)
      end
    end
    // If not enabled, always clear to no result.
    if (!mubi4_test_true_strict(mubi_es_enable)) begin
      ht_state_d = HtStNoResult;
    end
  end

  // Track when entropy is expected to get dropped instead of pushed into the esfinal FIFO: when the
  // esfinal FIFO is full and either routing to SW and the SW read FIFO is full or not routing to SW
  // and no request on the hardware interface.
  logic esfinal_exp_drop;
  assign esfinal_exp_drop = sfifo_esfinal_full & (es_route_to_sw ?
                                                  ~pfifo_swread_not_full :      // SW read FIFO full
                                                  ~entropy_src_hw_if_i.es_req); // no HW request

  // Count number of bits that are expected to have gotten pushed into precon FIFO and into esfinal
  // FIFO after boot and startup checks and while bypass mode was disabled.
  logic [63:0] precon_post_startup_exp_push_bit_cnt_d, precon_post_startup_exp_push_bit_cnt_q;
  logic [63:0] esfinal_post_startup_exp_push_bit_cnt_d, esfinal_post_startup_exp_push_bit_cnt_q;
  always_comb begin
    esfinal_post_startup_exp_push_bit_cnt_d = esfinal_post_startup_exp_push_bit_cnt_q;
    precon_post_startup_exp_push_bit_cnt_d = precon_post_startup_exp_push_bit_cnt_q;
    if (bsc_state_q == BscStPassed && bsc_state_d == BscStPushed) begin
      // On the completion of boot and startup checks, SeedLen bits are expected to be pushed into
      // the esfinal FIFO.
      esfinal_post_startup_exp_push_bit_cnt_d += SeedLen;
    end
    if (bsc_state_q != BscStIncomplete && health_test_done_pulse) begin
      // Once boot and startup checks have completed, (4 * health_test_window) bits are expected to
      // have gotten pushed into the precon FIFO.
      precon_post_startup_exp_push_bit_cnt_d += 4 * health_test_window;
    end
    if (ht_state_q == HtStPassed && main_stage_push_raw && !esfinal_exp_drop) begin
      // If none of the health tests failed and the alert threshold has not been exceeded, SeedLen
      // bits are expected to be pushed into the esfinal FIFO -- unless we expect them to get
      // dropped (see above).
      esfinal_post_startup_exp_push_bit_cnt_d += SeedLen;
    end
    // When Entropy Source gets disabled after boot and startup checks have been completed, add the
    // number of bits that have been pushed into precon FIFO since the last conditioner output to
    // the expected number of bits.
    if ((bsc_state_q != BscStIncomplete) && (bsc_state_d == BscStIncomplete)) begin
      logic [63:0] diff_;
      diff_ = precon_post_startup_push_bit_cnt_q - precon_post_startup_exp_push_bit_cnt_q;
      // Assert that the difference is not negative.
      `ASSERT_I(PreconPostStartupDiffNonNegative_A,
                rst_ni !== 1'b1 || (precon_post_startup_push_bit_cnt_q >=
                                    precon_post_startup_exp_push_bit_cnt_q))
      // Assert that the difference is smaller than the number of bits that would have sufficed to
      // get pushed into the conditioner.
      `ASSERT_I(PreconPostStartupDiffSmall_A, rst_ni !== 1'b1 || diff_ < (4 * health_test_window))
      precon_post_startup_exp_push_bit_cnt_d += diff_;
    end
  end
  // This code assumes that `health_test_window` does not change dynamically; capture that in an
  // assertion ensuring it only changes when entropy_src is not enabled.
  `ASSERT(HealthTestWindowStableWhenEnabled_A,
          mubi4_test_true_strict(mubi_es_enable) |-> $stable(health_test_window))

  // Assert that all bits pushed into the esfinal FIFO after startup checks were expected.
  `ASSERT_AT_RESET_AND_FINAL(EsfinalFifoPushedPostStartup_A,
                             esfinal_post_startup_push_bit_cnt_q ==
                             esfinal_post_startup_exp_push_bit_cnt_q)

  // Assert that the expected number of bits pushed into the precon FIFO based on the number of
  // outputs of the conditioner matches the actual number of bits pushed into the precon FIFO after
  // startup checks.  Add a margin (allowed more) as the simulation may end when bits in the precon
  // FIFO have not resulted in conditioner output and Entropy Source has not been disabled.
  logic [63:0] ppspb_allowed_more;
  assign ppspb_allowed_more = bsc_state_q != BscStIncomplete ? 4 * health_test_window : '0;
  `ASSERT_AT_RESET_AND_FINAL(PreconFifoPushedPostStartup_A,
                             `WITHIN_MARGIN(precon_post_startup_push_bit_cnt_q,     // actual
                                            precon_post_startup_exp_push_bit_cnt_q, // expected
                                            0,                                      // allowed less
                                            ppspb_allowed_more))                    // allowed more

  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      esbit_push_bit_cnt_q                <= '0;
      esfinal_non_bypass_push_cnt_q       <= '0;
      esfinal_post_startup_push_bit_cnt_q <= '0;
      esrng_push_bit_cnt_q                <= '0;
      postht_from_esbit_push_bit_cnt_q    <= '0;
      postht_from_esrng_push_bit_cnt_q    <= '0;
      postht_non_bypass_pop_bit_cnt_q     <= '0;
      postht_push_bit_cnt_q               <= '0;
      precon_post_startup_push_bit_cnt_q  <= '0;
      precon_push_bit_cnt_q               <= '0;
      rng_valid_bit_cnt_q                 <= '0;
    end else if (mubi4_test_true_strict(mubi_es_enable) & !fw_ov_mode_entropy_insert) begin
      // All these counters get updated if and only if entropy_src is enabled and the firmware
      // override entropy insertion mode is disabled.  Otherwise, there are no guarantees on how
      // much entropy from the noise source gets dropped due to backpressure.
      esbit_push_bit_cnt_q                <= esbit_push_bit_cnt_d;
      esfinal_non_bypass_push_cnt_q       <= esfinal_non_bypass_push_cnt_d;
      esfinal_post_startup_push_bit_cnt_q <= esfinal_post_startup_push_bit_cnt_d;
      esrng_push_bit_cnt_q                <= esrng_push_bit_cnt_d;
      postht_from_esbit_push_bit_cnt_q    <= postht_from_esbit_push_bit_cnt_d;
      postht_from_esrng_push_bit_cnt_q    <= postht_from_esrng_push_bit_cnt_d;
      postht_non_bypass_pop_bit_cnt_q     <= postht_non_bypass_pop_bit_cnt_d;
      postht_push_bit_cnt_q               <= postht_push_bit_cnt_d;
      precon_post_startup_push_bit_cnt_q  <= precon_post_startup_push_bit_cnt_d;
      precon_push_bit_cnt_q               <= precon_push_bit_cnt_d;
      rng_valid_bit_cnt_q                 <= rng_valid_bit_cnt_d;
    end
  end

  always_ff @(posedge clk_i, negedge rst_ni) begin
    if (!rst_ni) begin
      bsc_state_q                             <= BscStIncomplete;
      disable_cnt_q                           <= '0;
      es_delayed_enable_q                     <= '0;
      esfinal_post_startup_exp_push_bit_cnt_q <= '0;
      ht_state_q                              <= HtStNoResult;
      precon_post_startup_exp_push_bit_cnt_q  <= '0;
    end else begin
      bsc_state_q                             <= bsc_state_d;
      disable_cnt_q                           <= disable_cnt_d;
      es_delayed_enable_q                     <= es_delayed_enable_d;
      esfinal_post_startup_exp_push_bit_cnt_q <= esfinal_post_startup_exp_push_bit_cnt_d;
      ht_state_q                              <= ht_state_d;
      precon_post_startup_exp_push_bit_cnt_q  <= precon_post_startup_exp_push_bit_cnt_d;
    end
  end
`endif

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description: entropy_src top level wrapper file

`include "prim_assert.sv"


module entropy_src
  import entropy_src_pkg::*;
  import entropy_src_reg_pkg::*;
  import prim_mubi_pkg::mubi8_t;
#(
  parameter bit Stub = 1'b0,
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},
  parameter int EsFifoDepth = 4
) (
  input logic clk_i,
  input logic rst_ni,

  // Bus Interface
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // OTP Interface
  // SEC_CM: INTERSIG.MUBI
  input  mubi8_t otp_en_entropy_src_fw_read_i,
  // SEC_CM: INTERSIG.MUBI
  input  mubi8_t otp_en_entropy_src_fw_over_i,

  // RNG Interface
  output logic rng_fips_o,

  // Entropy Interface
  input  entropy_src_hw_if_req_t entropy_src_hw_if_i,
  output entropy_src_hw_if_rsp_t entropy_src_hw_if_o,

  // RNG Interface
  output entropy_src_rng_req_t entropy_src_rng_o,
  input  entropy_src_rng_rsp_t entropy_src_rng_i,

  // CSRNG Interface
  output cs_aes_halt_req_t cs_aes_halt_o,
  input  cs_aes_halt_rsp_t cs_aes_halt_i,

  // External Health Test Interface
  output entropy_src_xht_req_t entropy_src_xht_o,
  input  entropy_src_xht_rsp_t entropy_src_xht_i,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // Interrupts
  output logic    intr_es_entropy_valid_o,
  output logic    intr_es_health_test_failed_o,
  output logic    intr_es_observe_fifo_ready_o,
  output logic    intr_es_fatal_err_o
);

  localparam int RngBusWidth = 4; // AST RNG bus width
  localparam int NumBins = 2**RngBusWidth; // bucket health test bin count

  // common signals
  entropy_src_hw2reg_t hw2reg;
  entropy_src_reg2hw_t reg2hw;
  logic [NumAlerts-1:0] alert_test;
  logic [NumAlerts-1:0] alert;

  // core signals
  logic core_rst_n;
  entropy_src_hw2reg_t core_hw2reg;
  entropy_src_hw_if_rsp_t core_entropy_hw_if;
  entropy_src_rng_req_t core_rng;
  cs_aes_halt_req_t core_aes_halt;
  entropy_src_xht_req_t core_xht;
  logic core_intr_es_entropy_valid;
  logic core_intr_es_health_test_failed;
  logic core_intr_es_observe_fifo_ready;
  logic core_intr_es_fatal_err;
  logic [NumAlerts-1:0] core_alert_test;
  logic [NumAlerts-1:0] core_alert;

  //stub signals
  localparam int StubLfsrWidth = 64;
  localparam int Copies = CSRNG_BUS_WIDTH / StubLfsrWidth;
  entropy_src_hw2reg_t stub_hw2reg;
  entropy_src_hw_if_rsp_t stub_entropy_hw_if;
  logic stub_es_valid;
  logic [NumAlerts-1:0] stub_alert_test;
  logic [NumAlerts-1:0] stub_alert;
  logic [StubLfsrWidth-1:0] stub_lfsr_value;

  ///////////////////////////
  // Selecting between core and stub
  ///////////////////////////

  assign hw2reg                       = Stub ? stub_hw2reg        : core_hw2reg;
  assign core_rst_n                   = Stub ? '0                 : rst_ni;
  assign entropy_src_hw_if_o          = Stub ? stub_entropy_hw_if : core_entropy_hw_if;
  assign entropy_src_rng_o            = Stub ? '1                 : core_rng;
  assign cs_aes_halt_o                = Stub ? '0                 : core_aes_halt;
  assign entropy_src_xht_o            = Stub ? '0                 : core_xht;
  assign intr_es_entropy_valid_o      = Stub ? stub_es_valid      : core_intr_es_entropy_valid;
  assign intr_es_health_test_failed_o = Stub ? '0                 : core_intr_es_health_test_failed;
  assign intr_es_observe_fifo_ready_o = Stub ? '0                 : core_intr_es_observe_fifo_ready;
  assign intr_es_fatal_err_o          = Stub ? '0                 : core_intr_es_fatal_err;
  assign alert_test                   = Stub ? stub_alert_test    : core_alert_test;
  assign alert                        = Stub ? stub_alert         : core_alert;

  ///////////////////////////
  // core entropy operation
  ///////////////////////////

  logic [NumAlerts-1:0] intg_err_alert;
  assign intg_err_alert[0] = 1'b0;

  // SEC_CM: CONFIG.REGWEN
  // SEC_CM: TILE_LINK.BUS.INTEGRITY

  entropy_src_reg_top u_reg (
    .clk_i,
    .rst_ni,
    .tl_i,
    .tl_o,
    .reg2hw,
    .hw2reg(hw2reg),
    .intg_err_o(intg_err_alert[1]), // Assign this alert to the fatal alert index.
    .devmode_i(1'b1)
  );

  entropy_src_core #(
    .EsFifoDepth(EsFifoDepth)
  ) u_entropy_src_core (
    .clk_i,
    .rst_ni(core_rst_n),
    .reg2hw,
    .hw2reg(core_hw2reg),

    .otp_en_entropy_src_fw_read_i(otp_en_entropy_src_fw_read_i),
    .otp_en_entropy_src_fw_over_i(otp_en_entropy_src_fw_over_i),
    .rng_fips_o,

    .entropy_src_hw_if_o(core_entropy_hw_if),
    .entropy_src_hw_if_i,

    .entropy_src_xht_o(core_xht),
    .entropy_src_xht_i,

    .entropy_src_rng_o(core_rng),
    .entropy_src_rng_i,

    .cs_aes_halt_o(core_aes_halt),
    .cs_aes_halt_i,

    .recov_alert_o(core_alert[0]),
    .fatal_alert_o(core_alert[1]),

    .recov_alert_test_o(core_alert_test[0]),
    .fatal_alert_test_o(core_alert_test[1]),

    .intr_es_entropy_valid_o(core_intr_es_entropy_valid),
    .intr_es_health_test_failed_o(core_intr_es_health_test_failed),
    .intr_es_observe_fifo_ready_o(core_intr_es_observe_fifo_ready),
    .intr_es_fatal_err_o(core_intr_es_fatal_err)
  );

  ///////////////////////////
  // stub entropy operation
  ///////////////////////////

  assign stub_alert = '0;
  assign stub_alert_test = '0;
  assign stub_entropy_hw_if = '{
    es_ack:  '1,
    es_bits:  {Copies{stub_lfsr_value}},
    es_fips: '1
  };
  // once enabled, stub entropy is always available

  import prim_mubi_pkg::mubi4_t;
  import prim_mubi_pkg::mubi4_test_true_strict;

  mubi4_t mubi_module_en;
  assign mubi_module_en  = mubi4_t'(reg2hw.module_enable.q);
  assign stub_es_valid = mubi4_test_true_strict(mubi_module_en);

  if (Stub) begin : gen_stub_entropy_src
    prim_lfsr #(
      .LfsrDw(StubLfsrWidth),
      .StateOutDw(StubLfsrWidth)
    ) u_prim_lfsr (
      .clk_i          (clk_i),
      .rst_ni         (rst_ni),
      .seed_en_i      ('0),
      .seed_i         ('0),
      .lfsr_en_i      (stub_es_valid),
      .entropy_i      ('0),
      .state_o        (stub_lfsr_value)
    );

    // hardwire hw2reg inputs
    always_comb begin
      stub_hw2reg = '0;

      // as long as enable is 1, do not allow registers to be written
      stub_hw2reg.fw_ov_rd_data.d = stub_lfsr_value[31:0];
      stub_hw2reg.entropy_data.d = stub_lfsr_value[31:0];
      stub_hw2reg.debug_status.main_sm_idle.d = 1'b1;
      // need to move this to package so that it can be referenced
      stub_hw2reg.debug_status.main_sm_state.d = 8'b01110110;

      stub_hw2reg.intr_state.es_entropy_valid.de = stub_es_valid;
      stub_hw2reg.intr_state.es_entropy_valid.d = 1'b1;

    end
  end else begin : gen_stub_tieoff
    assign stub_hw2reg = '0;
    assign stub_lfsr_value = '0;
  end

  ///////////////////////////
  // Alert generation
  ///////////////////////////
  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i)
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i]                 ),
      .alert_req_i   ( alert[i] || intg_err_alert[i] ),
      .alert_ack_o   (                               ),
      .alert_state_o (                               ),
      .alert_rx_i    ( alert_rx_i[i]                 ),
      .alert_tx_o    ( alert_tx_o[i]                 )
    );
  end

  // Outputs should have a known value after reset
  `ASSERT_KNOWN(TlDValidKnownO_A, tl_o.d_valid)
  `ASSERT_KNOWN(TlAReadyKnownO_A, tl_o.a_ready)

  // Entropy Interface
  `ASSERT_KNOWN(EsHwIfEsAckKnownO_A, entropy_src_hw_if_o.es_ack)
  `ASSERT_KNOWN_IF(EsHwIfEsBitsKnownO_A, entropy_src_hw_if_o.es_bits,
      entropy_src_hw_if_o.es_ack)
  `ASSERT_KNOWN_IF(EsHwIfEsFipsKnownO_A, entropy_src_hw_if_o.es_fips,
      entropy_src_hw_if_o.es_ack)

  // RNG Interface
  `ASSERT_KNOWN(EsRngEnableKnownO_A, entropy_src_rng_o.rng_enable)

  // External Health Test Interface
  `ASSERT_KNOWN_IF(EsXhtEntropyBitKnownO_A, entropy_src_xht_o.entropy_bit,
      entropy_src_xht_o.entropy_bit_valid)
  `ASSERT_KNOWN(EsXhtEntropyBitValidKnownO_A, entropy_src_xht_o.entropy_bit_valid)
  `ASSERT_KNOWN(EsXhtClearKnownO_A, entropy_src_xht_o.clear)
  `ASSERT_KNOWN(EsXhtActiveKnownO_A, entropy_src_xht_o.active)
  `ASSERT_KNOWN(EsXhtThreshHiKnownO_A, entropy_src_xht_o.thresh_hi)
  `ASSERT_KNOWN(EsXhtThreshLoKnownO_A, entropy_src_xht_o.thresh_lo)
  `ASSERT_KNOWN(EsXhtWindowKnownO_A, entropy_src_xht_o.window_wrap_pulse)

  // Alerts
  `ASSERT_KNOWN(AlertTxKnownO_A, alert_tx_o)

  // Interrupts
  `ASSERT_KNOWN(IntrEsEntropyValidKnownO_A, intr_es_entropy_valid_o)
  `ASSERT_KNOWN(IntrEsHealthTestFailedKnownO_A, intr_es_health_test_failed_o)
  `ASSERT_KNOWN(IntrEsFifoErrKnownO_A, intr_es_fatal_err_o)

  // prim_count alerts
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck0_A,
    u_entropy_src_core.u_prim_count_window_cntr,
    alert_tx_o[1])

  for (genvar sh = 0; sh < RngBusWidth; sh = sh+1) begin : gen_bit_cntrs
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck1_A,
      u_entropy_src_core.u_entropy_src_adaptp_ht.gen_cntrs[sh].u_prim_count_test_cnt,
      alert_tx_o[1])
  end : gen_bit_cntrs

  for (genvar i = 0; i < NumBins; i = i + 1) begin : gen_symbol_match
   `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck_A,
     u_entropy_src_core.u_entropy_src_bucket_ht.gen_symbol_match[i].u_prim_count_bin_cntr,
     alert_tx_o[1])
  end : gen_symbol_match

  for (genvar sh = 0; sh < RngBusWidth; sh = sh+1) begin : gen_pair_cntrs
   `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck_A,
     u_entropy_src_core.u_entropy_src_markov_ht.gen_cntrs[sh].u_prim_count_pair_cntr,
     alert_tx_o[1])
  end : gen_pair_cntrs

  for (genvar sh = 0; sh < RngBusWidth; sh = sh+1) begin : gen_rep_cntrs
   `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck_A,
     u_entropy_src_core.u_entropy_src_repcnt_ht.gen_cntrs[sh].u_prim_count_rep_cntr,
     alert_tx_o[1])
  end : gen_rep_cntrs

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck7_A,
    u_entropy_src_core.u_entropy_src_repcnts_ht.u_prim_count_rep_cntr,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlMainFsmCheck_A,
    u_entropy_src_core.u_entropy_src_main_sm.u_state_regs,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlAckFsmCheck_A,
    u_entropy_src_core.u_entropy_src_ack_sm.u_state_regs,
    alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(SHA3FsmCheck_A,
    u_entropy_src_core.u_sha3.u_state_regs, alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(KeccakRoundFsmCheck_A,
    u_entropy_src_core.u_sha3.u_keccak.u_state_regs, alert_tx_o[1])

  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(SHA3padFsmCheck_A,
    u_entropy_src_core.u_sha3.u_pad.u_state_regs, alert_tx_o[1])


  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(SentMsgCountCheck_A,
    u_entropy_src_core.u_sha3.u_pad.u_sentmsg_count, alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(RoundCountCheck_A,
    u_entropy_src_core.u_sha3.u_keccak.u_round_count, alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck8_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_repcnt.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck9_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_repcnts.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck10_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_adaptp_hi.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck11_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_adaptp_lo.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck12_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_bucket.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck13_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_markov_hi.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck14_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_markov_lo.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck15_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_extht_hi.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck16_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_extht_lo.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck17_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_any_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck18_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_repcnt_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck19_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_repcnts_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck20_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_adaptp_hi_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck21_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_adaptp_lo_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck22_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_bucket_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck23_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_markov_hi_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck24_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_markov_lo_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck25_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_extht_hi_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CntAlertCheck26_A,
    u_entropy_src_core.u_entropy_src_cntr_reg_extht_lo_alert_fails.u_prim_count_cntr_reg,
    alert_tx_o[1])

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// kmac_pkg

package kmac_pkg;
  parameter int MsgWidth = sha3_pkg::MsgWidth;
  parameter int MsgStrbW = sha3_pkg::MsgStrbW;

  // Message FIFO depth
  //
  // Assume entropy is ready always (if Share is reused as an entropy in Chi)
  // Then it takes 72 cycles to complete the Keccak round. While Keccak is in
  // operation, the module need to store the incoming messages to not degrade
  // the throughput.
  //
  // Based on the observation from HMAC case, the core usually takes 5 clocks
  // to fetch data and store into KMAC. So the core can push at most 14.5 X 4B
  // which is 58B. After that, Keccak can fetch the data from MSG_FIFO faster
  // rate than the core can push. To fetch 58B, it takes around 7~8 cycles.
  // For that time, the core only can push at most 2 DW. After that Keccak
  // waits the incoming message.
  //
  // So Message FIFO doesn't need full block size except the KMAC case, which
  // is delayed the operation by processing Function Name N, customization S,
  // and secret keys. But KMAC doesn't need high throughput anyway (72Mb/s).
  parameter int RegIntfWidth = 32; // 32bit interface
  parameter int RegLatency   = 5;  // 5 cycle to write one Word
  parameter int Sha3Latency  = 72; // Expected masked sha3 processing time 24x3

  // Total required buffer size while SHA3 is in processing
  parameter int BufferCycles   = (Sha3Latency + RegLatency - 1)/RegLatency;
  parameter int BufferSizeBits = RegIntfWidth * BufferCycles;

  // Required MsgFifoDepth. Adding slightly more buffer for margin
  parameter int MsgFifoDepth   = 2 + ((BufferSizeBits + MsgWidth - 1)/MsgWidth);
  parameter int MsgFifoDepthW  = $clog2(MsgFifoDepth+1);

  parameter int MsgWindowWidth = 32; // Register width
  parameter int MsgWindowDepth = 512; // 2kB space

  // Key related definitions
  // If this value is changed, please modify the logic inside kmac_core
  // that assigns the value into `encoded_key`
  parameter int MaxKeyLen = 512;

  // size of encode_string(Key)
  // $ceil($clog2(MaxKeyLen+1)/8)
  parameter int MaxEncodedKeyLenW = $clog2(MaxKeyLen+1);
  parameter int MaxEncodedKeyLenByte = (MaxEncodedKeyLenW + 8 - 1) / 8;
  parameter int MaxEncodedKeyLenSize = MaxEncodedKeyLenByte * 8;

  //                             Secret Key  left_encode(len(Key))
  //                             ----------  ------------------------
  parameter int MaxEncodedKeyW = MaxKeyLen + MaxEncodedKeyLenSize + 8;

  // key_len is SW configurable CSR.
  // Current KMAC allows 5 key length options.
  // This value determines the KMAC core how to map the value
  // from Secret Key register to key size block
  typedef enum logic [2:0] {
    Key128 = 3'b 000, // 128 bit secret key
    Key192 = 3'b 001, // 192 bit secret key
    Key256 = 3'b 010, // 256 bit secret key
    Key384 = 3'b 011, // 384 bit secret key
    Key512 = 3'b 100  // 512 bit secret key
  } key_len_e;


  // kmac_cmd_e defines the possible command sets that software issues via
  // !!CMD register. This is mainly to limit the error scenario that SW writes
  // multiple commands at once. Additionally they are sparse encoded to harden
  // against FI attacks
  //
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 5 -n 6 \
  //      -s 1891656028 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (50.00%)
  //  4: |||||||||||||||| (40.00%)
  //  5: |||| (10.00%)
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 5
  // Minimum Hamming weight: 3
  // Maximum Hamming weight: 4
  //
  typedef enum logic [5:0] {
    //CmdNone      = 6'b001011, // dec 10
    // CmdNone is manually set to all zero by design!
    // The minimum Hamming distance is still 3
    CmdNone      = 6'b000000, // dec  0
    CmdStart     = 6'b011101, // dec 29
    CmdProcess   = 6'b101110, // dec 46
    CmdManualRun = 6'b110001, // dec 49
    CmdDone      = 6'b010110  // dec 22
  } kmac_cmd_e;

  // Timer
  parameter int unsigned TimerPrescalerW = 10;
  parameter int unsigned EdnWaitTimerW   = 16;

  // Entropy Mode Selection : Should be matched to register package Enum value
  typedef enum logic [1:0] {
    EntropyModeNone = 2'h 0,
    EntropyModeEdn  = 2'h 1,
    EntropyModeSw   = 2'h 2
  } entropy_mode_e;

  // PRNG (kmac_entropy)
  parameter int unsigned EntropyLfsrW = 800;
  parameter int unsigned ChunkSizeEntropyLfsr = 32;
  parameter int unsigned NumChunksEntropyLfsr = EntropyLfsrW / ChunkSizeEntropyLfsr;

  // We use a single seed that is split down into chunks internally.
  // These LFSR parameters have been generated with
  // $ ./util/design/gen-lfsr-seed.py --width 800 --seed 3369807298 --prefix ""
  typedef logic [EntropyLfsrW-1:0] lfsr_seed_t;
  typedef logic [EntropyLfsrW-1:0][$clog2(EntropyLfsrW)-1:0] lfsr_perm_t;
  parameter lfsr_seed_t RndCnstLfsrSeedDefault = {
    32'h34a19ca3,
    256'he514d8e17a5630c287247dff3d354c022f581ace4b6c5736b5efa4160261ab0f,
    256'h6cb2915197ab3588982bcffc9cf3b46a250cebf728c0e76f0e680420d7f428f2,
    256'h092c1e308f7c8f9d8bacc20cd18fd586d58879654aa4851de224033bfdcbc578
  };
  parameter lfsr_perm_t RndCnstLfsrPermDefault = {
    64'hb1a3e87aeb4e69f0,
    256'h2d8a6ee2c9ac567b2aa401a639a2a8ea2553614c0a8daf672c06546fc0d35267,
    256'hc4572024bc116458dd0f1c10a8aef5c4ad9a788968d0d7ca7345c6b8f277a5d3,
    256'hec5da20f261826ed3c8992724e70db897060be51b07a96902e14a42d12d320f8,
    256'h187049b6c25f35d0e485cc4b9ef01dad2865b5e558926f380718b74394fe0f82,
    256'hd5395a7d0aa4845af814e8681107a4c793758572c9467493bf1248a48f1b40c2,
    256'h09319b55111d0401819685a43a06f0da441021a8c220b14f01d44e49c1683a82,
    256'hafeb980964aa050641f4205131d9d4741eb5dd658e603b8ed438cb1096628d42,
    256'h62c9d75ced78ed09a3ddbb60f533eef10aa5a54b478d61a06a4b326eb3402105,
    256'hc27d562c6d91b48440d6d06e543be9871628a4aa9b3d2e51fa0ac2eb89a17f6d,
    256'h207ad96caf25d1fcffab210c1aff12252346fe4d56a7cd9b8605c7fa638895a9,
    256'h60158cd3a1ce4f2f6cf5d48579ac14b1e5219ca8914e0507b635dc712554f6bb,
    256'h0ae412943a7596f4644a0c13646adc91d02c406a10d232791d3de9919eec5424,
    256'haa2cac5f556c15c647eb29365062daf6aa848e10b3f665abccca713036d9f1cb,
    256'h1c9bd4aaeb19c5ac01b1805e0d5479860870da49a55e8f386ca8232c728e2f61,
    256'h3007aa420758818e5312401372eaa00d21c70c7e1158d2e08a1b6ac0b820cb67,
    256'hf0ba4b5c0865ff04f0f9d0175817c65d81918e43e14b2f83d574bfa9c6e6deae,
    256'h64c22c2974a1d5c55e2367004b249d5a02fc566685ea33b6f73aaa0244b34412,
    256'hb1a12230adb1748dc1d956f9f10c8e1aa52f4702e06a16680d92226c830ec4ce,
    256'h4c2eead21f08c387c3f1de89eb33b983c748e848f68b54f256715221177c5a4a,
    256'h0a47d82741955626755ba1cc24e2ba40504111b9e26136be714c5bc0d330c3f7,
    256'h75e863de763270a993890d633c6897218e151943edd8b79ae145cf564b774613,
    256'h0b0a76c40e7e84c876640dc78260c09a85e92e5ab56c22c0e72a8669fe88ba10,
    256'h8b99e437c776f0cea0d144f285b6ab7259e12284f380ae3410171cd6a8b04415,
    256'he95081c8c57e3e526ad5b38019a5c1b5505540462157e7c7e68e6a6a16ac460a,
    256'h5d5578da28092c7cc927cb9c0ed614a79b0e32b4c5b6a269a40743bef42b5e29,
    256'hd9a75ecb5548a29e9d34ddda07c8404aabbf5479456731ece3785f6090c3f862,
    256'h6eb1a5119e8b8e56b1455d820b46e20e15bb7d185a636b10ab8565732c59a302,
    256'h329925186604edbd5029a9f865268e90003b5b69d3e99240c3432291a60c62a4,
    256'hebad1ed028cd021b27260db22089e0c44481b1a4c120134ac63dc52fbc4cafb2,
    256'he065add2665fb361665267b53024329d96587d661f724171155ee73a3f0c47a8,
    256'h149751a5903c8bbcaf1782e415dfda531eb2af67c25e190330a12000e1fbb9cd
  };

  // These LFSR parameters have been generated with
  // $ ./util/design/gen-lfsr-seed.py --width 32 --seed 2336700764 --prefix ""
  parameter int LfsrFwdWidth = 32;
  typedef logic [LfsrFwdWidth-1:0][$clog2(LfsrFwdWidth)-1:0] lfsr_fwd_perm_t;
  parameter lfsr_fwd_perm_t RndCnstLfsrFwdPermDefault = {
    160'h7f3ac6d173d78678d84908157fba482e76685704
  };

  // Message permutation
  // These LFSR parameters have been generated with
  // $ ./util/design/gen-lfsr-seed.py --width 64 --seed 1201202158 --prefix ""
  // And changed the type name from lfsr_perm_t to msg_perm_t
  typedef logic [MsgWidth-1:0][$clog2(MsgWidth)-1:0] msg_perm_t;
  parameter msg_perm_t RndCnstMsgPermDefault = {
    128'h382af41849db4cfb9c885f72f118c102,
    256'hcb5526978defac799192f65f54148379af21d7e10d82a5a33c3f31a1eaf964b8
  };

  ///////////////////////////
  // Application interface //
  ///////////////////////////

  // Number of the application interface
  // Currently KMAC has three interface.
  // 0: KeyMgr
  // 1: LC_CTRL
  // 2: ROM_CTRL
  // Make sure to change `width` of app inter-module signal definition
  // if this value is changed.
  parameter int unsigned NumAppIntf = 3;

  // Application Algorithm
  // Each interface can choose algorithms among SHA3, cSHAKE, KMAC
  typedef enum bit [1:0] {
    // SHA3 mode doer not nees any additional information.
    // Prefix will be tied to all zero and not used.
    AppSHA3   = 0,

    // In CShake/ KMAC mode, the Prefix can be determined by the compile-time
    // parameter or through CSRs.
    AppCShake = 1,

    // In KMAC mode, the secret key always comes from sideload.
    // KMAC mode needs uniformly distributed entropy. The request will be
    // silently discarded in Reset state.
    AppKMAC   = 2
  } app_mode_e;

  // Predefined encoded_string
  parameter logic [15:0] EncodedStringEmpty   = 16'h                     0001;
  parameter logic [47:0] EncodedStringKMAC    = 48'h           4341_4D4B_2001;
  // encoded_string("LC_CTRL")
  parameter logic [71:0] EncodedStringLcCtrl  = 72'h   4c_5254_435f_434C_3801;
  // encoded_string("ROM_CTRL")
  parameter logic [79:0] EncodedStringRomCtrl = 80'h 4c52_5443_5f4d_4f52_4001;
  parameter int unsigned NSPrefixW = sha3_pkg::NSRegisterSize*8;

  typedef struct packed {
    app_mode_e Mode;

    sha3_pkg::keccak_strength_e Strength;

    // PrefixMode determines the origin value of Prefix that is used in KMAC
    // and cSHAKE operations.
    // Choose **0** for CSRs (!!PREFIX), or **1** to use `Prefix` parameter
    // below.
    bit PrefixMode;

    // If `PrefixMode` is 1'b 1, then this `Prefix` value will be used in
    // cSHAKE or KMAC operation.
    logic [NSPrefixW-1:0] Prefix;
  } app_config_t;

  parameter app_config_t AppCfg [NumAppIntf] = '{
    // KeyMgr
    '{
      Mode:       AppKMAC, // KeyMgr uses KMAC operation
      Strength:   sha3_pkg::L256,
      PrefixMode: 1'b 1,   // Use prefix parameter
      // {fname: encoded_string("KMAC"), custom_str: encoded_string("")}
      Prefix:     NSPrefixW'({EncodedStringEmpty, EncodedStringKMAC})
    },

    // LC_CTRL
    '{
      Mode:       AppCShake,
      Strength:   sha3_pkg::L128,
      PrefixMode: 1'b 1,     // Use prefix parameter
      // {fname: encode_string(""), custom_str: encode_string("LC_CTRL")}
      Prefix: NSPrefixW'({EncodedStringLcCtrl, EncodedStringEmpty})
    },

    // ROM_CTRL
    '{
      Mode:       AppCShake,
      Strength:   sha3_pkg::L256,
      PrefixMode: 1'b 1,     // Use prefix parameter
      // {fname: encode_string(""), custom_str: encode_string("ROM_CTRL")}
      Prefix: NSPrefixW'({EncodedStringRomCtrl, EncodedStringEmpty})
    }
  };

  // Exporting the app internal mux selection enum into the package. So that DV
  // can use this enum in its scoreboard.
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 4 -n 5 \
  //      -s 713832113 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (66.67%)
  //  4: |||||||||| (33.33%)
  //  5: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4
  //
  localparam int AppMuxWidth = 5;
  typedef enum logic [AppMuxWidth-1:0] {
    SelNone   = 5'b10100,
    SelApp    = 5'b11001,
    SelOutLen = 5'b00010,
    SelSw     = 5'b01111
  } app_mux_sel_e ;



  // MsgWidth : 64
  // MsgStrbW : 8
  parameter int unsigned AppDigestW = 384;
  parameter int unsigned AppKeyW = 256;

  typedef struct packed {
    logic valid;
    logic [MsgWidth-1:0] data;
    logic [MsgStrbW-1:0] strb;
    logic last;
  } app_req_t;

  typedef struct packed {
    logic ready;
    logic done;
    logic [AppDigestW-1:0] digest_share0;
    logic [AppDigestW-1:0] digest_share1;
    // Error is valid when done is high. If any error occurs during KDF, KMAC
    // returns the garbage digest data with error. The KeyMgr discards the
    // digest and may re-initiate the process.
    logic error;
  } app_rsp_t;

  parameter app_req_t APP_REQ_DEFAULT = '{
    valid: 1'b 0,
    data: '0,
    strb: '0,
    last: 1'b 0
  };
  parameter app_rsp_t APP_RSP_DEFAULT = '{
    ready: 1'b1,
    done:  1'b1,
    digest_share0: AppDigestW'(32'hDEADBEEF),
    digest_share1: AppDigestW'(32'hFACEBEEF),
    error: 1'b1
  };


  ////////////////////
  // Error Handling //
  ////////////////////

  // Error structure is same to the SHA3 one. The codes do not overlap.
  typedef enum logic [7:0] {
    ErrNone = 8'h 00,

    // ErrSha3SwControl occurs when software sent wrong flow signal.
    // e.g) Sw set `process_i` without `start_i`. The state machine ignores
    //      the signal and report through the error FIFO.
    //ErrSha3SwControl = 8'h 80

    // ErrKeyNotValid: KeyMgr interface raises an error if the secret key is
    // not valid when KeyMgr initiates KDF.
    ErrKeyNotValid = 8'h 01,

    // ErrSwPushMsgFifo: Sw writes data into Msg FIFO abruptly.
    // This error occurs in below scenario:
    //   - Sw does not send "Start" command to KMAC then writes data into
    //     Msg FIFO
    //   - Sw writes data into Msg FIFO when KeyMgr is in operation
    ErrSwPushedMsgFifo = 8'h 02,

    // ErrSwIssuedCmdInAppActive
    //  - Sw writes any command while AppIntf is in active.
    ErrSwIssuedCmdInAppActive = 8'h 03,

    // ErrWaitTimerExpired
    // Entropy Wait timer expired. Something wrong on EDN i/f
    ErrWaitTimerExpired = 8'h 04,

    // ErrIncorrectEntropyMode
    // Incorrect Entropy mode when entropy is ready
    ErrIncorrectEntropyMode = 8'h 05,

    // ErrUnexpectedModeStrength
    ErrUnexpectedModeStrength = 8'h 06,

    // ErrIncorrectFunctionName "KMAC"
    ErrIncorrectFunctionName = 8'h 07,

    // ErrSwCmdSequence
    ErrSwCmdSequence = 8'h 08,

    // ErrSwHashingWithoutEntropyReady
    //  - Sw issues KMAC op without Entropy setting.
    ErrSwHashingWithoutEntropyReady = 8'h 09,

    // Error Shadow register update
    ErrShadowRegUpdate = 8'h C0,

    // Error due to lc_escalation_en_i or fatal fault
    ErrFatalError = 8'h C1,

    // Error due to the counter integrity check failure inside MsgFifo.Packer
    ErrPackerIntegrity = 8'h C2,

    // Error due to the counter integrity check failure inside MsgFifo.Fifo
    ErrMsgFifoIntegrity = 8'h C3
  } err_code_e;

  typedef struct packed {
    logic        valid;
    err_code_e   code; // Type of error
    logic [23:0] info; // Additional Debug info
  } err_t;
  parameter int unsigned ErrInfoW = 24 ; // err_t::info

  typedef struct packed {
    logic [AppDigestW-1:0] digest_share0;
    logic [AppDigestW-1:0] digest_share1;
  } rsp_digest_t;
  ///////////////////////
  // Library Functions //
  ///////////////////////

  // Endian conversion functions (32-bit, 64-bit)
  function automatic logic [31:0] conv_endian32( input logic [31:0] v, input logic swap);
    logic [31:0] conv_data = {<<8{v}};
    conv_endian32 = (swap) ? conv_data : v ;
  endfunction : conv_endian32

  function automatic logic [63:0] conv_endian64( input logic [63:0] v, input logic swap);
    logic [63:0] conv_data = {<<8{v}};
    conv_endian64 = (swap) ? conv_data : v ;
  endfunction : conv_endian64

endpackage : kmac_pkg


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager top level
//

`include "prim_assert.sv"

module keymgr
  import keymgr_pkg::*;
  import keymgr_reg_pkg::*;
#(
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},
  parameter bit KmacEnMasking                  = 1'b1,
  parameter lfsr_seed_t RndCnstLfsrSeed        = RndCnstLfsrSeedDefault,
  parameter lfsr_perm_t RndCnstLfsrPerm        = RndCnstLfsrPermDefault,
  parameter rand_perm_t RndCnstRandPerm        = RndCnstRandPermDefault,
  parameter seed_t RndCnstRevisionSeed         = RndCnstRevisionSeedDefault,
  parameter seed_t RndCnstCreatorIdentitySeed  = RndCnstCreatorIdentitySeedDefault,
  parameter seed_t RndCnstOwnerIntIdentitySeed = RndCnstOwnerIntIdentitySeedDefault,
  parameter seed_t RndCnstOwnerIdentitySeed    = RndCnstOwnerIdentitySeedDefault,
  parameter seed_t RndCnstSoftOutputSeed       = RndCnstSoftOutputSeedDefault,
  parameter seed_t RndCnstHardOutputSeed       = RndCnstHardOutputSeedDefault,
  parameter seed_t RndCnstNoneSeed             = RndCnstNoneSeedDefault,
  parameter seed_t RndCnstAesSeed              = RndCnstAesSeedDefault,
  parameter seed_t RndCnstOtbnSeed             = RndCnstOtbnSeedDefault,
  parameter seed_t RndCnstKmacSeed             = RndCnstKmacSeedDefault,
  parameter seed_t RndCnstCdi                  = RndCnstCdiDefault
) (
  input clk_i,
  input rst_ni,
  input rst_shadowed_ni,
  input clk_edn_i,
  input rst_edn_ni,

  // Bus Interface
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // key interface to crypto modules
  output hw_key_req_t aes_key_o,
  output hw_key_req_t kmac_key_o,
  output otbn_key_req_t otbn_key_o,

  // data interface to/from crypto modules
  output kmac_pkg::app_req_t kmac_data_o,
  input  kmac_pkg::app_rsp_t kmac_data_i,

  // whether kmac is masked
  // Note this input is not driving ANY logic directly.  Instead it is only used
  // as part of assertions.  This is done because if boundary optimization were
  // ever disabled, it would provide a VERY obvious location for attacks.
  input kmac_en_masking_i,

  // the following signals should eventually be wrapped into structs from other modules
  // SEC_CM: LC_CTRL.INTERSIG.MUBI
  input lc_ctrl_pkg::lc_tx_t lc_keymgr_en_i,
  input lc_ctrl_pkg::lc_keymgr_div_t lc_keymgr_div_i,
  input otp_ctrl_pkg::otp_keymgr_key_t otp_key_i,
  input otp_ctrl_pkg::otp_device_id_t otp_device_id_i,
  input flash_ctrl_pkg::keymgr_flash_t flash_i,

  // connection to edn
  output edn_pkg::edn_req_t edn_o,
  input edn_pkg::edn_rsp_t edn_i,

  // connection to rom_ctrl
  input rom_ctrl_pkg::keymgr_data_t rom_digest_i,

  // interrupts and alerts
  output logic intr_op_done_o,
  input  prim_alert_pkg::alert_rx_t [keymgr_reg_pkg::NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [keymgr_reg_pkg::NumAlerts-1:0] alert_tx_o
);

  `ASSERT_INIT(AdvDataWidth_A, AdvDataWidth <= KDFMaxWidth)
  `ASSERT_INIT(IdDataWidth_A,  IdDataWidth  <= KDFMaxWidth)
  `ASSERT_INIT(GenDataWidth_A, GenDataWidth <= KDFMaxWidth)
  `ASSERT_INIT(OutputKeyDiff_A, RndCnstHardOutputSeed != RndCnstSoftOutputSeed)

  import prim_mubi_pkg::mubi4_test_true_strict;
  import prim_mubi_pkg::mubi4_test_false_strict;

  /////////////////////////////////////
  // Anchor incoming seeds and constants
  /////////////////////////////////////
  localparam int TotalSeedWidth = KeyWidth * 10;
  seed_t revision_seed;
  seed_t creator_identity_seed;
  seed_t owner_int_identity_seed;
  seed_t owner_identity_seed;
  seed_t soft_output_seed;
  seed_t hard_output_seed;
  seed_t aes_seed;
  seed_t otbn_seed;
  seed_t kmac_seed;
  seed_t none_seed;

  prim_sec_anchor_buf #(
    .Width(TotalSeedWidth)
  ) u_seed_anchor (
    .in_i({RndCnstRevisionSeed,
           RndCnstCreatorIdentitySeed,
           RndCnstOwnerIntIdentitySeed,
           RndCnstOwnerIdentitySeed,
           RndCnstSoftOutputSeed,
           RndCnstHardOutputSeed,
           RndCnstAesSeed,
           RndCnstOtbnSeed,
           RndCnstKmacSeed,
           RndCnstNoneSeed}),
    .out_o({revision_seed,
            creator_identity_seed,
            owner_int_identity_seed,
            owner_identity_seed,
            soft_output_seed,
            hard_output_seed,
            aes_seed,
            otbn_seed,
            kmac_seed,
            none_seed})
  );

  // Register module
  keymgr_reg2hw_t reg2hw;
  keymgr_hw2reg_t hw2reg;

  logic regfile_intg_err;
  logic shadowed_storage_err;
  logic shadowed_update_err;
  // SEC_CM: BUS.INTEGRITY
  // SEC_CM: CONFIG.SHADOW
  // SEC_CM: OP.CONFIG.REGWEN, RESEED.CONFIG.REGWEN, SW_BINDING.CONFIG.REGWEN
  // SEC_CM: MAX_KEY_VER.CONFIG.REGWEN
  keymgr_reg_top u_reg (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,
    .tl_i,
    .tl_o,
    .reg2hw,
    .hw2reg,
    .shadowed_storage_err_o (shadowed_storage_err),
    .shadowed_update_err_o  (shadowed_update_err),
    .intg_err_o             (regfile_intg_err),

    .devmode_i (1'b1) // connect to real devmode signal in the future
  );

  /////////////////////////////////////
  //  Synchronize lc_ctrl control inputs
  //  Data inputs are not synchronized and assumed quasi-static
  /////////////////////////////////////
  lc_ctrl_pkg::lc_tx_t [KeyMgrEnLast-1:0] lc_keymgr_en;

  prim_lc_sync #(
    .NumCopies(int'(KeyMgrEnLast))
  ) u_lc_keymgr_en_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i(lc_keymgr_en_i),
    .lc_en_o(lc_keymgr_en)
  );


  /////////////////////////////////////
  //  LFSR
  /////////////////////////////////////

  // A farily large lfsr is used here as entropy in multiple places.
  // - populate the default working state
  // - generate random inputs when a bad input is selected
  //
  // The first case is sensitive, and thus the working state is constructed
  // through multiple rounds of the Lfsr
  // The second case is less sensitive and is applied directly.  If the inputs
  // have more bits than the lfsr output, the lfsr value is simply replicated

  logic seed_en;
  logic [LfsrWidth-1:0] seed;
  logic reseed_req;
  logic reseed_ack;
  logic reseed_cnt_err;

  keymgr_reseed_ctrl u_reseed_ctrl (
    .clk_i,
    .rst_ni,
    .clk_edn_i,
    .rst_edn_ni,
    .reseed_req_i(reseed_req),
    .reseed_ack_o(reseed_ack),
    .reseed_interval_i(reg2hw.reseed_interval_shadowed.q),
    .edn_o,
    .edn_i,
    .seed_en_o(seed_en),
    .seed_o(seed),
    .cnt_err_o(reseed_cnt_err)
  );

  logic [63:0] lfsr;
  logic ctrl_lfsr_en, data_lfsr_en, sideload_lfsr_en;

  prim_lfsr #(
    .LfsrDw(LfsrWidth),
    .StateOutDw(LfsrWidth),
    .DefaultSeed(RndCnstLfsrSeed),
    .StatePermEn(1'b1),
    .StatePerm(RndCnstLfsrPerm),
    .NonLinearOut(1'b1)
  ) u_lfsr (
    .clk_i,
    .rst_ni,
    .lfsr_en_i(ctrl_lfsr_en | data_lfsr_en | sideload_lfsr_en),
    // The seed update is skipped if there is an ongoing keymgr transaction.
    // This is not really done for any functional purpose but more to simplify
    // DV. When an invalid operation is selected, the keymgr just starts transmitting
    // whatever is at the prng output, however, this may cause a dv protocol violation
    // if a reseed happens to coincide.
    .seed_en_i(seed_en & ~reg2hw.start.q),
    .seed_i(seed),
    .entropy_i('0),
    .state_o(lfsr)
  );
  `ASSERT_INIT(LfsrWidth_A, LfsrWidth == 64)


  logic [Shares-1:0][RandWidth-1:0] ctrl_rand;
  logic [Shares-1:0][RandWidth-1:0] data_rand;

  assign ctrl_rand[0] = lfsr[63:32];
  assign ctrl_rand[1] = perm_data(lfsr[31:0], RndCnstRandPerm);

  assign data_rand[0] = lfsr[31:0];
  assign data_rand[1] = perm_data(lfsr[63:32], RndCnstRandPerm);

  /////////////////////////////////////
  //  Key Manager Control
  /////////////////////////////////////

  keymgr_stage_e stage_sel;
  logic invalid_stage_sel;
  prim_mubi_pkg::mubi4_t hw_key_sel;
  logic adv_en, id_en, gen_en;
  logic wipe_key;
  hw_key_req_t kmac_key;
  logic op_done;
  logic init;
  logic data_valid;
  logic data_hw_en;
  logic data_sw_en;
  logic kmac_done;
  logic kmac_input_invalid;
  logic kmac_cmd_err;
  logic kmac_fsm_err;
  logic kmac_op_err;
  logic kmac_done_err;
  logic [Shares-1:0][kmac_pkg::AppDigestW-1:0] kmac_data;
  logic [Shares-1:0][KeyWidth-1:0] kmac_data_truncated;
  logic [ErrLastPos-1:0] err_code;
  logic [FaultLastPos-1:0] fault_code;
  logic sw_binding_unlock;
  logic [CdiWidth-1:0] cdi_sel;
  logic sideload_fsm_err;
  logic sideload_sel_err;

  for (genvar i = 0; i < Shares; i++) begin : gen_truncate_data
    assign kmac_data_truncated[i] = kmac_data[i][KeyWidth-1:0];
  end

  logic op_start;
  assign op_start = reg2hw.start.q;
  keymgr_ctrl #(
    .KmacEnMasking(KmacEnMasking)
  ) u_ctrl (
    .clk_i,
    .rst_ni,
    .en_i(lc_keymgr_en[KeyMgrEnCtrl] == lc_ctrl_pkg::On),
    .regfile_intg_err_i(regfile_intg_err),
    .shadowed_update_err_i(shadowed_update_err),
    .shadowed_storage_err_i(shadowed_storage_err),
    .reseed_cnt_err_i(reseed_cnt_err),
    .sideload_sel_err_i(sideload_sel_err),
    .sideload_fsm_err_i(sideload_fsm_err),
    .prng_reseed_req_o(reseed_req),
    .prng_reseed_ack_i(reseed_ack),
    .prng_en_o(ctrl_lfsr_en),
    .entropy_i(ctrl_rand),
    .op_i(keymgr_ops_e'(reg2hw.control_shadowed.operation.q)),
    .op_start_i(op_start),
    .op_cdi_sel_i(reg2hw.control_shadowed.cdi_sel.q),
    .op_done_o(op_done),
    .init_o(init),
    .sw_binding_unlock_o(sw_binding_unlock),
    .status_o(hw2reg.op_status.d),
    .fault_o(fault_code),
    .error_o(err_code),
    .data_hw_en_o(data_hw_en),
    .data_sw_en_o(data_sw_en),
    .data_valid_o(data_valid),
    .working_state_o(hw2reg.working_state.d),
    .root_key_i(otp_key_i),
    .hw_sel_o(hw_key_sel),
    .stage_sel_o(stage_sel),
    .invalid_stage_sel_o(invalid_stage_sel),
    .cdi_sel_o(cdi_sel),
    .wipe_key_o(wipe_key),
    .adv_en_o(adv_en),
    .id_en_o(id_en),
    .gen_en_o(gen_en),
    .key_o(kmac_key),
    .kmac_done_i(kmac_done),
    .kmac_input_invalid_i(kmac_input_invalid),
    .kmac_fsm_err_i(kmac_fsm_err),
    .kmac_op_err_i(kmac_op_err),
    .kmac_done_err_i(kmac_done_err),
    .kmac_cmd_err_i(kmac_cmd_err),
    .kmac_data_i(kmac_data_truncated)
  );

  assign hw2reg.start.d  = '0;
  assign hw2reg.start.de = op_done;
  // as long as operation is ongoing, capture status
  assign hw2reg.op_status.de = op_start;

  // working state is always visible
  assign hw2reg.working_state.de = 1'b1;

  logic cfg_regwen;

  // key manager registers cannot be changed once an operation starts
  keymgr_cfg_en u_cfgen (
    .clk_i,
    .rst_ni,
    .init_i(1'b1), // cfg_regwen does not care about init
    .en_i(lc_keymgr_en[KeyMgrEnCfgEn] == lc_ctrl_pkg::On),
    .set_i(op_start & op_done),
    .clr_i(op_start),
    .out_o(cfg_regwen)
  );

  assign hw2reg.cfg_regwen.d = cfg_regwen;


  logic sw_binding_clr;
  logic sw_binding_regwen;

  // this is w0c
  assign sw_binding_clr = reg2hw.sw_binding_regwen.qe & ~reg2hw.sw_binding_regwen.q;

  // software clears the enable
  // hardware restores it upon successful advance
  keymgr_cfg_en #(
    .NonInitClr(1'b1)  // clear has an effect regardless of init state
  ) u_sw_binding_regwen (
    .clk_i,
    .rst_ni,
    .init_i(init),
    .en_i(lc_keymgr_en[KeyMgrEnSwBindingEn] == lc_ctrl_pkg::On),
    .set_i(sw_binding_unlock),
    .clr_i(sw_binding_clr),
    .out_o(sw_binding_regwen)
  );

  assign hw2reg.sw_binding_regwen.d = sw_binding_regwen & cfg_regwen;

  /////////////////////////////////////
  //  Key Manager Input Construction
  /////////////////////////////////////

  // The various arrays of inputs for each operation
  logic rom_digest_vld;
  logic [2**StageWidth-1:0][AdvDataWidth-1:0] adv_matrix;
  logic [2**StageWidth-1:0] adv_dvalid;
  logic [2**StageWidth-1:0][IdDataWidth-1:0] id_matrix;
  logic [GenDataWidth-1:0] gen_in;

  // The max key version for each stage
  logic [2**StageWidth-1:0][31:0] max_key_versions;

  // Number of times the lfsr output fits into the inputs
  localparam int AdvLfsrCopies = AdvDataWidth / 32;
  localparam int IdLfsrCopies = IdDataWidth / 32;
  localparam int GenLfsrCopies = GenDataWidth / 32;

  // input checking
  logic creator_seed_vld;
  logic owner_seed_vld;
  logic devid_vld;
  logic health_state_vld;
  logic key_version_vld;

  // software binding
  logic [SwBindingWidth-1:0] sw_binding;
  assign sw_binding = (cdi_sel == 0) ? reg2hw.sealing_sw_binding :
                      (cdi_sel == 1) ? reg2hw.attest_sw_binding  : RndCnstCdi;

  // Advance state operation input construction
  for (genvar i = KeyMgrStages; i < 2**StageWidth; i++) begin : gen_adv_matrix_fill
    assign adv_matrix[i] = {AdvLfsrCopies{data_rand[0]}};
    assign adv_dvalid[i] = 1'b1;
  end

  // Advance to creator_root_key
  // The values coming from otp_ctrl / lc_ctrl are treat as quasi-static for CDC purposes
  logic [KeyWidth-1:0] creator_seed;
  assign creator_seed = flash_i.seeds[flash_ctrl_pkg::CreatorSeedIdx];
  assign adv_matrix[Creator] = AdvDataWidth'({sw_binding,
                                              revision_seed,
                                              otp_device_id_i,
                                              lc_keymgr_div_i,
                                              rom_digest_i.data,
                                              creator_seed});

  assign adv_dvalid[Creator] = creator_seed_vld &
                               devid_vld &
                               health_state_vld &
                               rom_digest_vld;

  // Advance to owner_intermediate_key
  logic [KeyWidth-1:0] owner_seed;
  assign owner_seed = flash_i.seeds[flash_ctrl_pkg::OwnerSeedIdx];
  assign adv_matrix[OwnerInt] = AdvDataWidth'({sw_binding,owner_seed});
  assign adv_dvalid[OwnerInt] = owner_seed_vld;

  // Advance to owner_key
  assign adv_matrix[Owner] = AdvDataWidth'(sw_binding);
  assign adv_dvalid[Owner] = 1'b1;

  // Generate Identity operation input construction
  for (genvar i = KeyMgrStages; i < 2**StageWidth; i++) begin : gen_id_matrix_fill
    assign id_matrix[i] = {IdLfsrCopies{data_rand[0]}};
  end

  assign id_matrix[Creator]  = creator_identity_seed;
  assign id_matrix[OwnerInt] = owner_int_identity_seed;
  assign id_matrix[Owner]    = owner_identity_seed;


  // Generate output operation input construction
  logic [KeyWidth-1:0] output_key;
  keymgr_key_dest_e dest_sel;
  logic [KeyWidth-1:0] dest_seed;

  assign dest_sel = keymgr_key_dest_e'(reg2hw.control_shadowed.dest_sel.q);
  assign dest_seed = dest_sel == Aes  ? aes_seed  :
                       dest_sel == Kmac ? kmac_seed :
                       dest_sel == Otbn ? otbn_seed : none_seed;
  assign output_key = mubi4_test_true_strict(hw_key_sel) ? hard_output_seed :
                      soft_output_seed;
  assign gen_in = invalid_stage_sel ? {GenLfsrCopies{lfsr[31:0]}} : {reg2hw.key_version,
                                                                     reg2hw.salt,
                                                                     dest_seed,
                                                                     output_key};

  // Advance state operation input construction
  for (genvar i = KeyMgrStages; i < 2**StageWidth; i++) begin : gen_key_version_fill
    assign max_key_versions[i] = '0;
  end

  assign max_key_versions[Creator]  = reg2hw.max_creator_key_ver_shadowed.q;
  assign max_key_versions[OwnerInt] = reg2hw.max_owner_int_key_ver_shadowed.q;
  assign max_key_versions[Owner]    = reg2hw.max_owner_key_ver_shadowed.q;


  // General module for checking inputs
  logic key_vld;
  // SEC_CM: CONSTANTS.CONSISTENCY
  // SEC_CM: INTERSIG.CONSISTENCY
  keymgr_input_checks #(
    .KmacEnMasking(KmacEnMasking)
  ) u_checks (
    .rom_digest_i,
    .max_key_versions_i(max_key_versions),
    .stage_sel_i(stage_sel),
    .key_version_i(reg2hw.key_version),
    .creator_seed_i(creator_seed),
    .owner_seed_i(owner_seed),
    .key_i(kmac_key_o),
    .devid_i(otp_device_id_i),
    .health_state_i(HealthStateWidth'(lc_keymgr_div_i)),
    .creator_seed_vld_o(creator_seed_vld),
    .owner_seed_vld_o(owner_seed_vld),
    .devid_vld_o(devid_vld),
    .health_state_vld_o(health_state_vld),
    .key_version_vld_o(key_version_vld),
    .key_vld_o(key_vld),
    .rom_digest_vld_o(rom_digest_vld)
  );

  assign hw2reg.debug.invalid_creator_seed.d = 1'b1;
  assign hw2reg.debug.invalid_owner_seed.d = 1'b1;
  assign hw2reg.debug.invalid_dev_id.d = 1'b1;
  assign hw2reg.debug.invalid_health_state.d = 1'b1;
  assign hw2reg.debug.invalid_key_version.d = 1'b1;
  assign hw2reg.debug.invalid_key.d = 1'b1;
  assign hw2reg.debug.invalid_digest.d = 1'b1;

  logic valid_op;
  assign valid_op = adv_en | id_en | gen_en;
  assign hw2reg.debug.invalid_creator_seed.de = adv_en & (stage_sel == Creator) & ~creator_seed_vld;
  assign hw2reg.debug.invalid_owner_seed.de = adv_en & (stage_sel == OwnerInt) & ~owner_seed_vld;
  assign hw2reg.debug.invalid_dev_id.de = adv_en & (stage_sel == Creator) & ~devid_vld;
  assign hw2reg.debug.invalid_health_state.de = adv_en & (stage_sel == Creator) & ~health_state_vld;
  assign hw2reg.debug.invalid_key_version.de = gen_en & ~key_version_vld;
  assign hw2reg.debug.invalid_key.de = valid_op & ~key_vld;
  assign hw2reg.debug.invalid_digest.de = adv_en & (stage_sel == Creator) & ~rom_digest_vld;

  /////////////////////////////////////
  //  KMAC Control
  /////////////////////////////////////

  logic [3:0] invalid_data;
  assign invalid_data[OpAdvance]  = ~key_vld | ~adv_dvalid[stage_sel];
  assign invalid_data[OpGenId]    = ~key_vld;
  assign invalid_data[OpGenSwOut] = ~key_vld | ~key_version_vld;
  assign invalid_data[OpGenHwOut] = ~key_vld | ~key_version_vld;

  keymgr_kmac_if u_kmac_if (
    .clk_i,
    .rst_ni,
    .prng_en_o(data_lfsr_en),
    .adv_data_i(adv_matrix[stage_sel]),
    .id_data_i(id_matrix[stage_sel]),
    .gen_data_i(gen_in),
    .inputs_invalid_i(invalid_data),
    .inputs_invalid_o(kmac_input_invalid),
    .adv_en_i(adv_en),
    .id_en_i(id_en),
    .gen_en_i(gen_en),
    .done_o(kmac_done),
    .data_o(kmac_data),
    .kmac_data_o,
    .kmac_data_i,
    .entropy_i(data_rand),
    .fsm_error_o(kmac_fsm_err),
    .kmac_error_o(kmac_op_err),
    .kmac_done_error_o(kmac_done_err),
    .cmd_error_o(kmac_cmd_err)
  );


  /////////////////////////////////////
  //  Side load key storage
  /////////////////////////////////////
  // SEC_CM: HW.KEY.SW_NOACCESS
  keymgr_sideload_key_ctrl u_sideload_ctrl (
    .clk_i,
    .rst_ni,
    .init_i(init),
    .entropy_i(data_rand),
    .clr_key_i(keymgr_sideload_clr_e'(reg2hw.sideload_clear.q)),
    .wipe_key_i(wipe_key),
    .dest_sel_i(dest_sel),
    .hw_key_sel_i(hw_key_sel),
    // SEC_CM: OUTPUT_KEYS.CTRL.REDUN
    .data_en_i(data_hw_en),
    .data_valid_i(data_valid),
    .key_i(kmac_key),
    .data_i(kmac_data),
    .prng_en_o(sideload_lfsr_en),
    .aes_key_o,
    .otbn_key_o,
    .kmac_key_o,
    .sideload_sel_err_o(sideload_sel_err),
    .fsm_err_o(sideload_fsm_err)
  );

  for (genvar i = 0; i < 8; i++) begin : gen_sw_assigns

    prim_mubi_pkg::mubi4_t [1:0] hw_key_sel_buf;
    prim_mubi4_sync #(
      .NumCopies(2),
      .AsyncOn(0)
    ) u_mubi_buf (
      .clk_i,
      .rst_ni,
      .mubi_i(hw_key_sel),
      .mubi_o(hw_key_sel_buf)
    );

    // SEC_CM: OUTPUT_KEYS.CTRL.REDUN
    prim_sec_anchor_buf #(
     .Width(32)
    ) u_prim_buf_share0_d (
      .in_i(~data_sw_en | wipe_key ? data_rand[0] : kmac_data[0][i*32 +: 32]),
      .out_o(hw2reg.sw_share0_output[i].d)
    );

    prim_sec_anchor_buf #(
     .Width(32)
    ) u_prim_buf_share1_d (
      .in_i(~data_sw_en | wipe_key ? data_rand[1] : kmac_data[1][i*32 +: 32]),
      .out_o(hw2reg.sw_share1_output[i].d)
    );

    prim_sec_anchor_buf #(
     .Width(1)
    ) u_prim_buf_share0_de (
      .in_i(wipe_key | data_valid & mubi4_test_false_strict(hw_key_sel_buf[0])),
      .out_o(hw2reg.sw_share0_output[i].de)
    );

    prim_sec_anchor_buf #(
     .Width(1)
    ) u_prim_buf_share1_de (
      .in_i(wipe_key | data_valid & mubi4_test_false_strict(hw_key_sel_buf[1])),
      .out_o(hw2reg.sw_share1_output[i].de)
    );
  end

  /////////////////////////////////////
  //  Alerts and Interrupts
  /////////////////////////////////////

  prim_intr_hw #(.Width(1)) u_intr_op_done (
    .clk_i,
    .rst_ni,
    .event_intr_i           (op_done),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.d),
    .intr_o                 (intr_op_done_o)
  );

  assign hw2reg.err_code.invalid_op.d             = 1'b1;
  assign hw2reg.err_code.invalid_kmac_input.d     = 1'b1;
  assign hw2reg.err_code.invalid_shadow_update.d  = 1'b1;
  assign hw2reg.err_code.invalid_op.de            = err_code[ErrInvalidOp];
  assign hw2reg.err_code.invalid_kmac_input.de    = err_code[ErrInvalidIn];
  assign hw2reg.err_code.invalid_shadow_update.de = err_code[ErrShadowUpdate];

  assign hw2reg.fault_status.cmd.de           = fault_code[FaultKmacCmd];
  assign hw2reg.fault_status.kmac_fsm.de      = fault_code[FaultKmacFsm];
  assign hw2reg.fault_status.kmac_op.de       = fault_code[FaultKmacOp];
  assign hw2reg.fault_status.kmac_done.de     = fault_code[FaultKmacDone];
  assign hw2reg.fault_status.kmac_out.de      = fault_code[FaultKmacOut];
  assign hw2reg.fault_status.regfile_intg.de  = fault_code[FaultRegIntg];
  assign hw2reg.fault_status.shadow.de        = fault_code[FaultShadow];
  assign hw2reg.fault_status.ctrl_fsm_intg.de = fault_code[FaultCtrlFsm];
  assign hw2reg.fault_status.ctrl_fsm_chk.de  = fault_code[FaultCtrlFsmChk];
  assign hw2reg.fault_status.ctrl_fsm_cnt.de  = fault_code[FaultCtrlCnt];
  assign hw2reg.fault_status.reseed_cnt.de    = fault_code[FaultReseedCnt];
  assign hw2reg.fault_status.side_ctrl_fsm.de = fault_code[FaultSideFsm];
  assign hw2reg.fault_status.side_ctrl_sel.de = fault_code[FaultSideSel];
  assign hw2reg.fault_status.key_ecc.de       = fault_code[FaultKeyEcc];
  assign hw2reg.fault_status.cmd.d            = 1'b1;
  assign hw2reg.fault_status.kmac_fsm.d       = 1'b1;
  assign hw2reg.fault_status.kmac_done.d      = 1'b1;
  assign hw2reg.fault_status.kmac_op.d        = 1'b1;
  assign hw2reg.fault_status.kmac_out.d       = 1'b1;
  assign hw2reg.fault_status.regfile_intg.d   = 1'b1;
  assign hw2reg.fault_status.shadow.d         = 1'b1;
  assign hw2reg.fault_status.ctrl_fsm_intg.d  = 1'b1;
  assign hw2reg.fault_status.ctrl_fsm_chk.d   = 1'b1;
  assign hw2reg.fault_status.ctrl_fsm_cnt.d   = 1'b1;
  assign hw2reg.fault_status.reseed_cnt.d     = 1'b1;
  assign hw2reg.fault_status.side_ctrl_fsm.d  = 1'b1;
  assign hw2reg.fault_status.side_ctrl_sel.d  = 1'b1;
  assign hw2reg.fault_status.key_ecc.d        = 1'b1;

  // There are two types of alerts
  // - alerts for hardware errors, these could not have been generated by software.
  // - alerts for errors that may have been generated by software.

  logic fault_errs, fault_err_req_q, fault_err_req_d, fault_err_ack;
  logic op_errs, op_err_req_q, op_err_req_d, op_err_ack;

  // Fault status can happen independently of any operation
  assign fault_errs = |reg2hw.fault_status;

  assign fault_err_req_d = fault_errs    ? 1'b1 :
                           fault_err_ack ? 1'b0 : fault_err_req_q;

  assign op_errs = |err_code;
  assign op_err_req_d = op_errs    ? 1'b1 :
                        op_err_ack ? 1'b0 : op_err_req_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      fault_err_req_q <= '0;
      op_err_req_q <= '0;
    end else begin
      fault_err_req_q <= fault_err_req_d;
      op_err_req_q <= op_err_req_d;
    end
  end

  logic fault_alert_test;
  assign fault_alert_test = reg2hw.alert_test.fatal_fault_err.q &
                            reg2hw.alert_test.fatal_fault_err.qe;
  prim_alert_sender #(
    .AsyncOn(AlertAsyncOn[1]),
    .IsFatal(1)
  ) u_fault_alert (
    .clk_i,
    .rst_ni,
    .alert_test_i(fault_alert_test),
    .alert_req_i(fault_err_req_q),
    .alert_ack_o(fault_err_ack),
    .alert_state_o(),
    .alert_rx_i(alert_rx_i[1]),
    .alert_tx_o(alert_tx_o[1])
  );

  logic op_err_alert_test;
  assign op_err_alert_test = reg2hw.alert_test.recov_operation_err.q &
                             reg2hw.alert_test.recov_operation_err.qe;
  prim_alert_sender #(
    .AsyncOn(AlertAsyncOn[0]),
    .IsFatal(0)
  ) u_op_err_alert (
    .clk_i,
    .rst_ni,
    .alert_test_i(op_err_alert_test),
    .alert_req_i(op_err_req_q),
    .alert_ack_o(op_err_ack),
    .alert_state_o(),
    .alert_rx_i(alert_rx_i[0]),
    .alert_tx_o(alert_tx_o[0])
  );

  // known asserts
  `ASSERT_KNOWN(TlDValidKnownO_A, tl_o.d_valid)
  `ASSERT_KNOWN(TlAReadyKnownO_A, tl_o.a_ready)
  `ASSERT_KNOWN(IntrKnownO_A, intr_op_done_o)
  `ASSERT_KNOWN(AlertKnownO_A, alert_tx_o)

  `ASSERT_KNOWN(AesKeyKnownO_A,  aes_key_o)
  `ASSERT_KNOWN(KmacKeyKnownO_A, kmac_key_o)
  `ASSERT_KNOWN(OtbnKeyKnownO_A, otbn_key_o)
  `ASSERT_KNOWN(KmacDataKnownO_A, kmac_data_o)


  // kmac parameter consistency
  // Both modules must be consistent with regards to masking assumptions
  logic unused_kmac_en_masking;
  assign unused_kmac_en_masking = kmac_en_masking_i;

  `ASSERT_INIT_NET(KmacMaskCheck_A, KmacEnMasking == kmac_en_masking_i)

  // Ensure all parameters are consistent
  `ASSERT_INIT(FaultCntMatch_A, FaultLastPos == AsyncFaultLastIdx + SyncFaultLastIdx)
  `ASSERT_INIT(ErrCntMatch_A, ErrLastPos == AsyncErrLastIdx + SyncErrLastIdx)
  `ASSERT_INIT(StageMatch_A, KeyMgrStages == Disable)

  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CtrlCntAlertCheck_A, u_ctrl.u_cnt, alert_tx_o[1])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(KmacIfCntAlertCheck_A, u_kmac_if.u_cnt, alert_tx_o[1])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(ReseedCtrlCntAlertCheck_A, u_reseed_ctrl.u_reseed_cnt,
                                         alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlMainFsmCheck_A, u_ctrl.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlDataFsmCheck_A,
      u_ctrl.u_data_en.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CtrlOpFsmCheck_A,
      u_ctrl.u_op_state.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(KmacIfFsmCheck_A, u_kmac_if.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(SideloadCtrlFsmCheck_A,
      u_sideload_ctrl.u_state_regs, alert_tx_o[1])

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule // keymgr


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager top level
//

`include "prim_assert.sv"

module keymgr_ctrl
  import keymgr_pkg::*;
  import keymgr_reg_pkg::*;
#(
  parameter bit KmacEnMasking = 1'b1
) (
  input clk_i,
  input rst_ni,

  // lifecycle enforcement
  // SEC_CM: CTRL.FSM.GLOBAL_ESC
  input en_i,

  // faults that can occur outside of operations
  input regfile_intg_err_i,
  input shadowed_update_err_i,
  input shadowed_storage_err_i,
  input reseed_cnt_err_i,
  input sideload_sel_err_i,
  input sideload_fsm_err_i,

  // Software interface
  input op_start_i,
  input keymgr_ops_e op_i,
  input [CdiWidth-1:0] op_cdi_sel_i,
  output logic op_done_o,
  output keymgr_op_status_e status_o,
  output logic [ErrLastPos-1:0] error_o,
  output logic [FaultLastPos-1:0] fault_o,
  output logic data_hw_en_o,
  output logic data_sw_en_o,
  output logic data_valid_o,
  output logic wipe_key_o,
  output keymgr_working_state_e working_state_o,
  output logic sw_binding_unlock_o,
  output logic init_o,

  // Data input
  input  otp_ctrl_pkg::otp_keymgr_key_t root_key_i,
  output prim_mubi_pkg::mubi4_t hw_sel_o,
  output keymgr_stage_e stage_sel_o,
  output logic invalid_stage_sel_o,
  output logic [CdiWidth-1:0] cdi_sel_o,

  // KMAC ctrl interface
  output logic adv_en_o,
  output logic id_en_o,
  output logic gen_en_o,
  output hw_key_req_t key_o,
  input kmac_done_i,
  input kmac_input_invalid_i, // asserted when selected data fails criteria check
  input kmac_fsm_err_i, // asserted when kmac fsm reaches unexpected state
  input kmac_op_err_i,  // asserted when kmac itself reports an error
  input kmac_done_err_i,// asserted when kmac unexpectedly toggles done
  input kmac_cmd_err_i, // asserted when more than one command given to kmac
  input [Shares-1:0][KeyWidth-1:0] kmac_data_i,

  // prng control interface
  input [Shares-1:0][RandWidth-1:0] entropy_i,
  input prng_reseed_ack_i,
  output logic prng_reseed_req_o,
  output logic prng_en_o
);

  localparam int EntropyWidth = LfsrWidth / 2;
  localparam int EntropyRounds = KeyWidth / EntropyWidth;
  localparam int EntropyRndWidth = prim_util_pkg::vbits(EntropyRounds);
  localparam int CntWidth = EntropyRounds > CDIs ? EntropyRndWidth : CdiWidth;
  localparam int EccDataWidth = 64;
  localparam int EccWidth = 8;
  localparam int EccWords = KeyWidth / EccDataWidth;
  localparam int TotalEccWords = EccWords * Shares * CDIs;


  // Enumeration for working state
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 11 -n 10 \
  //      -s 4101887575 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||||||| (54.55%)
  //  6: |||||||||||||||| (45.45%)
  //  7: --
  //  8: --
  //  9: --
  // 10: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 6
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 8
  //
  localparam int StateWidth = 10;
  typedef enum logic [StateWidth-1:0] {
    StCtrlReset          = 10'b1101100001,
    StCtrlEntropyReseed  = 10'b1110010010,
    StCtrlRandom         = 10'b0011110100,
    StCtrlRootKey        = 10'b0110101111,
    StCtrlInit           = 10'b0100000100,
    StCtrlCreatorRootKey = 10'b1000011101,
    StCtrlOwnerIntKey    = 10'b0001001010,
    StCtrlOwnerKey       = 10'b1101111110,
    StCtrlDisabled       = 10'b1010101000,
    StCtrlWipe           = 10'b0000110011,
    StCtrlInvalid        = 10'b1011000111
  } state_e;
  state_e state_q, state_d;

  // A variable that represents differentiates states before root key and after root key.
  logic initialized;

  // There are two versions of the key state, one for sealing one for attestation
  // Among each version, there are multiple shares
  // Each share is a fixed multiple of the entropy width
  logic [CDIs-1:0][Shares-1:0][EntropyRounds-1:0][EntropyWidth-1:0] key_state_d;
  logic [CDIs-1:0][Shares-1:0][EccWords-1:0][EccDataWidth-1:0] key_state_ecc_words_d;
  logic [CDIs-1:0][Shares-1:0][EccWords-1:0][EccDataWidth-1:0] key_state_q;
  logic [CDIs-1:0][Shares-1:0][EccWords-1:0][EccWidth-1:0] key_state_ecc_q;
  logic [CntWidth-1:0] cnt;
  logic [CdiWidth-1:0] cdi_cnt;

  // error conditions
  logic invalid_kmac_out;
  logic invalid_op;
  logic cnt_err;
  // states fall out of sparsely encoded range
  logic state_intg_err_q, state_intg_err_d;

  ///////////////////////////
  //  General operation decode
  ///////////////////////////

  logic adv_op, dis_op, gen_id_op, gen_sw_op, gen_hw_op, gen_op;
  assign adv_op    = (op_i == OpAdvance);
  assign gen_id_op = (op_i == OpGenId);
  assign gen_sw_op = (op_i == OpGenSwOut);
  assign gen_hw_op = (op_i == OpGenHwOut);
  assign dis_op    = ~(op_i inside {OpAdvance, OpGenId, OpGenSwOut, OpGenHwOut});
  assign gen_op    = (gen_id_op | gen_sw_op | gen_hw_op);

  ///////////////////////////
  //  interaction between software and main fsm
  ///////////////////////////
  // disable is treated like an advanced call
  logic advance_sel;
  logic disable_sel;
  logic gen_out_hw_sel;

  assign advance_sel    = op_start_i & adv_op    & en_i;
  assign gen_out_hw_sel = op_start_i & gen_hw_op & en_i;

  // disable is selected whenever a normal operation is not set
  assign disable_sel    = (op_start_i & dis_op) | !en_i;


  ///////////////////////////
  //  interaction between main control fsm and operation fsm
  ///////////////////////////

  // req/ack interface with op handling fsm
  logic op_req;
  logic op_ack;
  logic op_update;
  logic op_busy;
  logic disabled;
  logic invalid;

  logic adv_req, dis_req, id_req, gen_req;
  assign adv_req = op_req & adv_op;
  assign dis_req = op_req & dis_op;
  assign id_req  = op_req & gen_id_op;
  assign gen_req = op_req & (gen_sw_op | gen_hw_op);

  ///////////////////////////
  //  interaction between operation fsm and software
  ///////////////////////////
  // categories of keymgr errors
  logic [SyncErrLastIdx-1:0] sync_err;
  logic [SyncFaultLastIdx-1:0] sync_fault;
  logic [AsyncFaultLastIdx-1:0] async_fault;

  logic op_err;
  logic op_fault_err;

  // unlock sw binding configuration whenever an advance call is made without errors
  assign sw_binding_unlock_o = adv_req & op_ack & ~(op_err | op_fault_err);

  // error definition
  // check incoming kmac data validity
  // Only check during the periods when there is actual kmac output
  assign invalid_kmac_out = (op_update | op_ack) &
                            (~valid_data_chk(kmac_data_i[0]) |
                            (~valid_data_chk(kmac_data_i[1]) & KmacEnMasking));

  // async errors have nothing to do with the operation and thus should not
  // impact operation results.
  assign op_err = |sync_err;

  assign op_fault_err = |{sync_fault, async_fault};

  ///////////////////////////
  //  key update controls
  ///////////////////////////

  // update select can come from both main and operation fsm's
  keymgr_key_update_e update_sel, op_update_sel;

  // req from main control fsm to key update controls
  logic wipe_req;
  logic random_req;
  logic random_ack;

  // wipe and initialize take precedence
  assign update_sel = wipe_req             ? KeyUpdateWipe   :
                      random_req           ? KeyUpdateRandom :
                      init_o               ? KeyUpdateRoot   : op_update_sel;

  ///////////////////////////
  //  interaction between main fsm and prng
  ///////////////////////////

  assign prng_en_o = random_req | disabled | invalid | wipe_req;

  //////////////////////////
  // Main Control FSM
  //////////////////////////
  // SEC_CM: CTRL.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, StCtrlReset)

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      state_intg_err_q <= '0;
    end else begin
      state_intg_err_q <= state_intg_err_d;
    end
  end

  // prevents unknowns from reaching the outside world.
  // - whatever operation causes the input data select to be disabled should not expose the key
  //   state.
  // - when there are no operations, the key state also should be exposed.
  assign key_o.valid = op_req;

  assign cdi_sel_o = advance_sel ? cdi_cnt : op_cdi_sel_i;

  assign invalid_stage_sel_o = ~(stage_sel_o inside {Creator, OwnerInt, Owner});
  for (genvar i = 0; i < Shares; i++) begin : gen_key_out_assign
    assign key_o.key[i] = invalid_stage_sel_o ?
                          {EntropyRounds{entropy_i[i]}} :
                          key_state_q[cdi_sel_o][i];
  end


  //SEC_CM: CTRL.KEY.INTEGRITY
  assign key_state_ecc_words_d = key_state_d;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      key_state_q <= '0;
      key_state_ecc_q <= {TotalEccWords{prim_secded_pkg::SecdedInv7264ZeroEcc}};
    end else begin
      for (int i = 0; i < CDIs; i++) begin
        for (int j = 0; j < Shares; j++) begin
          for (int k = 0; k < EccWords; k++) begin
            {key_state_ecc_q[i][j][k], key_state_q[i][j][k]} <=
                prim_secded_pkg::prim_secded_inv_72_64_enc(key_state_ecc_words_d[i][j][k]);
          end
        end
      end
    end
  end

  logic [CDIs-1:0][Shares-1:0][EccWords-1:0] ecc_errs;
  for (genvar i = 0; i < CDIs; i++) begin : gen_ecc_loop_cdi
    for (genvar j = 0; j < Shares; j++) begin : gen_ecc_loop_shares
      for (genvar k = 0; k < EccWords; k++) begin : gen_ecc_loop_words
        logic [1:0] errs;
        prim_secded_inv_72_64_dec u_dec (
          .data_i({key_state_ecc_q[i][j][k], key_state_q[i][j][k]}),
          .data_o(),
          .syndrome_o(),
          .err_o(errs)
        );
        assign ecc_errs[i][j][k] = |errs;
      end
    end
  end

  // root key valid sync
  logic root_key_valid_q;

  prim_flop_2sync # (
    .Width(1)
  ) u_key_valid_sync (
    .clk_i,
    .rst_ni,
    .d_i(root_key_i.valid),
    .q_o(root_key_valid_q)
  );

  // Do not let the count toggle unless an advance operation is
  // selected
  assign cdi_cnt = op_req ? cnt[CdiWidth-1:0] : '0;

  always_comb begin
    key_state_d = key_state_q;
    data_valid_o = 1'b0;
    wipe_key_o = 1'b0;

    // if a wipe request arrives, immediately destroy the
    // keys regardless of current state
    unique case (update_sel)
      KeyUpdateRandom: begin
        for (int i = 0; i < CDIs; i++) begin
          for (int j = 0; j < Shares; j++) begin
            // Load each share with the same randomness so we can
            // later simply XOR root key on them
            key_state_d[i][j][cnt[EntropyRndWidth-1:0]] = entropy_i[i];
          end
        end
      end

      KeyUpdateRoot: begin
        if (root_key_valid_q) begin
          for (int i = 0; i < CDIs; i++) begin
            if (KmacEnMasking) begin : gen_two_share_key
              key_state_d[i][0] ^= root_key_i.key_share0;
              key_state_d[i][1] ^= root_key_i.key_share1;
            end else begin : gen_one_share_key
              key_state_d[i][0] = root_key_i.key_share0 ^ root_key_i.key_share1;
              key_state_d[i][1] = '0;
            end
          end
        end else begin
          // if root key is not valid, load and invalid value
          for (int i = 0; i < CDIs; i++) begin
              key_state_d[i][0] = '0;
              key_state_d[i][1] = '{default: '1};
          end
        end
      end

      KeyUpdateKmac: begin
        data_valid_o = gen_op;
        key_state_d[cdi_sel_o] = (adv_op || dis_op) ? kmac_data_i : key_state_q[cdi_sel_o];
      end

      KeyUpdateWipe: begin
        wipe_key_o = 1'b1;
        for (int i = 0; i < CDIs; i++) begin
          for (int j = 0; j < Shares; j++) begin
            key_state_d[i][j] = {EntropyRounds{entropy_i[j]}};
          end
        end
      end

      default:;
    endcase // unique case (update_sel)
  end

  // SEC_CM: CTRL.CTR.REDUN
  prim_count #(
    .Width(CntWidth)
  ) u_cnt (
    .clk_i,
    .rst_ni,
    .clr_i(op_ack | random_ack),
    .set_i('0),
    .set_cnt_i('0),
    .incr_en_i(op_update | random_req),
    .decr_en_i(1'b0),
    .step_i(CntWidth'(1'b1)),
    .cnt_o(cnt),
    .cnt_next_o(),
    .err_o(cnt_err)
  );


  prim_mubi4_sender u_hw_sel (
    .clk_i,
    .rst_ni,
    .mubi_i (prim_mubi_pkg::mubi4_bool_to_mubi(gen_out_hw_sel)),
    .mubi_o (hw_sel_o)
  );

  // when in a state that accepts commands, look at op_ack for completion
  // when in a state that does not accept commands, wait for other triggers.
  assign op_done_o = op_req ? op_ack :
                     (init_o | invalid_op);


  // There are 3 possibilities
  // advance to next state (software command)
  // advance to disabled state (software command)
  // advance to invalid state (detected fault)
  logic adv_state;
  logic dis_state;
  logic inv_state;
  assign adv_state = op_ack & adv_req & ~op_err;
  assign dis_state = op_ack & dis_req;

  // SEC_CM: CTRL.FSM.LOCAL_ESC
  // begin invalidation when faults are observed.
  // sync faults only invalidate on transaction boudaries
  // async faults begin invalidating immediately
  assign inv_state = |fault_o;

  always_comb begin
    // persistent data
    state_d = state_q;

    // request to op handling
    op_req = 1'b0;
    random_req = 1'b0;
    random_ack = 1'b0;

    // request to key updates
    wipe_req = 1'b0;

    // invalid operation issued
    invalid_op = '0;

    // data update and select signals
    stage_sel_o = Disable;

    // indication that state is disabled
    disabled = 1'b0;

    // indication that state is invalid
    invalid = 1'b0;

    // enable prng toggling
    prng_reseed_req_o = 1'b0;

    // initialization complete
    init_o = 1'b0;

    // Most states are initialized, mark the exceptions
    initialized = 1'b1;

    // if state is ever faulted, hold on to this indication
    // until reset.
    state_intg_err_d = state_intg_err_q;

    unique case (state_q)
      // Only advance can be called from reset state
      StCtrlReset: begin
        initialized = 1'b0;

        // always use random data for advance, since out of reset state
        // the key state will be randomized.
        stage_sel_o = Disable;

        // key state is updated when it is an advance call
        // all other operations are invalid, including disable
        invalid_op = op_start_i & ~advance_sel;

        // if there was a structural fault before anything began, wipe immediately
        if (inv_state) begin
          state_d = StCtrlWipe;
        end else if (advance_sel) begin
          state_d = StCtrlEntropyReseed;
        end
      end

      // reseed entropy
      StCtrlEntropyReseed: begin
        initialized = 1'b0;
        prng_reseed_req_o = 1'b1;

        if (prng_reseed_ack_i) begin
          state_d = StCtrlRandom;
        end
      end

      // This state does not accept any command.
      StCtrlRandom: begin
        initialized = 1'b0;
        random_req = 1'b1;

        // when mask population is complete, xor the root_key into the zero share
        // if in the future the root key is updated to 2 shares, it will direclty overwrite
        // the values here
        if (int'(cnt) == EntropyRounds-1) begin
          random_ack = 1'b1;
          state_d = StCtrlRootKey;
        end
      end

      // load the root key.
      StCtrlRootKey: begin
        init_o = 1'b1;
        initialized = 1'b1;
        state_d = en_i ? StCtrlInit : StCtrlWipe;
      end

      // Beginning from the Init state, operations are accepted.
      // Only valid operation is advance state. If invalid command received,
      // random data is selected for operation and no persistent state is changed.
      StCtrlInit: begin
        op_req = op_start_i;

        // when advancing select creator data, otherwise use random input
        stage_sel_o = advance_sel ? Creator : Disable;
        invalid_op = op_start_i & ~(advance_sel | disable_sel);

        if (!en_i || inv_state) begin
          state_d = StCtrlWipe;
        end else if (dis_state) begin
          state_d = StCtrlDisabled;
        end else if (adv_state) begin
          state_d = StCtrlCreatorRootKey;
        end
      end

      // all commands  are valid during this stage
      StCtrlCreatorRootKey: begin
        op_req = op_start_i;

        // when generating, select creator data input
        // when advancing, select owner intermediate key as target
        // when disabling, select random data input
        stage_sel_o = disable_sel ? Disable  :
                      advance_sel ? OwnerInt : Creator;

        if (!en_i || inv_state) begin
          state_d = StCtrlWipe;
        end else if (dis_state) begin
          state_d = StCtrlDisabled;
        end else if (adv_state) begin
          state_d = StCtrlOwnerIntKey;
        end
      end

      // all commands are valid during this stage
      StCtrlOwnerIntKey: begin
        op_req = op_start_i;

        // when generating, select owner intermediate data input
        // when advancing, select owner as target
        // when disabling, select random data input
        stage_sel_o = disable_sel ? Disable  :
                      advance_sel ? Owner : OwnerInt;

        if (!en_i || inv_state) begin
          state_d = StCtrlWipe;
        end else if (dis_state) begin
          state_d = StCtrlDisabled;
        end else if (adv_state) begin
          state_d = StCtrlOwnerKey;
        end
      end

      // all commands are valid during this stage
      // however advance goes directly to disabled state
      StCtrlOwnerKey: begin
        op_req = op_start_i;

        // when generating, select owner data input
        // when advancing, select disable as target
        // when disabling, select random data input
        stage_sel_o = disable_sel | advance_sel ? Disable : Owner;

        if (!en_i || inv_state) begin
          state_d = StCtrlWipe;
        end else if (adv_state || dis_state) begin
          state_d = StCtrlDisabled;
        end
      end

      // The wipe state immediately clears out the key state, but waits for any ongoing
      // transaction to finish before going to disabled state.
      // Unlike the random state, this is an immedaite shutdown request, so all parts of the
      // key are wiped.
      StCtrlWipe: begin
        wipe_req = 1'b1;
        // if there was already an operation ongoing, maintain the request until completion
        op_req = op_busy;
        invalid_op = op_start_i;

        // If the enable is dropped during the middle of a transaction, we clear and wait for that
        // transaction to gracefully complete (if it can).
        // There are two scenarios:
        // 1. the operation completed right when we started wiping, in which case the done would
        //    clear the start.
        // 2. the operation completed before we started wiping, or there was never an operation to
        //    begin with (op_start_i == 0), in this case, don't wait and immediately transition
        if (!op_start_i) begin
          state_d = StCtrlInvalid;
        end
      end

      // StCtrlDisabled and StCtrlInvalid are almost functionally equivalent
      // The only difference is that Disabled is entered through software invocation,
      // while Invalid is entered through life cycle disable or operational fault.
      //
      // Both states continue to kick off random transactions
      // All transactions are treated as invalid despite completing
      StCtrlDisabled: begin
        op_req = op_start_i;
        disabled = 1'b1;

        if (!en_i || inv_state) begin
          state_d = StCtrlWipe;
        end
      end

      StCtrlInvalid: begin
        op_req = op_start_i;
        invalid = 1'b1;
      end

      // latch the fault indication and start to wipe the key manager
      default: begin
        state_intg_err_d = 1'b1;
        state_d = StCtrlWipe;
      end

    endcase // unique case (state_q)
  end // always_comb

  // Current working state provided for software read
  // Certain states are collapsed for simplicity
  keymgr_working_state_e last_working_st;
  logic update_en;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      last_working_st <= StReset;
    end else if (update_en) begin
      last_working_st <= working_state_o;
    end
  end

  always_comb begin
    update_en = 1'b1;
    working_state_o = StInvalid;

    unique case (state_q)
      StCtrlReset, StCtrlEntropyReseed, StCtrlRandom:
        working_state_o = StReset;

      StCtrlRootKey, StCtrlInit:
        working_state_o = StInit;

      StCtrlCreatorRootKey:
        working_state_o = StCreatorRootKey;

      StCtrlOwnerIntKey:
        working_state_o = StOwnerIntKey;

      StCtrlOwnerKey:
        working_state_o = StOwnerKey;

      StCtrlDisabled:
        working_state_o = StDisabled;

      StCtrlWipe: begin
        update_en = 1'b0;
        working_state_o = last_working_st;
      end

      StCtrlInvalid:
        working_state_o = StInvalid;

      default:
        working_state_o = StInvalid;
    endcase // unique case (state_q)
  end

  always_comb begin
    status_o = OpIdle;
    if (op_done_o) begin
      // It is possible for an operation to finish the same cycle en_i goes low.
      // The main fsm handling is one cycle behind, but still report operation
      // fail.
      status_o = |{error_o, fault_o} ? OpDoneFail : OpDoneSuccess;
    end else if (op_start_i) begin
      status_o = OpWip;
    end
  end


  /////////////////////////
  // Operateion state, handle advance and generate
  /////////////////////////

  logic op_fsm_err;
  keymgr_op_state_ctrl u_op_state (
    .clk_i,
    .rst_ni,
    .adv_req_i(adv_req),
    .dis_req_i(dis_req),
    .id_req_i(id_req),
    .gen_req_i(gen_req),
    .cnt_i(cdi_cnt),
    .op_ack_o(op_ack),
    .op_busy_o(op_busy),
    .op_update_o(op_update),
    .kmac_done_i,
    .adv_en_o,
    .id_en_o,
    .gen_en_o,
    .op_fsm_err_o(op_fsm_err)
  );

  // operational state cross check.  The state value must be consistent with
  // the input operations.
  logic op_state_cmd_err;
  assign op_state_cmd_err = (adv_en_o & ~(advance_sel | disable_sel)) |
                            (gen_en_o & ~gen_op);

  // operations fsm update precedence
  // when in invalid state, always update.
  // when in disabled state, always update unless a fault is encountered.
  assign op_update_sel = (op_ack | op_update) & invalid      ? KeyUpdateKmac :
                         (op_ack | op_update) & op_fault_err ? KeyUpdateWipe :
                         (op_ack | op_update) & disabled     ? KeyUpdateKmac :
                         (op_ack | op_update) & op_err       ? KeyUpdateIdle :
                         (op_ack | op_update)                ? KeyUpdateKmac : KeyUpdateIdle;


  ///////////////////////////////
  // Suppress kmac return data
  ///////////////////////////////

  logic data_fsm_err;
  keymgr_data_en_state u_data_en (
    .clk_i,
    .rst_ni,
    .hw_sel_i(hw_sel_o),
    .adv_en_i(adv_en_o),
    .id_en_i(id_en_o),
    .gen_en_i(gen_en_o),
    .op_done_i(op_done_o),
    .op_start_i,
    .data_hw_en_o,
    .data_sw_en_o,
    .fsm_err_o(data_fsm_err)
  );

  /////////////////////////
  // Cross-checks, errors and faults
  /////////////////////////

  logic vld_state_change_d, vld_state_change_q;
  assign vld_state_change_d = (state_d != state_q) &
                              (state_d inside {StCtrlRootKey,
                                               StCtrlCreatorRootKey,
                                               StCtrlOwnerIntKey,
                                               StCtrlOwnerKey});

  // capture for cross check in following cycle
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      vld_state_change_q <= '0;
    end else begin
      vld_state_change_q <= vld_state_change_d;
    end
  end

  // state cross check
  // if the state advanced, ensure that it was due to an advanced operation
  logic state_change_err;
  assign state_change_err = vld_state_change_q & !adv_op;

  keymgr_err u_err (
    .clk_i,
    .rst_ni,
    .invalid_op_i(invalid_op),
    .disabled_i(disabled | (initialized & ~en_i)),
    .invalid_i(invalid),
    .kmac_input_invalid_i,
    .shadowed_update_err_i,
    .kmac_op_err_i,
    .invalid_kmac_out_i(invalid_kmac_out),
    .sideload_sel_err_i,
    .kmac_cmd_err_i,
    .kmac_fsm_err_i,
    .kmac_done_err_i,
    .regfile_intg_err_i,
    .shadowed_storage_err_i,
    .ctrl_fsm_err_i(state_intg_err_q | state_intg_err_d),
    .data_fsm_err_i(data_fsm_err),
    .op_fsm_err_i(op_fsm_err),
    .ecc_err_i(|ecc_errs),
    .state_change_err_i(state_change_err),
    .op_state_cmd_err_i(op_state_cmd_err),
    .cnt_err_i(cnt_err),
    .reseed_cnt_err_i,
    .sideload_fsm_err_i,

    .op_update_i(op_update),
    .op_done_i(op_done_o),

    .sync_err_o(sync_err),
    .async_err_o(),
    .sync_fault_o(sync_fault),
    .async_fault_o(async_fault),
    .error_o,
    .fault_o
  );

  ///////////////////////////////
  // Functions
  ///////////////////////////////

  // unclear what this is supposed to be yet
  // right now just check to see if it not all 0's and not all 1's
 function automatic logic valid_data_chk (logic [KeyWidth-1:0] value);

    return |value & ~&value;

  endfunction // byte_mask

  /////////////////////////////////
  // Assertions
  /////////////////////////////////

  // This assertion will not work if fault_status ever takes on metafields such as
  // qe / re etc.
  `ASSERT_INIT(SameErrCnt_A, $bits(keymgr_reg2hw_fault_status_reg_t) ==
                             (SyncFaultLastIdx + AsyncFaultLastIdx))

  // stage select should always be Disable whenever it is not enabled
  `ASSERT(StageDisableSel_A, !en_i |-> stage_sel_o == Disable)

  // Unless it is a legal command, only select disable
  `ASSERT(InitLegalCommands_A, op_start_i & en_i & state_q inside {StCtrlInit} &
                               !(op_i inside {OpAdvance}) |-> stage_sel_o == Disable)

  // All commands are legal, so select disable only if operation is disable
  `ASSERT(GeneralLegalCommands_A, op_start_i & en_i &
                                  state_q inside {StCtrlCreatorRootKey, StCtrlOwnerIntKey} &
                                  (op_i inside {OpDisable}) |-> stage_sel_o == Disable)

  `ASSERT(OwnerLegalCommands_A, op_start_i & en_i & state_q inside {StCtrlOwnerKey} &
                                (op_i inside {OpAdvance, OpDisable}) |-> stage_sel_o == Disable)

  // load_key should not be high if there is no ongoing operation
  `ASSERT(LoadKey_A, key_o.valid |-> op_start_i)

  // The count value should always be 0 when a transaction start
  `ASSERT(CntZero_A, $rose(op_start_i) |-> cnt == '0)

  // Whenever a transaction completes, data_en must return to 0 on the next cycle
  `ASSERT(DataEnDis_A, op_start_i & op_done_o |=> ~data_hw_en_o && ~data_sw_en_o)

  // Whenever data enable asserts, it must be the case that there was a generate or
  // id operation
  `ASSERT(DataEn_A, data_hw_en_o | data_sw_en_o |-> (id_en_o | gen_en_o) & ~adv_en_o)

  // Check that the FSM is linear and does not contain any loops
  `ASSERT_FPV_LINEAR_FSM(SecCmCFILinear_A, state_q, state_e)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager CFGEN
// TBD This should be enhanced in the future to contain a shadow copy

`include "prim_assert.sv"

module keymgr_cfg_en #(
  // controls whether clear has an effect on output value during non-init
  parameter bit NonInitClr = 1'b1
) (
  input clk_i,
  input rst_ni,
  input init_i,
  input en_i,
  input set_i,
  input clr_i,
  output logic out_o
);

  logic out_q;
  logic init_q;

  logic vld_clr;
  logic vld_set;
  logic vld_dis;

  assign vld_clr = init_q && clr_i;
  assign vld_set = init_q && set_i;
  assign vld_dis = init_q && !en_i;

  // the same cycle where clear is asserted should already block future
  // configuration
  logic out_clr;
  assign out_clr = NonInitClr ? clr_i : vld_clr;
  assign out_o = ~out_clr & out_q & en_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      init_q <= '0;
    end else if (init_q && !en_i) begin
      init_q <= '0;
    end else if (init_i && en_i) begin
      init_q <= 1'b1;
    end
  end

  // clearing the configure enable always has higher priority than setting
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      out_q <= 1'b1;
    end else if (vld_dis) begin
      out_q <= 1'b0;
    end else if (vld_set) begin
      out_q <= 1'b1;
    end else if (out_clr) begin
      out_q <= 1'b0;
    end
  end

endmodule // keymgr_cfg_en


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager date enable generation
// This is a redundant alternative to data_valid

`include "prim_assert.sv"

module keymgr_data_en_state
  import keymgr_pkg::*;
  import keymgr_reg_pkg::*;
(
  input clk_i,
  input rst_ni,
  input prim_mubi_pkg::mubi4_t hw_sel_i,
  input adv_en_i,
  input id_en_i,
  input gen_en_i,
  input op_done_i,
  input op_start_i,
  output logic data_hw_en_o,
  output logic data_sw_en_o,
  output logic fsm_err_o
);

  import prim_mubi_pkg::mubi4_test_true_strict;
  import prim_mubi_pkg::mubi4_test_true_loose;
  import prim_mubi_pkg::mubi4_test_false_strict;
  import prim_mubi_pkg::mubi4_test_false_loose;

  // This is a separate data path from the FSM used to control the data_en outputs
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 6 -n 10 \
  //      -s 2015444891 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||| (33.33%)
  //  6: |||||||||||||||||||| (40.00%)
  //  7: ||||||||||||| (26.67%)
  //  8: --
  //  9: --
  // 10: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 7
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 7
  //
  localparam int DataStateWidth = 10;
  typedef enum logic [DataStateWidth-1:0] {
    StCtrlDataIdle    = 10'b1000010000,
    StCtrlDataHwEn    = 10'b0001100100,
    StCtrlDataSwEn    = 10'b1110101110,
    StCtrlDataDis     = 10'b0010011111,
    StCtrlDataWait    = 10'b0111110011,
    StCtrlDataInvalid = 10'b1111001001
  } state_e;

  state_e state_d, state_q;

  // SEC_CM: DATA.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, StCtrlDataIdle)

  // The below control path is used for modulating the datapath to sideload and sw keys.
  // This path is separate from the data_valid_o path, thus creating two separate attack points.
  // The data is only enabled when a non-advance operation is invoked.
  // When an advance operation is called, the data is disabled. It will stay disabled until an
  // entire completion sequence is seen (op_done_o assert -> start_i de-assertion).
  // When a generate operation is called, the data is enabled.  However, any indication of this
  // supposedly being an advance call will force the path to disable again.
  always_comb begin
    state_d = state_q;
    fsm_err_o = 1'b0;
    data_hw_en_o = 1'b0;
    data_sw_en_o = 1'b0;
    unique case (state_q)

      StCtrlDataIdle: begin
        if (adv_en_i) begin
          state_d = StCtrlDataDis;
        end else if ((id_en_i || gen_en_i) && mubi4_test_true_strict(hw_sel_i)) begin
          state_d = StCtrlDataHwEn;
        end else if ((id_en_i || gen_en_i) && mubi4_test_false_strict(hw_sel_i)) begin
          state_d = StCtrlDataSwEn;
        end else if (id_en_i || gen_en_i) begin
          state_d = StCtrlDataDis;
        end
      end

      StCtrlDataHwEn: begin
        data_hw_en_o = 1'b1;
        if (op_done_i) begin
          state_d = StCtrlDataWait;
        end else if (adv_en_i || mubi4_test_false_loose(hw_sel_i)) begin
          state_d = StCtrlDataDis;
        end
      end

      StCtrlDataSwEn: begin
        data_sw_en_o = 1'b1;
        if (op_done_i) begin
          state_d = StCtrlDataWait;
        end else if (adv_en_i || mubi4_test_true_loose(hw_sel_i)) begin
          state_d = StCtrlDataDis;
        end
      end

      StCtrlDataDis: begin
        if (op_done_i) begin
          state_d = StCtrlDataWait;
        end
      end

      StCtrlDataWait: begin
        if (!op_start_i) begin
          state_d = StCtrlDataIdle;
        end
      end

      default: begin
        fsm_err_o = 1'b1;
      end


    endcase // unique case (state_q)
  end


endmodule // keymgr_data_en_state


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager error and fault collection
//

`include "prim_assert.sv"

module keymgr_err
  import keymgr_pkg::*;
  import keymgr_reg_pkg::*;
(
  input clk_i,
  input rst_ni,

  input invalid_op_i,
  input disabled_i,
  input invalid_i,
  input kmac_input_invalid_i,
  input shadowed_update_err_i,
  input kmac_op_err_i,
  input invalid_kmac_out_i,
  input sideload_sel_err_i,
  input kmac_cmd_err_i,
  input kmac_fsm_err_i,
  input kmac_done_err_i,
  input regfile_intg_err_i,
  input shadowed_storage_err_i,
  input ctrl_fsm_err_i,
  input data_fsm_err_i,
  input op_fsm_err_i,
  input ecc_err_i,
  input state_change_err_i,
  input op_state_cmd_err_i,
  input cnt_err_i,
  input reseed_cnt_err_i,
  input sideload_fsm_err_i,

  input op_update_i,
  input op_done_i,

  // The following outputs are very similar, but have slightly different timing for
  // for CDIs on sync errors/faults.
  // Advance operations must go through for all CDIs.
  // The sync_err/fault outputs register when any CDI completes and helps with
  // the appropriate behavior on key state change.
  // The sync error_o/fault_o outputs on the other hand only output when the entire
  // operation is complete, which could be multiple CDIs.
  output logic [SyncErrLastIdx-1:0] sync_err_o,
  output logic [AsyncErrLastIdx-1:0] async_err_o,
  output logic [SyncFaultLastIdx-1:0] sync_fault_o,
  output logic [AsyncFaultLastIdx-1:0] async_fault_o,
  output logic [ErrLastPos-1:0] error_o,
  output logic [FaultLastPos-1:0] fault_o
);

  // Advance calls are made up of multiple rounds of kmac operations.
  // Any sync error that occurs is treated as an error of the entire call.
  // Therefore sync errors that happen before the end of the call must be
  // latched.
  logic[SyncErrLastIdx-1:0] sync_err_q, sync_err_d;
  logic[SyncFaultLastIdx-1:0] sync_fault_q, sync_fault_d;

  logic err_vld;
  assign err_vld = op_update_i | op_done_i;

  // sync errors
  // When an operation encounters a fault, the operation is always rejected as the FSM
  // transitions to wipe.  When an operation is ongoing and en drops, it is also rejected.
  assign sync_err_d[SyncErrInvalidOp] = err_vld & (invalid_op_i |
                                                   disabled_i |
                                                   invalid_i |
                                                   (|fault_o));
  assign sync_err_d[SyncErrInvalidIn] = err_vld & kmac_input_invalid_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      sync_err_q <= '0;
    end else if (op_done_i) begin
      sync_err_q <= '0;
    end else if (op_update_i) begin
      sync_err_q <= sync_err_d;
    end
  end
  assign sync_err_o = sync_err_q | sync_err_d;

  // async errors
  assign async_err_o[AsyncErrShadowUpdate] = shadowed_update_err_i;

  // sync faults
  assign sync_fault_d[SyncFaultKmacOp] = err_vld & kmac_op_err_i;
  assign sync_fault_d[SyncFaultKmacOut] = err_vld & invalid_kmac_out_i;
  assign sync_fault_d[SyncFaultSideSel] = err_vld & sideload_sel_err_i;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      sync_fault_q <= '0;
    end else if (op_done_i) begin
      sync_fault_q <= '0;
    end else if (op_update_i) begin
      sync_fault_q <= sync_fault_d;
    end
  end
  assign sync_fault_o = sync_fault_q | sync_fault_d;

  // async faults
  logic [AsyncFaultLastIdx-1:0] async_fault_q, async_fault_d;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      async_fault_q <= '0;
    end else begin
      async_fault_q <= async_fault_o;
    end
  end
  assign async_fault_o = async_fault_q | async_fault_d;
  assign async_fault_d[AsyncFaultKmacCmd]  = kmac_cmd_err_i;
  assign async_fault_d[AsyncFaultKmacFsm]  = kmac_fsm_err_i;
  assign async_fault_d[AsyncFaultKmacDone] = kmac_done_err_i;
  assign async_fault_d[AsyncFaultRegIntg]  = regfile_intg_err_i;
  assign async_fault_d[AsyncFaultShadow ]  = shadowed_storage_err_i;
  assign async_fault_d[AsyncFaultFsmIntg]  = ctrl_fsm_err_i | data_fsm_err_i | op_fsm_err_i;
  assign async_fault_d[AsyncFaultKeyEcc]   = ecc_err_i;

  // SEC_CM: CTRL.FSM.CONSISTENCY
  assign async_fault_d[AsyncFaultFsmChk]   = state_change_err_i | op_state_cmd_err_i;
  assign async_fault_d[AsyncFaultCntErr ]  = cnt_err_i;
  assign async_fault_d[AsyncFaultRCntErr]  = reseed_cnt_err_i;
  assign async_fault_d[AsyncFaultSideErr]  = sideload_fsm_err_i;

  // certain errors/faults can only happen when there's an actual kmac transaction,
  // others can happen with or without.
  assign error_o[ErrInvalidOp]    = op_done_i & sync_err_o[SyncErrInvalidOp];
  assign error_o[ErrInvalidIn]    = op_done_i & sync_err_o[SyncErrInvalidIn];
  assign error_o[ErrShadowUpdate] = async_err_o[AsyncErrShadowUpdate];

  // output to fault code register
  assign fault_o[FaultKmacOp]     = op_done_i & sync_fault_o[SyncFaultKmacOp];
  assign fault_o[FaultKmacOut]    = op_done_i & sync_fault_o[SyncFaultKmacOut];
  assign fault_o[FaultSideSel]    = op_done_i & sync_fault_o[SyncFaultSideSel];
  assign fault_o[FaultKmacCmd]    = async_fault_o[AsyncFaultKmacCmd];
  assign fault_o[FaultKmacFsm]    = async_fault_o[AsyncFaultKmacFsm];
  assign fault_o[FaultKmacDone]   = async_fault_o[AsyncFaultKmacDone];
  assign fault_o[FaultRegIntg]    = async_fault_o[AsyncFaultRegIntg];
  assign fault_o[FaultShadow]     = async_fault_o[AsyncFaultShadow];
  assign fault_o[FaultCtrlFsm]    = async_fault_o[AsyncFaultFsmIntg];
  assign fault_o[FaultCtrlFsmChk] = async_fault_o[AsyncFaultFsmChk];
  assign fault_o[FaultCtrlCnt]    = async_fault_o[AsyncFaultCntErr];
  assign fault_o[FaultReseedCnt]  = async_fault_o[AsyncFaultRCntErr];
  assign fault_o[FaultSideFsm]    = async_fault_o[AsyncFaultSideErr];
  assign fault_o[FaultKeyEcc]     = async_fault_o[AsyncFaultKeyEcc];


endmodule // keymgr_err


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager input checks
// Checks input data for errors

`include "prim_assert.sv"

// We should also check for input validity
module keymgr_input_checks import keymgr_pkg::*; #(
  parameter bit KmacEnMasking = 1'b1
) (
  input rom_ctrl_pkg::keymgr_data_t rom_digest_i,
  input [2**StageWidth-1:0][31:0] max_key_versions_i,
  input keymgr_stage_e stage_sel_i,
  input hw_key_req_t key_i,
  input [31:0] key_version_i,
  input [KeyWidth-1:0] creator_seed_i,
  input [KeyWidth-1:0] owner_seed_i,
  input [DevIdWidth-1:0] devid_i,
  input [HealthStateWidth-1:0] health_state_i,
  output logic creator_seed_vld_o,
  output logic owner_seed_vld_o,
  output logic devid_vld_o,
  output logic health_state_vld_o,
  output logic key_version_vld_o,
  output logic key_vld_o,
  output logic rom_digest_vld_o
);

  logic [31:0] cur_max_key_version;
  assign cur_max_key_version = max_key_versions_i[stage_sel_i];

  // key version must be smaller than or equal to max version
  assign key_version_vld_o = key_version_i <= cur_max_key_version;

  // general data check
  logic [MaxWidth-1:0] creator_seed_padded, owner_seed_padded, devid_padded, health_state_padded;

  prim_msb_extend #(
    .InWidth(KeyWidth),
    .OutWidth(MaxWidth)
  ) u_creator_seed (
    .in_i(creator_seed_i),
    .out_o(creator_seed_padded)
  );

  prim_msb_extend #(
    .InWidth(KeyWidth),
    .OutWidth(MaxWidth)
  ) u_owner_seed (
    .in_i(owner_seed_i),
    .out_o(owner_seed_padded)
  );

  prim_msb_extend #(
    .InWidth(DevIdWidth),
    .OutWidth(MaxWidth)
  ) u_devid (
    .in_i(devid_i),
    .out_o(devid_padded)
  );

  prim_msb_extend #(
    .InWidth(HealthStateWidth),
    .OutWidth(MaxWidth)
  ) u_health_state (
    .in_i(health_state_i),
    .out_o(health_state_padded)
  );

  assign creator_seed_vld_o = valid_chk(creator_seed_padded);
  assign owner_seed_vld_o = valid_chk(owner_seed_padded);
  assign devid_vld_o = valid_chk(devid_padded);
  assign health_state_vld_o = valid_chk(health_state_padded);

  // key check
  logic unused_key_vld;
  assign unused_key_vld = key_i.valid;

  localparam int KeyShares = KmacEnMasking ? Shares : 1;
  logic [KeyShares-1:0][MaxWidth-1:0] key_padded;
  logic [KeyShares-1:0] key_chk;

  for (genvar i = 0; i < KeyShares; i++) begin : gen_key_chk
    prim_msb_extend #(
      .InWidth(KeyWidth),
      .OutWidth(MaxWidth)
    ) u_key_pad (
      .in_i(key_i.key[i]),
      .out_o(key_padded[i])
    );

    assign key_chk[i] = valid_chk(key_padded[i]);
  end

  assign key_vld_o = &key_chk;

  // rom digest check
  assign rom_digest_vld_o = rom_digest_i.valid &
                            valid_chk(MaxWidth'(rom_digest_i.data));

  // checks for all 0's or all 1's of value
  function automatic logic valid_chk (logic [MaxWidth-1:0] value);

    return |value & ~&value;

  endfunction // valid_chk


endmodule // keymgr_input_checks


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager interface to kmac
//

`include "prim_assert.sv"

module keymgr_kmac_if import keymgr_pkg::*;(
  input clk_i,
  input rst_ni,

  // data input interfaces
  input [AdvDataWidth-1:0] adv_data_i,
  input [IdDataWidth-1:0] id_data_i,
  input [GenDataWidth-1:0] gen_data_i,
  input [3:0] inputs_invalid_i,
  output logic inputs_invalid_o,

  // keymgr control to select appropriate inputs
  input adv_en_i,
  input id_en_i,
  input gen_en_i,
  output logic done_o,
  output logic [Shares-1:0][kmac_pkg::AppDigestW-1:0] data_o,

  // actual connection to kmac
  output kmac_pkg::app_req_t kmac_data_o,
  input  kmac_pkg::app_rsp_t kmac_data_i,

  // entropy input
  output logic prng_en_o,
  input [Shares-1:0][RandWidth-1:0] entropy_i,

  // error outputs
  output logic fsm_error_o,
  output logic kmac_error_o,
  output logic kmac_done_error_o,
  output logic cmd_error_o
);


  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 6 -n 10 \
  //      -s 2292624416 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||||||| (46.67%)
  //  6: ||||||||||||||||| (40.00%)
  //  7: ||||| (13.33%)
  //  8: --
  //  9: --
  // 10: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 7
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 9
  //
  localparam int StateWidth = 10;
  typedef enum logic [StateWidth-1:0] {
    StIdle    = 10'b1110100010,
    StTx      = 10'b0010011011,
    StTxLast  = 10'b0101000000,
    StOpWait  = 10'b1000101001,
    StClean   = 10'b1111111101,
    StError   = 10'b0011101110
  } data_state_e;

  localparam int AdvRem = AdvDataWidth % KmacDataIfWidth;
  localparam int IdRem  = IdDataWidth  % KmacDataIfWidth;
  localparam int GenRem = GenDataWidth % KmacDataIfWidth;

  // the remainder must be in number of bytes
  `ASSERT_INIT(AdvRemBytes_A, AdvRem % 8 == 0)
  `ASSERT_INIT(IdRemBytes_A,  IdRem  % 8 == 0)
  `ASSERT_INIT(GenRemBytes_A, GenRem % 8 == 0)

  // Number of kmac transactions required
  localparam int AdvRounds = (AdvDataWidth + KmacDataIfWidth - 1) / KmacDataIfWidth;
  localparam int IdRounds  = (IdDataWidth + KmacDataIfWidth - 1) / KmacDataIfWidth;
  localparam int GenRounds = (GenDataWidth + KmacDataIfWidth - 1) / KmacDataIfWidth;
  localparam int MaxRounds = KDFMaxWidth  / KmacDataIfWidth;

  // calculated parameters for number of roudns and interface width
  localparam int CntWidth = $clog2(MaxRounds);
  localparam int IfBytes = KmacDataIfWidth / 8;
  localparam int DecoyCopies = KmacDataIfWidth / RandWidth;
  localparam int DecoyOutputCopies = (kmac_pkg::AppDigestW / RandWidth) * Shares;

  localparam int unsigned LastAdvRoundInt = AdvRounds - 1;
  localparam int unsigned LastIdRoundInt = IdRounds - 1;
  localparam int unsigned LastGenRoundInt = GenRounds - 1;
  localparam bit [CntWidth-1:0] LastAdvRound = LastAdvRoundInt[CntWidth-1:0];
  localparam bit [CntWidth-1:0] LastIdRound = LastIdRoundInt[CntWidth-1:0];
  localparam bit [CntWidth-1:0] LastGenRound = LastGenRoundInt[CntWidth-1:0];

  // byte mask for the last transfer
  localparam logic [IfBytes-1:0] AdvByteMask = (AdvRem > 0) ? (2**(AdvRem/8)-1) : {IfBytes{1'b1}};
  localparam logic [IfBytes-1:0] IdByteMask  = (IdRem > 0)  ? (2**(IdRem/8)-1)  : {IfBytes{1'b1}};
  localparam logic [IfBytes-1:0] GenByteMask = (GenRem > 0) ? (2**(GenRem/8)-1) : {IfBytes{1'b1}};

  logic [MaxRounds-1:0][KmacDataIfWidth-1:0] adv_data;
  logic [MaxRounds-1:0][KmacDataIfWidth-1:0] id_data;
  logic [MaxRounds-1:0][KmacDataIfWidth-1:0] gen_data;
  logic [CntWidth-1:0] cnt;
  logic [CntWidth-1:0] rounds;
  logic [KmacDataIfWidth-1:0] decoy_data;
  logic valid;
  logic last;
  logic [IfBytes-1:0] strb;
  logic cnt_clr, cnt_set, cnt_en;
  logic start;
  logic [3:0] inputs_invalid_d, inputs_invalid_q;
  logic clr_err;
  logic kmac_done_vld;
  logic cmd_chk;

  data_state_e state_q, state_d;

  // 0 pad to the appropriate width
  // this is basically for scenarios where *DataWidth % KmacDataIfWidth != 0
  assign adv_data = KDFMaxWidth'(adv_data_i);
  assign id_data  = KDFMaxWidth'(id_data_i);
  assign gen_data = KDFMaxWidth'(gen_data_i);

  assign start = adv_en_i | id_en_i | gen_en_i;

  logic cnt_err;
  // SEC_CM: KMAC_IF.CTR.REDUN
  prim_count #(
    .Width(CntWidth),
    .ResetValue({CntWidth{1'b1}})
  ) u_cnt (
    .clk_i,
    .rst_ni,
    .clr_i(cnt_clr),
    .set_i(cnt_set),
    .set_cnt_i(rounds),
    .incr_en_i(1'b0),
    .decr_en_i(cnt_en),
    .step_i(CntWidth'(1'b1)),
    .cnt_o(cnt),
    .cnt_next_o(),
    .err_o(cnt_err)
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      inputs_invalid_q <= '0;
    end else begin
      inputs_invalid_q <= inputs_invalid_d;
    end
   end

  // SEC_CM: KMAC_IF.FSM.SPARSE
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, data_state_e, StIdle)

  always_comb begin
    cnt_clr = 1'b0;
    cnt_set = 1'b0;
    cnt_en  = 1'b0;
    valid   = 1'b0;
    last    = 1'b0;
    strb    = '0;
    done_o  = 1'b0;
    state_d = state_q;
    rounds  = '0;

    clr_err = '0;
    fsm_error_o = '0;
    kmac_error_o = '0;

    kmac_done_vld = '0;

    cmd_chk = 1'b1;

    unique case (state_q)

      StIdle: begin
        // if for some reason multiple bits are set, adv_en has priority
        // as the current key state will be destroyed

        // cross check for commands once transaction begins
        cmd_chk = '0;
        if (start) begin
          cnt_set = 1'b1;
          if (adv_en_i) begin
            rounds = LastAdvRound;
          end else if (id_en_i) begin
            rounds = LastIdRound;
          end else if (gen_en_i) begin
            rounds = LastGenRound;
          end
          // in case we are sending only 1 entry
          state_d = (rounds == 0) ? StTxLast : StTx;
        end
      end

      StTx: begin
        valid = 1'b1;
        strb = {IfBytes{1'b1}};

        // transaction accepted
        if (kmac_data_i.ready) begin
          cnt_en = 1'b1;

          // second to last beat
          if (cnt == CntWidth'(1'b1)) begin
            state_d = StTxLast;
          end
        end

      end

      StTxLast: begin
        valid = 1'b1;
        last = 1'b1;

        if (adv_en_i) begin
          strb = AdvByteMask;
        end else if (id_en_i) begin
          strb = IdByteMask;
        end else if (gen_en_i) begin
          strb = GenByteMask;
        end

        // transaction accepted
        cnt_clr = kmac_data_i.ready;
        state_d = kmac_data_i.ready ? StOpWait : StTxLast;

      end

      StOpWait: begin
        kmac_done_vld = 1'b1;
        if (kmac_data_i.done) begin
          kmac_error_o = kmac_data_i.error;
          done_o = 1'b1;
          state_d = StClean;
        end
      end

      StClean: begin
        cmd_chk = '0;
        done_o = 1'b1;

        // wait for control side to ack done by waiting start de-assertion
        if (!start) begin
          done_o = 1'b0;
          clr_err = 1'b1;
          state_d = StIdle;
        end
      end

      // trigger error
      default: begin
        // This state is terminal
        done_o = 1'b1;
        fsm_error_o = 1'b1;
      end

    endcase // unique case (state_q)

    // unconditional error transitions
    // counter errors may disturb the fsm flow and are
    // treated like fsm errors
    if (cnt_err) begin
      state_d = StError;
      fsm_error_o = 1;
      done_o = 1'b1;
    end
  end

  // when transaction is not complete, populate the data with random
  assign data_o = start && done_o ?
                  {kmac_data_i.digest_share1,
                   kmac_data_i.digest_share0} :
                  {DecoyOutputCopies{entropy_i[0]}};

  // The input invalid check is done whenever transactions are ongoing with kmac
  // once set, it cannot be unset until transactions are fully complete
  always_comb begin
    inputs_invalid_d = inputs_invalid_q;

    if (clr_err) begin
      inputs_invalid_d = '0;
    end else if (valid) begin
      inputs_invalid_d[OpAdvance]  = adv_en_i & (inputs_invalid_i[OpAdvance] |
                                                 inputs_invalid_q[OpAdvance]);
      inputs_invalid_d[OpGenId]    = id_en_i  & (inputs_invalid_i[OpGenId]   |
                                                 inputs_invalid_q[OpGenId]);
      inputs_invalid_d[OpGenSwOut] = gen_en_i & (inputs_invalid_i[OpGenSwOut]|
                                                 inputs_invalid_q[OpGenSwOut]);
      inputs_invalid_d[OpGenHwOut] = gen_en_i & (inputs_invalid_i[OpGenHwOut]|
                                                 inputs_invalid_q[OpGenHwOut]);
    end
  end

  // immediately assert errors
  assign inputs_invalid_o = |inputs_invalid_d;

  logic [CntWidth-1:0] adv_sel, id_sel, gen_sel;
  assign adv_sel = LastAdvRound - cnt;
  assign id_sel = LastIdRound - cnt;
  assign gen_sel = LastGenRound - cnt;

  // The count is maintained as a downcount
  // so a subtract is necessary to send the right byte
  // alternatively we can also reverse the order of the input
  assign decoy_data = {DecoyCopies{entropy_i[1]}};
  always_comb begin
    kmac_data_o.data  = decoy_data;
    if (|cmd_error_o || inputs_invalid_o || fsm_error_o) begin
      kmac_data_o.data  = decoy_data;
    end else if (valid && adv_en_i) begin
      kmac_data_o.data  = adv_data[adv_sel];
    end else if (valid && id_en_i) begin
      kmac_data_o.data  = id_data[id_sel];
    end else if (valid && gen_en_i) begin
      kmac_data_o.data  = gen_data[gen_sel];
    end
  end

  assign kmac_data_o.valid = valid;
  assign kmac_data_o.last  = last;
  assign kmac_data_o.strb  = strb;

  // kmac done is asserted outside of expected window
  // SEC_CM: KMAC_IF_DONE.CTRL.CONSISTENCY
  logic kmac_done_err_q, kmac_done_err_d;
  assign kmac_done_err_d = ~kmac_done_vld & kmac_data_i.done |
                           kmac_done_err_q;
  assign kmac_done_error_o = kmac_done_err_q;


  // the enables must be 1 hot
  logic [2:0] enables_d, enables_q, enables_sub;
  assign enables_d = {adv_en_i, id_en_i, gen_en_i};
  assign enables_sub = enables_d - 1'b1;

  // cross check to ensure the one-hot command that kicked off
  // the transaction remains consistent throughout.
  logic cmd_consty_err_q, cmd_consty_err_d;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      enables_q <= '0;
    end else if (cnt_set) begin
      enables_q <= enables_d;
    end
  end
  assign cmd_consty_err_d = (cmd_chk & (enables_q != enables_d)) |
                            cmd_consty_err_q;

  // if a one hot error occurs, latch onto it permanently
  // SEC_CM: KMAC_IF_CMD.CTRL.CONSISTENCY
  logic one_hot_err_q, one_hot_err_d;
  assign one_hot_err_d = |(enables_d & enables_sub) |
                         one_hot_err_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      one_hot_err_q <= '0;
      kmac_done_err_q <= '0;
      cmd_consty_err_q <= '0;
    end else begin
      one_hot_err_q <= one_hot_err_d;
      kmac_done_err_q <= kmac_done_err_d;
      cmd_consty_err_q <= cmd_consty_err_d;
    end
  end

  // command error occurs if kmac errors or if the command itself is invalid
  assign cmd_error_o = one_hot_err_q | cmd_consty_err_q;

  // request entropy to churn whenever a transaction is accepted
  assign prng_en_o = kmac_data_o.valid & kmac_data_i.ready;

  // as long as we are transmitting, the strobe should never be 0.
  `ASSERT(LastStrb_A, valid |-> strb != '0)


endmodule // keymgr_kmac_if


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager operation state control
//

`include "prim_assert.sv"

module keymgr_op_state_ctrl
  import keymgr_pkg::*;
  import keymgr_reg_pkg::*;
(
  input clk_i,
  input rst_ni,

  input adv_req_i,
  input dis_req_i,
  input id_req_i,
  input gen_req_i,
  input [CdiWidth-1:0] cnt_i,
  output logic op_ack_o,
  output logic op_busy_o,
  output logic op_update_o,

  input kmac_done_i,
  output logic adv_en_o,
  output logic id_en_o,
  output logic gen_en_o,

  output logic op_fsm_err_o

);

  localparam int OpStateWidth = 8;
  typedef enum logic [OpStateWidth-1:0] {
    StIdle   = 8'b10010101,
    StAdv    = 8'b00101000,
    StAdvAck = 8'b01000011,
    StWait   = 8'b11111110
  } state_e;

  state_e state_q, state_d;
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, StIdle)

  logic gen_en;
  assign id_en_o = gen_en & id_req_i;
  assign gen_en_o = gen_en & gen_req_i;

  always_comb begin
    state_d = state_q;
    op_update_o = 1'b0;
    op_ack_o = 1'b0;
    op_busy_o = 1'b1;

    // output to kmac interface
    adv_en_o = 1'b0;

    gen_en = 1'b0;
    op_fsm_err_o = 1'b0;

    unique case (state_q)
      StIdle: begin
        op_busy_o = '0;
        if (adv_req_i || dis_req_i) begin
          state_d = StAdv;
        end else if (id_req_i || gen_req_i) begin
          state_d = StWait;
        end
      end

      StAdv: begin
        adv_en_o = 1'b1;

        if (kmac_done_i && (int'(cnt_i) == CDIs-1)) begin
          op_ack_o = 1'b1;
          state_d = StIdle;
        end else if (kmac_done_i && (int'(cnt_i) < CDIs-1)) begin
          op_update_o = 1'b1;
          state_d = StAdvAck;
        end
      end

      // drop adv_en_o to allow kmac interface handshake
      StAdvAck: begin
        state_d = StAdv;
      end

      // Not an advanced operation
      StWait: begin
        gen_en = 1'b1;

        if (kmac_done_i) begin
          op_ack_o = 1'b1;
          state_d = StIdle;
        end
      end

      // error state
      default: begin
        // allow completion of transaction
        op_ack_o = 1'b1;
        op_fsm_err_o = 1'b1;
      end

    endcase // unique case (adv_state_q)
  end


endmodule // keymgr_op_state_ctrl


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module keymgr_reg_top (
  input clk_i,
  input rst_ni,
  input rst_shadowed_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output keymgr_reg_pkg::keymgr_reg2hw_t reg2hw, // Write
  input  keymgr_reg_pkg::keymgr_hw2reg_t hw2reg, // Read

  output logic shadowed_storage_err_o,
  output logic shadowed_update_err_o,

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import keymgr_reg_pkg::* ;

  localparam int AW = 8;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [62:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(63)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_qs;
  logic intr_state_wd;
  logic intr_enable_we;
  logic intr_enable_qs;
  logic intr_enable_wd;
  logic intr_test_we;
  logic intr_test_wd;
  logic alert_test_we;
  logic alert_test_recov_operation_err_wd;
  logic alert_test_fatal_fault_err_wd;
  logic cfg_regwen_re;
  logic cfg_regwen_qs;
  logic start_we;
  logic start_qs;
  logic start_wd;
  logic control_shadowed_re;
  logic control_shadowed_we;
  logic [2:0] control_shadowed_operation_qs;
  logic [2:0] control_shadowed_operation_wd;
  logic control_shadowed_operation_storage_err;
  logic control_shadowed_operation_update_err;
  logic control_shadowed_cdi_sel_qs;
  logic control_shadowed_cdi_sel_wd;
  logic control_shadowed_cdi_sel_storage_err;
  logic control_shadowed_cdi_sel_update_err;
  logic [1:0] control_shadowed_dest_sel_qs;
  logic [1:0] control_shadowed_dest_sel_wd;
  logic control_shadowed_dest_sel_storage_err;
  logic control_shadowed_dest_sel_update_err;
  logic sideload_clear_we;
  logic [2:0] sideload_clear_qs;
  logic [2:0] sideload_clear_wd;
  logic reseed_interval_regwen_we;
  logic reseed_interval_regwen_qs;
  logic reseed_interval_regwen_wd;
  logic reseed_interval_shadowed_re;
  logic reseed_interval_shadowed_we;
  logic [15:0] reseed_interval_shadowed_qs;
  logic [15:0] reseed_interval_shadowed_wd;
  logic reseed_interval_shadowed_storage_err;
  logic reseed_interval_shadowed_update_err;
  logic sw_binding_regwen_re;
  logic sw_binding_regwen_we;
  logic sw_binding_regwen_qs;
  logic sw_binding_regwen_wd;
  logic sealing_sw_binding_0_we;
  logic [31:0] sealing_sw_binding_0_qs;
  logic [31:0] sealing_sw_binding_0_wd;
  logic sealing_sw_binding_1_we;
  logic [31:0] sealing_sw_binding_1_qs;
  logic [31:0] sealing_sw_binding_1_wd;
  logic sealing_sw_binding_2_we;
  logic [31:0] sealing_sw_binding_2_qs;
  logic [31:0] sealing_sw_binding_2_wd;
  logic sealing_sw_binding_3_we;
  logic [31:0] sealing_sw_binding_3_qs;
  logic [31:0] sealing_sw_binding_3_wd;
  logic sealing_sw_binding_4_we;
  logic [31:0] sealing_sw_binding_4_qs;
  logic [31:0] sealing_sw_binding_4_wd;
  logic sealing_sw_binding_5_we;
  logic [31:0] sealing_sw_binding_5_qs;
  logic [31:0] sealing_sw_binding_5_wd;
  logic sealing_sw_binding_6_we;
  logic [31:0] sealing_sw_binding_6_qs;
  logic [31:0] sealing_sw_binding_6_wd;
  logic sealing_sw_binding_7_we;
  logic [31:0] sealing_sw_binding_7_qs;
  logic [31:0] sealing_sw_binding_7_wd;
  logic attest_sw_binding_0_we;
  logic [31:0] attest_sw_binding_0_qs;
  logic [31:0] attest_sw_binding_0_wd;
  logic attest_sw_binding_1_we;
  logic [31:0] attest_sw_binding_1_qs;
  logic [31:0] attest_sw_binding_1_wd;
  logic attest_sw_binding_2_we;
  logic [31:0] attest_sw_binding_2_qs;
  logic [31:0] attest_sw_binding_2_wd;
  logic attest_sw_binding_3_we;
  logic [31:0] attest_sw_binding_3_qs;
  logic [31:0] attest_sw_binding_3_wd;
  logic attest_sw_binding_4_we;
  logic [31:0] attest_sw_binding_4_qs;
  logic [31:0] attest_sw_binding_4_wd;
  logic attest_sw_binding_5_we;
  logic [31:0] attest_sw_binding_5_qs;
  logic [31:0] attest_sw_binding_5_wd;
  logic attest_sw_binding_6_we;
  logic [31:0] attest_sw_binding_6_qs;
  logic [31:0] attest_sw_binding_6_wd;
  logic attest_sw_binding_7_we;
  logic [31:0] attest_sw_binding_7_qs;
  logic [31:0] attest_sw_binding_7_wd;
  logic salt_0_we;
  logic [31:0] salt_0_qs;
  logic [31:0] salt_0_wd;
  logic salt_1_we;
  logic [31:0] salt_1_qs;
  logic [31:0] salt_1_wd;
  logic salt_2_we;
  logic [31:0] salt_2_qs;
  logic [31:0] salt_2_wd;
  logic salt_3_we;
  logic [31:0] salt_3_qs;
  logic [31:0] salt_3_wd;
  logic salt_4_we;
  logic [31:0] salt_4_qs;
  logic [31:0] salt_4_wd;
  logic salt_5_we;
  logic [31:0] salt_5_qs;
  logic [31:0] salt_5_wd;
  logic salt_6_we;
  logic [31:0] salt_6_qs;
  logic [31:0] salt_6_wd;
  logic salt_7_we;
  logic [31:0] salt_7_qs;
  logic [31:0] salt_7_wd;
  logic key_version_we;
  logic [31:0] key_version_qs;
  logic [31:0] key_version_wd;
  logic max_creator_key_ver_regwen_we;
  logic max_creator_key_ver_regwen_qs;
  logic max_creator_key_ver_regwen_wd;
  logic max_creator_key_ver_shadowed_re;
  logic max_creator_key_ver_shadowed_we;
  logic [31:0] max_creator_key_ver_shadowed_qs;
  logic [31:0] max_creator_key_ver_shadowed_wd;
  logic max_creator_key_ver_shadowed_storage_err;
  logic max_creator_key_ver_shadowed_update_err;
  logic max_owner_int_key_ver_regwen_we;
  logic max_owner_int_key_ver_regwen_qs;
  logic max_owner_int_key_ver_regwen_wd;
  logic max_owner_int_key_ver_shadowed_re;
  logic max_owner_int_key_ver_shadowed_we;
  logic [31:0] max_owner_int_key_ver_shadowed_qs;
  logic [31:0] max_owner_int_key_ver_shadowed_wd;
  logic max_owner_int_key_ver_shadowed_storage_err;
  logic max_owner_int_key_ver_shadowed_update_err;
  logic max_owner_key_ver_regwen_we;
  logic max_owner_key_ver_regwen_qs;
  logic max_owner_key_ver_regwen_wd;
  logic max_owner_key_ver_shadowed_re;
  logic max_owner_key_ver_shadowed_we;
  logic [31:0] max_owner_key_ver_shadowed_qs;
  logic [31:0] max_owner_key_ver_shadowed_wd;
  logic max_owner_key_ver_shadowed_storage_err;
  logic max_owner_key_ver_shadowed_update_err;
  logic sw_share0_output_0_re;
  logic [31:0] sw_share0_output_0_qs;
  logic [31:0] sw_share0_output_0_wd;
  logic sw_share0_output_1_re;
  logic [31:0] sw_share0_output_1_qs;
  logic [31:0] sw_share0_output_1_wd;
  logic sw_share0_output_2_re;
  logic [31:0] sw_share0_output_2_qs;
  logic [31:0] sw_share0_output_2_wd;
  logic sw_share0_output_3_re;
  logic [31:0] sw_share0_output_3_qs;
  logic [31:0] sw_share0_output_3_wd;
  logic sw_share0_output_4_re;
  logic [31:0] sw_share0_output_4_qs;
  logic [31:0] sw_share0_output_4_wd;
  logic sw_share0_output_5_re;
  logic [31:0] sw_share0_output_5_qs;
  logic [31:0] sw_share0_output_5_wd;
  logic sw_share0_output_6_re;
  logic [31:0] sw_share0_output_6_qs;
  logic [31:0] sw_share0_output_6_wd;
  logic sw_share0_output_7_re;
  logic [31:0] sw_share0_output_7_qs;
  logic [31:0] sw_share0_output_7_wd;
  logic sw_share1_output_0_re;
  logic [31:0] sw_share1_output_0_qs;
  logic [31:0] sw_share1_output_0_wd;
  logic sw_share1_output_1_re;
  logic [31:0] sw_share1_output_1_qs;
  logic [31:0] sw_share1_output_1_wd;
  logic sw_share1_output_2_re;
  logic [31:0] sw_share1_output_2_qs;
  logic [31:0] sw_share1_output_2_wd;
  logic sw_share1_output_3_re;
  logic [31:0] sw_share1_output_3_qs;
  logic [31:0] sw_share1_output_3_wd;
  logic sw_share1_output_4_re;
  logic [31:0] sw_share1_output_4_qs;
  logic [31:0] sw_share1_output_4_wd;
  logic sw_share1_output_5_re;
  logic [31:0] sw_share1_output_5_qs;
  logic [31:0] sw_share1_output_5_wd;
  logic sw_share1_output_6_re;
  logic [31:0] sw_share1_output_6_qs;
  logic [31:0] sw_share1_output_6_wd;
  logic sw_share1_output_7_re;
  logic [31:0] sw_share1_output_7_qs;
  logic [31:0] sw_share1_output_7_wd;
  logic [2:0] working_state_qs;
  logic op_status_we;
  logic [1:0] op_status_qs;
  logic [1:0] op_status_wd;
  logic err_code_we;
  logic err_code_invalid_op_qs;
  logic err_code_invalid_op_wd;
  logic err_code_invalid_kmac_input_qs;
  logic err_code_invalid_kmac_input_wd;
  logic err_code_invalid_shadow_update_qs;
  logic err_code_invalid_shadow_update_wd;
  logic fault_status_cmd_qs;
  logic fault_status_kmac_fsm_qs;
  logic fault_status_kmac_done_qs;
  logic fault_status_kmac_op_qs;
  logic fault_status_kmac_out_qs;
  logic fault_status_regfile_intg_qs;
  logic fault_status_shadow_qs;
  logic fault_status_ctrl_fsm_intg_qs;
  logic fault_status_ctrl_fsm_chk_qs;
  logic fault_status_ctrl_fsm_cnt_qs;
  logic fault_status_reseed_cnt_qs;
  logic fault_status_side_ctrl_fsm_qs;
  logic fault_status_side_ctrl_sel_qs;
  logic fault_status_key_ecc_qs;
  logic debug_we;
  logic debug_invalid_creator_seed_qs;
  logic debug_invalid_creator_seed_wd;
  logic debug_invalid_owner_seed_qs;
  logic debug_invalid_owner_seed_wd;
  logic debug_invalid_dev_id_qs;
  logic debug_invalid_dev_id_wd;
  logic debug_invalid_health_state_qs;
  logic debug_invalid_health_state_wd;
  logic debug_invalid_key_version_qs;
  logic debug_invalid_key_version_wd;
  logic debug_invalid_key_qs;
  logic debug_invalid_key_wd;
  logic debug_invalid_digest_qs;
  logic debug_invalid_digest_wd;

  // Register instances
  // R[intr_state]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.de),
    .d      (hw2reg.intr_state.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_qs)
  );


  // R[intr_enable]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [0:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[recov_operation_err]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov_operation_err (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_operation_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.recov_operation_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov_operation_err.qe = alert_test_qe;

  //   F[fatal_fault_err]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal_fault_err (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_fault_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.fatal_fault_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal_fault_err.qe = alert_test_qe;


  // R[cfg_regwen]: V(True)
  prim_subreg_ext #(
    .DW    (1)
  ) u_cfg_regwen (
    .re     (cfg_regwen_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.cfg_regwen.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (cfg_regwen_qs)
  );


  // R[start]: V(False)
  // Create REGWEN-gated WE signal
  logic start_gated_we;
  assign start_gated_we = start_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_start (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (start_gated_we),
    .wd     (start_wd),

    // from internal hardware
    .de     (hw2reg.start.de),
    .d      (hw2reg.start.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.start.q),
    .ds     (),

    // to register interface (read)
    .qs     (start_qs)
  );


  // R[control_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic control_shadowed_gated_we;
  assign control_shadowed_gated_we = control_shadowed_we & cfg_regwen_qs;
  //   F[operation]: 6:4
  prim_subreg_shadow #(
    .DW      (3),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (3'h1)
  ) u_control_shadowed_operation (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (control_shadowed_re),
    .we     (control_shadowed_gated_we),
    .wd     (control_shadowed_operation_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.control_shadowed.operation.q),
    .ds     (),

    // to register interface (read)
    .qs     (control_shadowed_operation_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (control_shadowed_operation_update_err),
    .err_storage (control_shadowed_operation_storage_err)
  );

  //   F[cdi_sel]: 7:7
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_control_shadowed_cdi_sel (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (control_shadowed_re),
    .we     (control_shadowed_gated_we),
    .wd     (control_shadowed_cdi_sel_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.control_shadowed.cdi_sel.q),
    .ds     (),

    // to register interface (read)
    .qs     (control_shadowed_cdi_sel_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (control_shadowed_cdi_sel_update_err),
    .err_storage (control_shadowed_cdi_sel_storage_err)
  );

  //   F[dest_sel]: 13:12
  prim_subreg_shadow #(
    .DW      (2),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (2'h0)
  ) u_control_shadowed_dest_sel (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (control_shadowed_re),
    .we     (control_shadowed_gated_we),
    .wd     (control_shadowed_dest_sel_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.control_shadowed.dest_sel.q),
    .ds     (),

    // to register interface (read)
    .qs     (control_shadowed_dest_sel_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (control_shadowed_dest_sel_update_err),
    .err_storage (control_shadowed_dest_sel_storage_err)
  );


  // R[sideload_clear]: V(False)
  // Create REGWEN-gated WE signal
  logic sideload_clear_gated_we;
  assign sideload_clear_gated_we = sideload_clear_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (3),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (3'h0)
  ) u_sideload_clear (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sideload_clear_gated_we),
    .wd     (sideload_clear_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sideload_clear.q),
    .ds     (),

    // to register interface (read)
    .qs     (sideload_clear_qs)
  );


  // R[reseed_interval_regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_reseed_interval_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (reseed_interval_regwen_we),
    .wd     (reseed_interval_regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (reseed_interval_regwen_qs)
  );


  // R[reseed_interval_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic reseed_interval_shadowed_gated_we;
  assign reseed_interval_shadowed_gated_we =
    reseed_interval_shadowed_we & reseed_interval_regwen_qs;
  prim_subreg_shadow #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h100)
  ) u_reseed_interval_shadowed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (reseed_interval_shadowed_re),
    .we     (reseed_interval_shadowed_gated_we),
    .wd     (reseed_interval_shadowed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.reseed_interval_shadowed.q),
    .ds     (),

    // to register interface (read)
    .qs     (reseed_interval_shadowed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (reseed_interval_shadowed_update_err),
    .err_storage (reseed_interval_shadowed_storage_err)
  );


  // R[sw_binding_regwen]: V(True)
  logic sw_binding_regwen_qe;
  logic [0:0] sw_binding_regwen_flds_we;
  assign sw_binding_regwen_qe = &sw_binding_regwen_flds_we;
  prim_subreg_ext #(
    .DW    (1)
  ) u_sw_binding_regwen (
    .re     (sw_binding_regwen_re),
    .we     (sw_binding_regwen_we),
    .wd     (sw_binding_regwen_wd),
    .d      (hw2reg.sw_binding_regwen.d),
    .qre    (),
    .qe     (sw_binding_regwen_flds_we[0]),
    .q      (reg2hw.sw_binding_regwen.q),
    .ds     (),
    .qs     (sw_binding_regwen_qs)
  );
  assign reg2hw.sw_binding_regwen.qe = sw_binding_regwen_qe;


  // Subregister 0 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_0]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_0_gated_we;
  assign sealing_sw_binding_0_gated_we = sealing_sw_binding_0_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_0_gated_we),
    .wd     (sealing_sw_binding_0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_0_qs)
  );


  // Subregister 1 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_1]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_1_gated_we;
  assign sealing_sw_binding_1_gated_we = sealing_sw_binding_1_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_1_gated_we),
    .wd     (sealing_sw_binding_1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_1_qs)
  );


  // Subregister 2 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_2]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_2_gated_we;
  assign sealing_sw_binding_2_gated_we = sealing_sw_binding_2_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_2_gated_we),
    .wd     (sealing_sw_binding_2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_2_qs)
  );


  // Subregister 3 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_3]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_3_gated_we;
  assign sealing_sw_binding_3_gated_we = sealing_sw_binding_3_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_3_gated_we),
    .wd     (sealing_sw_binding_3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_3_qs)
  );


  // Subregister 4 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_4]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_4_gated_we;
  assign sealing_sw_binding_4_gated_we = sealing_sw_binding_4_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_4_gated_we),
    .wd     (sealing_sw_binding_4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_4_qs)
  );


  // Subregister 5 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_5]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_5_gated_we;
  assign sealing_sw_binding_5_gated_we = sealing_sw_binding_5_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_5_gated_we),
    .wd     (sealing_sw_binding_5_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_5_qs)
  );


  // Subregister 6 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_6]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_6_gated_we;
  assign sealing_sw_binding_6_gated_we = sealing_sw_binding_6_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_6_gated_we),
    .wd     (sealing_sw_binding_6_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_6_qs)
  );


  // Subregister 7 of Multireg sealing_sw_binding
  // R[sealing_sw_binding_7]: V(False)
  // Create REGWEN-gated WE signal
  logic sealing_sw_binding_7_gated_we;
  assign sealing_sw_binding_7_gated_we = sealing_sw_binding_7_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_sealing_sw_binding_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sealing_sw_binding_7_gated_we),
    .wd     (sealing_sw_binding_7_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.sealing_sw_binding[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (sealing_sw_binding_7_qs)
  );


  // Subregister 0 of Multireg attest_sw_binding
  // R[attest_sw_binding_0]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_0_gated_we;
  assign attest_sw_binding_0_gated_we = attest_sw_binding_0_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_0_gated_we),
    .wd     (attest_sw_binding_0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_0_qs)
  );


  // Subregister 1 of Multireg attest_sw_binding
  // R[attest_sw_binding_1]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_1_gated_we;
  assign attest_sw_binding_1_gated_we = attest_sw_binding_1_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_1_gated_we),
    .wd     (attest_sw_binding_1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_1_qs)
  );


  // Subregister 2 of Multireg attest_sw_binding
  // R[attest_sw_binding_2]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_2_gated_we;
  assign attest_sw_binding_2_gated_we = attest_sw_binding_2_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_2_gated_we),
    .wd     (attest_sw_binding_2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_2_qs)
  );


  // Subregister 3 of Multireg attest_sw_binding
  // R[attest_sw_binding_3]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_3_gated_we;
  assign attest_sw_binding_3_gated_we = attest_sw_binding_3_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_3_gated_we),
    .wd     (attest_sw_binding_3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_3_qs)
  );


  // Subregister 4 of Multireg attest_sw_binding
  // R[attest_sw_binding_4]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_4_gated_we;
  assign attest_sw_binding_4_gated_we = attest_sw_binding_4_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_4_gated_we),
    .wd     (attest_sw_binding_4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_4_qs)
  );


  // Subregister 5 of Multireg attest_sw_binding
  // R[attest_sw_binding_5]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_5_gated_we;
  assign attest_sw_binding_5_gated_we = attest_sw_binding_5_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_5_gated_we),
    .wd     (attest_sw_binding_5_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_5_qs)
  );


  // Subregister 6 of Multireg attest_sw_binding
  // R[attest_sw_binding_6]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_6_gated_we;
  assign attest_sw_binding_6_gated_we = attest_sw_binding_6_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_6_gated_we),
    .wd     (attest_sw_binding_6_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_6_qs)
  );


  // Subregister 7 of Multireg attest_sw_binding
  // R[attest_sw_binding_7]: V(False)
  // Create REGWEN-gated WE signal
  logic attest_sw_binding_7_gated_we;
  assign attest_sw_binding_7_gated_we = attest_sw_binding_7_we & sw_binding_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_attest_sw_binding_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (attest_sw_binding_7_gated_we),
    .wd     (attest_sw_binding_7_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.attest_sw_binding[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (attest_sw_binding_7_qs)
  );


  // Subregister 0 of Multireg salt
  // R[salt_0]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_0_gated_we;
  assign salt_0_gated_we = salt_0_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_0_gated_we),
    .wd     (salt_0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_0_qs)
  );


  // Subregister 1 of Multireg salt
  // R[salt_1]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_1_gated_we;
  assign salt_1_gated_we = salt_1_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_1_gated_we),
    .wd     (salt_1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_1_qs)
  );


  // Subregister 2 of Multireg salt
  // R[salt_2]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_2_gated_we;
  assign salt_2_gated_we = salt_2_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_2_gated_we),
    .wd     (salt_2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_2_qs)
  );


  // Subregister 3 of Multireg salt
  // R[salt_3]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_3_gated_we;
  assign salt_3_gated_we = salt_3_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_3_gated_we),
    .wd     (salt_3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_3_qs)
  );


  // Subregister 4 of Multireg salt
  // R[salt_4]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_4_gated_we;
  assign salt_4_gated_we = salt_4_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_4_gated_we),
    .wd     (salt_4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_4_qs)
  );


  // Subregister 5 of Multireg salt
  // R[salt_5]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_5_gated_we;
  assign salt_5_gated_we = salt_5_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_5_gated_we),
    .wd     (salt_5_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_5_qs)
  );


  // Subregister 6 of Multireg salt
  // R[salt_6]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_6_gated_we;
  assign salt_6_gated_we = salt_6_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_6_gated_we),
    .wd     (salt_6_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_6_qs)
  );


  // Subregister 7 of Multireg salt
  // R[salt_7]: V(False)
  // Create REGWEN-gated WE signal
  logic salt_7_gated_we;
  assign salt_7_gated_we = salt_7_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_salt_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (salt_7_gated_we),
    .wd     (salt_7_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.salt[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (salt_7_qs)
  );


  // Subregister 0 of Multireg key_version
  // R[key_version]: V(False)
  // Create REGWEN-gated WE signal
  logic key_version_gated_we;
  assign key_version_gated_we = key_version_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_key_version (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (key_version_gated_we),
    .wd     (key_version_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.key_version[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (key_version_qs)
  );


  // R[max_creator_key_ver_regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_max_creator_key_ver_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (max_creator_key_ver_regwen_we),
    .wd     (max_creator_key_ver_regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (max_creator_key_ver_regwen_qs)
  );


  // R[max_creator_key_ver_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic max_creator_key_ver_shadowed_gated_we;
  assign max_creator_key_ver_shadowed_gated_we =
    max_creator_key_ver_shadowed_we & max_creator_key_ver_regwen_qs;
  prim_subreg_shadow #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_max_creator_key_ver_shadowed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (max_creator_key_ver_shadowed_re),
    .we     (max_creator_key_ver_shadowed_gated_we),
    .wd     (max_creator_key_ver_shadowed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.max_creator_key_ver_shadowed.q),
    .ds     (),

    // to register interface (read)
    .qs     (max_creator_key_ver_shadowed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (max_creator_key_ver_shadowed_update_err),
    .err_storage (max_creator_key_ver_shadowed_storage_err)
  );


  // R[max_owner_int_key_ver_regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_max_owner_int_key_ver_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (max_owner_int_key_ver_regwen_we),
    .wd     (max_owner_int_key_ver_regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (max_owner_int_key_ver_regwen_qs)
  );


  // R[max_owner_int_key_ver_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic max_owner_int_key_ver_shadowed_gated_we;
  assign max_owner_int_key_ver_shadowed_gated_we =
    max_owner_int_key_ver_shadowed_we & max_owner_int_key_ver_regwen_qs;
  prim_subreg_shadow #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h1)
  ) u_max_owner_int_key_ver_shadowed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (max_owner_int_key_ver_shadowed_re),
    .we     (max_owner_int_key_ver_shadowed_gated_we),
    .wd     (max_owner_int_key_ver_shadowed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.max_owner_int_key_ver_shadowed.q),
    .ds     (),

    // to register interface (read)
    .qs     (max_owner_int_key_ver_shadowed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (max_owner_int_key_ver_shadowed_update_err),
    .err_storage (max_owner_int_key_ver_shadowed_storage_err)
  );


  // R[max_owner_key_ver_regwen]: V(False)
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h1)
  ) u_max_owner_key_ver_regwen (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (max_owner_key_ver_regwen_we),
    .wd     (max_owner_key_ver_regwen_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (max_owner_key_ver_regwen_qs)
  );


  // R[max_owner_key_ver_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic max_owner_key_ver_shadowed_gated_we;
  assign max_owner_key_ver_shadowed_gated_we =
    max_owner_key_ver_shadowed_we & max_owner_key_ver_regwen_qs;
  prim_subreg_shadow #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_max_owner_key_ver_shadowed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (max_owner_key_ver_shadowed_re),
    .we     (max_owner_key_ver_shadowed_gated_we),
    .wd     (max_owner_key_ver_shadowed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.max_owner_key_ver_shadowed.q),
    .ds     (),

    // to register interface (read)
    .qs     (max_owner_key_ver_shadowed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (max_owner_key_ver_shadowed_update_err),
    .err_storage (max_owner_key_ver_shadowed_storage_err)
  );


  // Subregister 0 of Multireg sw_share0_output
  // R[sw_share0_output_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_0_re),
    .wd     (sw_share0_output_0_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[0].de),
    .d      (hw2reg.sw_share0_output[0].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_0_qs)
  );


  // Subregister 1 of Multireg sw_share0_output
  // R[sw_share0_output_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_1_re),
    .wd     (sw_share0_output_1_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[1].de),
    .d      (hw2reg.sw_share0_output[1].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_1_qs)
  );


  // Subregister 2 of Multireg sw_share0_output
  // R[sw_share0_output_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_2_re),
    .wd     (sw_share0_output_2_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[2].de),
    .d      (hw2reg.sw_share0_output[2].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_2_qs)
  );


  // Subregister 3 of Multireg sw_share0_output
  // R[sw_share0_output_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_3_re),
    .wd     (sw_share0_output_3_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[3].de),
    .d      (hw2reg.sw_share0_output[3].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_3_qs)
  );


  // Subregister 4 of Multireg sw_share0_output
  // R[sw_share0_output_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_4_re),
    .wd     (sw_share0_output_4_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[4].de),
    .d      (hw2reg.sw_share0_output[4].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_4_qs)
  );


  // Subregister 5 of Multireg sw_share0_output
  // R[sw_share0_output_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_5_re),
    .wd     (sw_share0_output_5_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[5].de),
    .d      (hw2reg.sw_share0_output[5].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_5_qs)
  );


  // Subregister 6 of Multireg sw_share0_output
  // R[sw_share0_output_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_6_re),
    .wd     (sw_share0_output_6_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[6].de),
    .d      (hw2reg.sw_share0_output[6].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_6_qs)
  );


  // Subregister 7 of Multireg sw_share0_output
  // R[sw_share0_output_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share0_output_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share0_output_7_re),
    .wd     (sw_share0_output_7_wd),

    // from internal hardware
    .de     (hw2reg.sw_share0_output[7].de),
    .d      (hw2reg.sw_share0_output[7].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share0_output_7_qs)
  );


  // Subregister 0 of Multireg sw_share1_output
  // R[sw_share1_output_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_0_re),
    .wd     (sw_share1_output_0_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[0].de),
    .d      (hw2reg.sw_share1_output[0].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_0_qs)
  );


  // Subregister 1 of Multireg sw_share1_output
  // R[sw_share1_output_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_1_re),
    .wd     (sw_share1_output_1_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[1].de),
    .d      (hw2reg.sw_share1_output[1].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_1_qs)
  );


  // Subregister 2 of Multireg sw_share1_output
  // R[sw_share1_output_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_2_re),
    .wd     (sw_share1_output_2_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[2].de),
    .d      (hw2reg.sw_share1_output[2].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_2_qs)
  );


  // Subregister 3 of Multireg sw_share1_output
  // R[sw_share1_output_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_3_re),
    .wd     (sw_share1_output_3_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[3].de),
    .d      (hw2reg.sw_share1_output[3].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_3_qs)
  );


  // Subregister 4 of Multireg sw_share1_output
  // R[sw_share1_output_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_4_re),
    .wd     (sw_share1_output_4_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[4].de),
    .d      (hw2reg.sw_share1_output[4].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_4_qs)
  );


  // Subregister 5 of Multireg sw_share1_output
  // R[sw_share1_output_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_5_re),
    .wd     (sw_share1_output_5_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[5].de),
    .d      (hw2reg.sw_share1_output[5].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_5_qs)
  );


  // Subregister 6 of Multireg sw_share1_output
  // R[sw_share1_output_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_6_re),
    .wd     (sw_share1_output_6_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[6].de),
    .d      (hw2reg.sw_share1_output[6].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_6_qs)
  );


  // Subregister 7 of Multireg sw_share1_output
  // R[sw_share1_output_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRC),
    .RESVAL  (32'h0)
  ) u_sw_share1_output_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (sw_share1_output_7_re),
    .wd     (sw_share1_output_7_wd),

    // from internal hardware
    .de     (hw2reg.sw_share1_output[7].de),
    .d      (hw2reg.sw_share1_output[7].d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (sw_share1_output_7_qs)
  );


  // R[working_state]: V(False)
  prim_subreg #(
    .DW      (3),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (3'h0)
  ) u_working_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.working_state.de),
    .d      (hw2reg.working_state.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (working_state_qs)
  );


  // R[op_status]: V(False)
  prim_subreg #(
    .DW      (2),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (2'h0)
  ) u_op_status (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (op_status_we),
    .wd     (op_status_wd),

    // from internal hardware
    .de     (hw2reg.op_status.de),
    .d      (hw2reg.op_status.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (op_status_qs)
  );


  // R[err_code]: V(False)
  //   F[invalid_op]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_err_code_invalid_op (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (err_code_we),
    .wd     (err_code_invalid_op_wd),

    // from internal hardware
    .de     (hw2reg.err_code.invalid_op.de),
    .d      (hw2reg.err_code.invalid_op.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_invalid_op_qs)
  );

  //   F[invalid_kmac_input]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_err_code_invalid_kmac_input (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (err_code_we),
    .wd     (err_code_invalid_kmac_input_wd),

    // from internal hardware
    .de     (hw2reg.err_code.invalid_kmac_input.de),
    .d      (hw2reg.err_code.invalid_kmac_input.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_invalid_kmac_input_qs)
  );

  //   F[invalid_shadow_update]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_err_code_invalid_shadow_update (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (err_code_we),
    .wd     (err_code_invalid_shadow_update_wd),

    // from internal hardware
    .de     (hw2reg.err_code.invalid_shadow_update.de),
    .d      (hw2reg.err_code.invalid_shadow_update.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_invalid_shadow_update_qs)
  );


  // R[fault_status]: V(False)
  //   F[cmd]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_cmd (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.cmd.de),
    .d      (hw2reg.fault_status.cmd.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.cmd.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_cmd_qs)
  );

  //   F[kmac_fsm]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_kmac_fsm (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.kmac_fsm.de),
    .d      (hw2reg.fault_status.kmac_fsm.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.kmac_fsm.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_kmac_fsm_qs)
  );

  //   F[kmac_done]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_kmac_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.kmac_done.de),
    .d      (hw2reg.fault_status.kmac_done.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.kmac_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_kmac_done_qs)
  );

  //   F[kmac_op]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_kmac_op (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.kmac_op.de),
    .d      (hw2reg.fault_status.kmac_op.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.kmac_op.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_kmac_op_qs)
  );

  //   F[kmac_out]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_kmac_out (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.kmac_out.de),
    .d      (hw2reg.fault_status.kmac_out.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.kmac_out.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_kmac_out_qs)
  );

  //   F[regfile_intg]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_regfile_intg (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.regfile_intg.de),
    .d      (hw2reg.fault_status.regfile_intg.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.regfile_intg.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_regfile_intg_qs)
  );

  //   F[shadow]: 6:6
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_shadow (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.shadow.de),
    .d      (hw2reg.fault_status.shadow.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.shadow.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_shadow_qs)
  );

  //   F[ctrl_fsm_intg]: 7:7
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_ctrl_fsm_intg (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.ctrl_fsm_intg.de),
    .d      (hw2reg.fault_status.ctrl_fsm_intg.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.ctrl_fsm_intg.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_ctrl_fsm_intg_qs)
  );

  //   F[ctrl_fsm_chk]: 8:8
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_ctrl_fsm_chk (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.ctrl_fsm_chk.de),
    .d      (hw2reg.fault_status.ctrl_fsm_chk.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.ctrl_fsm_chk.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_ctrl_fsm_chk_qs)
  );

  //   F[ctrl_fsm_cnt]: 9:9
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_ctrl_fsm_cnt (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.ctrl_fsm_cnt.de),
    .d      (hw2reg.fault_status.ctrl_fsm_cnt.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.ctrl_fsm_cnt.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_ctrl_fsm_cnt_qs)
  );

  //   F[reseed_cnt]: 10:10
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_reseed_cnt (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.reseed_cnt.de),
    .d      (hw2reg.fault_status.reseed_cnt.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.reseed_cnt.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_reseed_cnt_qs)
  );

  //   F[side_ctrl_fsm]: 11:11
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_side_ctrl_fsm (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.side_ctrl_fsm.de),
    .d      (hw2reg.fault_status.side_ctrl_fsm.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.side_ctrl_fsm.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_side_ctrl_fsm_qs)
  );

  //   F[side_ctrl_sel]: 12:12
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_side_ctrl_sel (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.side_ctrl_sel.de),
    .d      (hw2reg.fault_status.side_ctrl_sel.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.side_ctrl_sel.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_side_ctrl_sel_qs)
  );

  //   F[key_ecc]: 13:13
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fault_status_key_ecc (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fault_status.key_ecc.de),
    .d      (hw2reg.fault_status.key_ecc.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.fault_status.key_ecc.q),
    .ds     (),

    // to register interface (read)
    .qs     (fault_status_key_ecc_qs)
  );


  // R[debug]: V(False)
  //   F[invalid_creator_seed]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_creator_seed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_creator_seed_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_creator_seed.de),
    .d      (hw2reg.debug.invalid_creator_seed.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_creator_seed_qs)
  );

  //   F[invalid_owner_seed]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_owner_seed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_owner_seed_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_owner_seed.de),
    .d      (hw2reg.debug.invalid_owner_seed.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_owner_seed_qs)
  );

  //   F[invalid_dev_id]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_dev_id (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_dev_id_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_dev_id.de),
    .d      (hw2reg.debug.invalid_dev_id.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_dev_id_qs)
  );

  //   F[invalid_health_state]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_health_state (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_health_state_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_health_state.de),
    .d      (hw2reg.debug.invalid_health_state.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_health_state_qs)
  );

  //   F[invalid_key_version]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_key_version (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_key_version_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_key_version.de),
    .d      (hw2reg.debug.invalid_key_version.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_key_version_qs)
  );

  //   F[invalid_key]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_key (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_key_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_key.de),
    .d      (hw2reg.debug.invalid_key.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_key_qs)
  );

  //   F[invalid_digest]: 6:6
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW0C),
    .RESVAL  (1'h0)
  ) u_debug_invalid_digest (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (debug_we),
    .wd     (debug_invalid_digest_wd),

    // from internal hardware
    .de     (hw2reg.debug.invalid_digest.de),
    .d      (hw2reg.debug.invalid_digest.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (debug_invalid_digest_qs)
  );



  logic [62:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == KEYMGR_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == KEYMGR_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == KEYMGR_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == KEYMGR_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == KEYMGR_CFG_REGWEN_OFFSET);
    addr_hit[ 5] = (reg_addr == KEYMGR_START_OFFSET);
    addr_hit[ 6] = (reg_addr == KEYMGR_CONTROL_SHADOWED_OFFSET);
    addr_hit[ 7] = (reg_addr == KEYMGR_SIDELOAD_CLEAR_OFFSET);
    addr_hit[ 8] = (reg_addr == KEYMGR_RESEED_INTERVAL_REGWEN_OFFSET);
    addr_hit[ 9] = (reg_addr == KEYMGR_RESEED_INTERVAL_SHADOWED_OFFSET);
    addr_hit[10] = (reg_addr == KEYMGR_SW_BINDING_REGWEN_OFFSET);
    addr_hit[11] = (reg_addr == KEYMGR_SEALING_SW_BINDING_0_OFFSET);
    addr_hit[12] = (reg_addr == KEYMGR_SEALING_SW_BINDING_1_OFFSET);
    addr_hit[13] = (reg_addr == KEYMGR_SEALING_SW_BINDING_2_OFFSET);
    addr_hit[14] = (reg_addr == KEYMGR_SEALING_SW_BINDING_3_OFFSET);
    addr_hit[15] = (reg_addr == KEYMGR_SEALING_SW_BINDING_4_OFFSET);
    addr_hit[16] = (reg_addr == KEYMGR_SEALING_SW_BINDING_5_OFFSET);
    addr_hit[17] = (reg_addr == KEYMGR_SEALING_SW_BINDING_6_OFFSET);
    addr_hit[18] = (reg_addr == KEYMGR_SEALING_SW_BINDING_7_OFFSET);
    addr_hit[19] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_0_OFFSET);
    addr_hit[20] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_1_OFFSET);
    addr_hit[21] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_2_OFFSET);
    addr_hit[22] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_3_OFFSET);
    addr_hit[23] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_4_OFFSET);
    addr_hit[24] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_5_OFFSET);
    addr_hit[25] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_6_OFFSET);
    addr_hit[26] = (reg_addr == KEYMGR_ATTEST_SW_BINDING_7_OFFSET);
    addr_hit[27] = (reg_addr == KEYMGR_SALT_0_OFFSET);
    addr_hit[28] = (reg_addr == KEYMGR_SALT_1_OFFSET);
    addr_hit[29] = (reg_addr == KEYMGR_SALT_2_OFFSET);
    addr_hit[30] = (reg_addr == KEYMGR_SALT_3_OFFSET);
    addr_hit[31] = (reg_addr == KEYMGR_SALT_4_OFFSET);
    addr_hit[32] = (reg_addr == KEYMGR_SALT_5_OFFSET);
    addr_hit[33] = (reg_addr == KEYMGR_SALT_6_OFFSET);
    addr_hit[34] = (reg_addr == KEYMGR_SALT_7_OFFSET);
    addr_hit[35] = (reg_addr == KEYMGR_KEY_VERSION_OFFSET);
    addr_hit[36] = (reg_addr == KEYMGR_MAX_CREATOR_KEY_VER_REGWEN_OFFSET);
    addr_hit[37] = (reg_addr == KEYMGR_MAX_CREATOR_KEY_VER_SHADOWED_OFFSET);
    addr_hit[38] = (reg_addr == KEYMGR_MAX_OWNER_INT_KEY_VER_REGWEN_OFFSET);
    addr_hit[39] = (reg_addr == KEYMGR_MAX_OWNER_INT_KEY_VER_SHADOWED_OFFSET);
    addr_hit[40] = (reg_addr == KEYMGR_MAX_OWNER_KEY_VER_REGWEN_OFFSET);
    addr_hit[41] = (reg_addr == KEYMGR_MAX_OWNER_KEY_VER_SHADOWED_OFFSET);
    addr_hit[42] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_0_OFFSET);
    addr_hit[43] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_1_OFFSET);
    addr_hit[44] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_2_OFFSET);
    addr_hit[45] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_3_OFFSET);
    addr_hit[46] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_4_OFFSET);
    addr_hit[47] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_5_OFFSET);
    addr_hit[48] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_6_OFFSET);
    addr_hit[49] = (reg_addr == KEYMGR_SW_SHARE0_OUTPUT_7_OFFSET);
    addr_hit[50] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_0_OFFSET);
    addr_hit[51] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_1_OFFSET);
    addr_hit[52] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_2_OFFSET);
    addr_hit[53] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_3_OFFSET);
    addr_hit[54] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_4_OFFSET);
    addr_hit[55] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_5_OFFSET);
    addr_hit[56] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_6_OFFSET);
    addr_hit[57] = (reg_addr == KEYMGR_SW_SHARE1_OUTPUT_7_OFFSET);
    addr_hit[58] = (reg_addr == KEYMGR_WORKING_STATE_OFFSET);
    addr_hit[59] = (reg_addr == KEYMGR_OP_STATUS_OFFSET);
    addr_hit[60] = (reg_addr == KEYMGR_ERR_CODE_OFFSET);
    addr_hit[61] = (reg_addr == KEYMGR_FAULT_STATUS_OFFSET);
    addr_hit[62] = (reg_addr == KEYMGR_DEBUG_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(KEYMGR_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(KEYMGR_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(KEYMGR_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(KEYMGR_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(KEYMGR_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(KEYMGR_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(KEYMGR_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(KEYMGR_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(KEYMGR_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(KEYMGR_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(KEYMGR_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(KEYMGR_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(KEYMGR_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(KEYMGR_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(KEYMGR_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(KEYMGR_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(KEYMGR_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(KEYMGR_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(KEYMGR_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(KEYMGR_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(KEYMGR_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(KEYMGR_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(KEYMGR_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(KEYMGR_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(KEYMGR_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(KEYMGR_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(KEYMGR_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(KEYMGR_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(KEYMGR_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(KEYMGR_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(KEYMGR_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(KEYMGR_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(KEYMGR_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(KEYMGR_PERMIT[33] & ~reg_be))) |
               (addr_hit[34] & (|(KEYMGR_PERMIT[34] & ~reg_be))) |
               (addr_hit[35] & (|(KEYMGR_PERMIT[35] & ~reg_be))) |
               (addr_hit[36] & (|(KEYMGR_PERMIT[36] & ~reg_be))) |
               (addr_hit[37] & (|(KEYMGR_PERMIT[37] & ~reg_be))) |
               (addr_hit[38] & (|(KEYMGR_PERMIT[38] & ~reg_be))) |
               (addr_hit[39] & (|(KEYMGR_PERMIT[39] & ~reg_be))) |
               (addr_hit[40] & (|(KEYMGR_PERMIT[40] & ~reg_be))) |
               (addr_hit[41] & (|(KEYMGR_PERMIT[41] & ~reg_be))) |
               (addr_hit[42] & (|(KEYMGR_PERMIT[42] & ~reg_be))) |
               (addr_hit[43] & (|(KEYMGR_PERMIT[43] & ~reg_be))) |
               (addr_hit[44] & (|(KEYMGR_PERMIT[44] & ~reg_be))) |
               (addr_hit[45] & (|(KEYMGR_PERMIT[45] & ~reg_be))) |
               (addr_hit[46] & (|(KEYMGR_PERMIT[46] & ~reg_be))) |
               (addr_hit[47] & (|(KEYMGR_PERMIT[47] & ~reg_be))) |
               (addr_hit[48] & (|(KEYMGR_PERMIT[48] & ~reg_be))) |
               (addr_hit[49] & (|(KEYMGR_PERMIT[49] & ~reg_be))) |
               (addr_hit[50] & (|(KEYMGR_PERMIT[50] & ~reg_be))) |
               (addr_hit[51] & (|(KEYMGR_PERMIT[51] & ~reg_be))) |
               (addr_hit[52] & (|(KEYMGR_PERMIT[52] & ~reg_be))) |
               (addr_hit[53] & (|(KEYMGR_PERMIT[53] & ~reg_be))) |
               (addr_hit[54] & (|(KEYMGR_PERMIT[54] & ~reg_be))) |
               (addr_hit[55] & (|(KEYMGR_PERMIT[55] & ~reg_be))) |
               (addr_hit[56] & (|(KEYMGR_PERMIT[56] & ~reg_be))) |
               (addr_hit[57] & (|(KEYMGR_PERMIT[57] & ~reg_be))) |
               (addr_hit[58] & (|(KEYMGR_PERMIT[58] & ~reg_be))) |
               (addr_hit[59] & (|(KEYMGR_PERMIT[59] & ~reg_be))) |
               (addr_hit[60] & (|(KEYMGR_PERMIT[60] & ~reg_be))) |
               (addr_hit[61] & (|(KEYMGR_PERMIT[61] & ~reg_be))) |
               (addr_hit[62] & (|(KEYMGR_PERMIT[62] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_wd = reg_wdata[0];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_wd = reg_wdata[0];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_wd = reg_wdata[0];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_recov_operation_err_wd = reg_wdata[0];

  assign alert_test_fatal_fault_err_wd = reg_wdata[1];
  assign cfg_regwen_re = addr_hit[4] & reg_re & !reg_error;
  assign start_we = addr_hit[5] & reg_we & !reg_error;

  assign start_wd = reg_wdata[0];
  assign control_shadowed_re = addr_hit[6] & reg_re & !reg_error;
  assign control_shadowed_we = addr_hit[6] & reg_we & !reg_error;

  assign control_shadowed_operation_wd = reg_wdata[6:4];

  assign control_shadowed_cdi_sel_wd = reg_wdata[7];

  assign control_shadowed_dest_sel_wd = reg_wdata[13:12];
  assign sideload_clear_we = addr_hit[7] & reg_we & !reg_error;

  assign sideload_clear_wd = reg_wdata[2:0];
  assign reseed_interval_regwen_we = addr_hit[8] & reg_we & !reg_error;

  assign reseed_interval_regwen_wd = reg_wdata[0];
  assign reseed_interval_shadowed_re = addr_hit[9] & reg_re & !reg_error;
  assign reseed_interval_shadowed_we = addr_hit[9] & reg_we & !reg_error;

  assign reseed_interval_shadowed_wd = reg_wdata[15:0];
  assign sw_binding_regwen_re = addr_hit[10] & reg_re & !reg_error;
  assign sw_binding_regwen_we = addr_hit[10] & reg_we & !reg_error;

  assign sw_binding_regwen_wd = reg_wdata[0];
  assign sealing_sw_binding_0_we = addr_hit[11] & reg_we & !reg_error;

  assign sealing_sw_binding_0_wd = reg_wdata[31:0];
  assign sealing_sw_binding_1_we = addr_hit[12] & reg_we & !reg_error;

  assign sealing_sw_binding_1_wd = reg_wdata[31:0];
  assign sealing_sw_binding_2_we = addr_hit[13] & reg_we & !reg_error;

  assign sealing_sw_binding_2_wd = reg_wdata[31:0];
  assign sealing_sw_binding_3_we = addr_hit[14] & reg_we & !reg_error;

  assign sealing_sw_binding_3_wd = reg_wdata[31:0];
  assign sealing_sw_binding_4_we = addr_hit[15] & reg_we & !reg_error;

  assign sealing_sw_binding_4_wd = reg_wdata[31:0];
  assign sealing_sw_binding_5_we = addr_hit[16] & reg_we & !reg_error;

  assign sealing_sw_binding_5_wd = reg_wdata[31:0];
  assign sealing_sw_binding_6_we = addr_hit[17] & reg_we & !reg_error;

  assign sealing_sw_binding_6_wd = reg_wdata[31:0];
  assign sealing_sw_binding_7_we = addr_hit[18] & reg_we & !reg_error;

  assign sealing_sw_binding_7_wd = reg_wdata[31:0];
  assign attest_sw_binding_0_we = addr_hit[19] & reg_we & !reg_error;

  assign attest_sw_binding_0_wd = reg_wdata[31:0];
  assign attest_sw_binding_1_we = addr_hit[20] & reg_we & !reg_error;

  assign attest_sw_binding_1_wd = reg_wdata[31:0];
  assign attest_sw_binding_2_we = addr_hit[21] & reg_we & !reg_error;

  assign attest_sw_binding_2_wd = reg_wdata[31:0];
  assign attest_sw_binding_3_we = addr_hit[22] & reg_we & !reg_error;

  assign attest_sw_binding_3_wd = reg_wdata[31:0];
  assign attest_sw_binding_4_we = addr_hit[23] & reg_we & !reg_error;

  assign attest_sw_binding_4_wd = reg_wdata[31:0];
  assign attest_sw_binding_5_we = addr_hit[24] & reg_we & !reg_error;

  assign attest_sw_binding_5_wd = reg_wdata[31:0];
  assign attest_sw_binding_6_we = addr_hit[25] & reg_we & !reg_error;

  assign attest_sw_binding_6_wd = reg_wdata[31:0];
  assign attest_sw_binding_7_we = addr_hit[26] & reg_we & !reg_error;

  assign attest_sw_binding_7_wd = reg_wdata[31:0];
  assign salt_0_we = addr_hit[27] & reg_we & !reg_error;

  assign salt_0_wd = reg_wdata[31:0];
  assign salt_1_we = addr_hit[28] & reg_we & !reg_error;

  assign salt_1_wd = reg_wdata[31:0];
  assign salt_2_we = addr_hit[29] & reg_we & !reg_error;

  assign salt_2_wd = reg_wdata[31:0];
  assign salt_3_we = addr_hit[30] & reg_we & !reg_error;

  assign salt_3_wd = reg_wdata[31:0];
  assign salt_4_we = addr_hit[31] & reg_we & !reg_error;

  assign salt_4_wd = reg_wdata[31:0];
  assign salt_5_we = addr_hit[32] & reg_we & !reg_error;

  assign salt_5_wd = reg_wdata[31:0];
  assign salt_6_we = addr_hit[33] & reg_we & !reg_error;

  assign salt_6_wd = reg_wdata[31:0];
  assign salt_7_we = addr_hit[34] & reg_we & !reg_error;

  assign salt_7_wd = reg_wdata[31:0];
  assign key_version_we = addr_hit[35] & reg_we & !reg_error;

  assign key_version_wd = reg_wdata[31:0];
  assign max_creator_key_ver_regwen_we = addr_hit[36] & reg_we & !reg_error;

  assign max_creator_key_ver_regwen_wd = reg_wdata[0];
  assign max_creator_key_ver_shadowed_re = addr_hit[37] & reg_re & !reg_error;
  assign max_creator_key_ver_shadowed_we = addr_hit[37] & reg_we & !reg_error;

  assign max_creator_key_ver_shadowed_wd = reg_wdata[31:0];
  assign max_owner_int_key_ver_regwen_we = addr_hit[38] & reg_we & !reg_error;

  assign max_owner_int_key_ver_regwen_wd = reg_wdata[0];
  assign max_owner_int_key_ver_shadowed_re = addr_hit[39] & reg_re & !reg_error;
  assign max_owner_int_key_ver_shadowed_we = addr_hit[39] & reg_we & !reg_error;

  assign max_owner_int_key_ver_shadowed_wd = reg_wdata[31:0];
  assign max_owner_key_ver_regwen_we = addr_hit[40] & reg_we & !reg_error;

  assign max_owner_key_ver_regwen_wd = reg_wdata[0];
  assign max_owner_key_ver_shadowed_re = addr_hit[41] & reg_re & !reg_error;
  assign max_owner_key_ver_shadowed_we = addr_hit[41] & reg_we & !reg_error;

  assign max_owner_key_ver_shadowed_wd = reg_wdata[31:0];
  assign sw_share0_output_0_re = addr_hit[42] & reg_re & !reg_error;

  assign sw_share0_output_0_wd = '1;
  assign sw_share0_output_1_re = addr_hit[43] & reg_re & !reg_error;

  assign sw_share0_output_1_wd = '1;
  assign sw_share0_output_2_re = addr_hit[44] & reg_re & !reg_error;

  assign sw_share0_output_2_wd = '1;
  assign sw_share0_output_3_re = addr_hit[45] & reg_re & !reg_error;

  assign sw_share0_output_3_wd = '1;
  assign sw_share0_output_4_re = addr_hit[46] & reg_re & !reg_error;

  assign sw_share0_output_4_wd = '1;
  assign sw_share0_output_5_re = addr_hit[47] & reg_re & !reg_error;

  assign sw_share0_output_5_wd = '1;
  assign sw_share0_output_6_re = addr_hit[48] & reg_re & !reg_error;

  assign sw_share0_output_6_wd = '1;
  assign sw_share0_output_7_re = addr_hit[49] & reg_re & !reg_error;

  assign sw_share0_output_7_wd = '1;
  assign sw_share1_output_0_re = addr_hit[50] & reg_re & !reg_error;

  assign sw_share1_output_0_wd = '1;
  assign sw_share1_output_1_re = addr_hit[51] & reg_re & !reg_error;

  assign sw_share1_output_1_wd = '1;
  assign sw_share1_output_2_re = addr_hit[52] & reg_re & !reg_error;

  assign sw_share1_output_2_wd = '1;
  assign sw_share1_output_3_re = addr_hit[53] & reg_re & !reg_error;

  assign sw_share1_output_3_wd = '1;
  assign sw_share1_output_4_re = addr_hit[54] & reg_re & !reg_error;

  assign sw_share1_output_4_wd = '1;
  assign sw_share1_output_5_re = addr_hit[55] & reg_re & !reg_error;

  assign sw_share1_output_5_wd = '1;
  assign sw_share1_output_6_re = addr_hit[56] & reg_re & !reg_error;

  assign sw_share1_output_6_wd = '1;
  assign sw_share1_output_7_re = addr_hit[57] & reg_re & !reg_error;

  assign sw_share1_output_7_wd = '1;
  assign op_status_we = addr_hit[59] & reg_we & !reg_error;

  assign op_status_wd = reg_wdata[1:0];
  assign err_code_we = addr_hit[60] & reg_we & !reg_error;

  assign err_code_invalid_op_wd = reg_wdata[0];

  assign err_code_invalid_kmac_input_wd = reg_wdata[1];

  assign err_code_invalid_shadow_update_wd = reg_wdata[2];
  assign debug_we = addr_hit[62] & reg_we & !reg_error;

  assign debug_invalid_creator_seed_wd = reg_wdata[0];

  assign debug_invalid_owner_seed_wd = reg_wdata[1];

  assign debug_invalid_dev_id_wd = reg_wdata[2];

  assign debug_invalid_health_state_wd = reg_wdata[3];

  assign debug_invalid_key_version_wd = reg_wdata[4];

  assign debug_invalid_key_wd = reg_wdata[5];

  assign debug_invalid_digest_wd = reg_wdata[6];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = 1'b0;
    reg_we_check[5] = start_gated_we;
    reg_we_check[6] = control_shadowed_gated_we;
    reg_we_check[7] = sideload_clear_gated_we;
    reg_we_check[8] = reseed_interval_regwen_we;
    reg_we_check[9] = reseed_interval_shadowed_gated_we;
    reg_we_check[10] = sw_binding_regwen_we;
    reg_we_check[11] = sealing_sw_binding_0_gated_we;
    reg_we_check[12] = sealing_sw_binding_1_gated_we;
    reg_we_check[13] = sealing_sw_binding_2_gated_we;
    reg_we_check[14] = sealing_sw_binding_3_gated_we;
    reg_we_check[15] = sealing_sw_binding_4_gated_we;
    reg_we_check[16] = sealing_sw_binding_5_gated_we;
    reg_we_check[17] = sealing_sw_binding_6_gated_we;
    reg_we_check[18] = sealing_sw_binding_7_gated_we;
    reg_we_check[19] = attest_sw_binding_0_gated_we;
    reg_we_check[20] = attest_sw_binding_1_gated_we;
    reg_we_check[21] = attest_sw_binding_2_gated_we;
    reg_we_check[22] = attest_sw_binding_3_gated_we;
    reg_we_check[23] = attest_sw_binding_4_gated_we;
    reg_we_check[24] = attest_sw_binding_5_gated_we;
    reg_we_check[25] = attest_sw_binding_6_gated_we;
    reg_we_check[26] = attest_sw_binding_7_gated_we;
    reg_we_check[27] = salt_0_gated_we;
    reg_we_check[28] = salt_1_gated_we;
    reg_we_check[29] = salt_2_gated_we;
    reg_we_check[30] = salt_3_gated_we;
    reg_we_check[31] = salt_4_gated_we;
    reg_we_check[32] = salt_5_gated_we;
    reg_we_check[33] = salt_6_gated_we;
    reg_we_check[34] = salt_7_gated_we;
    reg_we_check[35] = key_version_gated_we;
    reg_we_check[36] = max_creator_key_ver_regwen_we;
    reg_we_check[37] = max_creator_key_ver_shadowed_gated_we;
    reg_we_check[38] = max_owner_int_key_ver_regwen_we;
    reg_we_check[39] = max_owner_int_key_ver_shadowed_gated_we;
    reg_we_check[40] = max_owner_key_ver_regwen_we;
    reg_we_check[41] = max_owner_key_ver_shadowed_gated_we;
    reg_we_check[42] = 1'b0;
    reg_we_check[43] = 1'b0;
    reg_we_check[44] = 1'b0;
    reg_we_check[45] = 1'b0;
    reg_we_check[46] = 1'b0;
    reg_we_check[47] = 1'b0;
    reg_we_check[48] = 1'b0;
    reg_we_check[49] = 1'b0;
    reg_we_check[50] = 1'b0;
    reg_we_check[51] = 1'b0;
    reg_we_check[52] = 1'b0;
    reg_we_check[53] = 1'b0;
    reg_we_check[54] = 1'b0;
    reg_we_check[55] = 1'b0;
    reg_we_check[56] = 1'b0;
    reg_we_check[57] = 1'b0;
    reg_we_check[58] = 1'b0;
    reg_we_check[59] = op_status_we;
    reg_we_check[60] = err_code_we;
    reg_we_check[61] = 1'b0;
    reg_we_check[62] = debug_we;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[0] = cfg_regwen_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[0] = start_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[6:4] = control_shadowed_operation_qs;
        reg_rdata_next[7] = control_shadowed_cdi_sel_qs;
        reg_rdata_next[13:12] = control_shadowed_dest_sel_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[2:0] = sideload_clear_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[0] = reseed_interval_regwen_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[15:0] = reseed_interval_shadowed_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[0] = sw_binding_regwen_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_0_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_1_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_2_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_3_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_4_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_5_qs;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_6_qs;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = sealing_sw_binding_7_qs;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = attest_sw_binding_0_qs;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = attest_sw_binding_1_qs;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = attest_sw_binding_2_qs;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = attest_sw_binding_3_qs;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = attest_sw_binding_4_qs;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = attest_sw_binding_5_qs;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = attest_sw_binding_6_qs;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = attest_sw_binding_7_qs;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = salt_0_qs;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = salt_1_qs;
      end

      addr_hit[29]: begin
        reg_rdata_next[31:0] = salt_2_qs;
      end

      addr_hit[30]: begin
        reg_rdata_next[31:0] = salt_3_qs;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = salt_4_qs;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = salt_5_qs;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = salt_6_qs;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = salt_7_qs;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = key_version_qs;
      end

      addr_hit[36]: begin
        reg_rdata_next[0] = max_creator_key_ver_regwen_qs;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = max_creator_key_ver_shadowed_qs;
      end

      addr_hit[38]: begin
        reg_rdata_next[0] = max_owner_int_key_ver_regwen_qs;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = max_owner_int_key_ver_shadowed_qs;
      end

      addr_hit[40]: begin
        reg_rdata_next[0] = max_owner_key_ver_regwen_qs;
      end

      addr_hit[41]: begin
        reg_rdata_next[31:0] = max_owner_key_ver_shadowed_qs;
      end

      addr_hit[42]: begin
        reg_rdata_next[31:0] = sw_share0_output_0_qs;
      end

      addr_hit[43]: begin
        reg_rdata_next[31:0] = sw_share0_output_1_qs;
      end

      addr_hit[44]: begin
        reg_rdata_next[31:0] = sw_share0_output_2_qs;
      end

      addr_hit[45]: begin
        reg_rdata_next[31:0] = sw_share0_output_3_qs;
      end

      addr_hit[46]: begin
        reg_rdata_next[31:0] = sw_share0_output_4_qs;
      end

      addr_hit[47]: begin
        reg_rdata_next[31:0] = sw_share0_output_5_qs;
      end

      addr_hit[48]: begin
        reg_rdata_next[31:0] = sw_share0_output_6_qs;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = sw_share0_output_7_qs;
      end

      addr_hit[50]: begin
        reg_rdata_next[31:0] = sw_share1_output_0_qs;
      end

      addr_hit[51]: begin
        reg_rdata_next[31:0] = sw_share1_output_1_qs;
      end

      addr_hit[52]: begin
        reg_rdata_next[31:0] = sw_share1_output_2_qs;
      end

      addr_hit[53]: begin
        reg_rdata_next[31:0] = sw_share1_output_3_qs;
      end

      addr_hit[54]: begin
        reg_rdata_next[31:0] = sw_share1_output_4_qs;
      end

      addr_hit[55]: begin
        reg_rdata_next[31:0] = sw_share1_output_5_qs;
      end

      addr_hit[56]: begin
        reg_rdata_next[31:0] = sw_share1_output_6_qs;
      end

      addr_hit[57]: begin
        reg_rdata_next[31:0] = sw_share1_output_7_qs;
      end

      addr_hit[58]: begin
        reg_rdata_next[2:0] = working_state_qs;
      end

      addr_hit[59]: begin
        reg_rdata_next[1:0] = op_status_qs;
      end

      addr_hit[60]: begin
        reg_rdata_next[0] = err_code_invalid_op_qs;
        reg_rdata_next[1] = err_code_invalid_kmac_input_qs;
        reg_rdata_next[2] = err_code_invalid_shadow_update_qs;
      end

      addr_hit[61]: begin
        reg_rdata_next[0] = fault_status_cmd_qs;
        reg_rdata_next[1] = fault_status_kmac_fsm_qs;
        reg_rdata_next[2] = fault_status_kmac_done_qs;
        reg_rdata_next[3] = fault_status_kmac_op_qs;
        reg_rdata_next[4] = fault_status_kmac_out_qs;
        reg_rdata_next[5] = fault_status_regfile_intg_qs;
        reg_rdata_next[6] = fault_status_shadow_qs;
        reg_rdata_next[7] = fault_status_ctrl_fsm_intg_qs;
        reg_rdata_next[8] = fault_status_ctrl_fsm_chk_qs;
        reg_rdata_next[9] = fault_status_ctrl_fsm_cnt_qs;
        reg_rdata_next[10] = fault_status_reseed_cnt_qs;
        reg_rdata_next[11] = fault_status_side_ctrl_fsm_qs;
        reg_rdata_next[12] = fault_status_side_ctrl_sel_qs;
        reg_rdata_next[13] = fault_status_key_ecc_qs;
      end

      addr_hit[62]: begin
        reg_rdata_next[0] = debug_invalid_creator_seed_qs;
        reg_rdata_next[1] = debug_invalid_owner_seed_qs;
        reg_rdata_next[2] = debug_invalid_dev_id_qs;
        reg_rdata_next[3] = debug_invalid_health_state_qs;
        reg_rdata_next[4] = debug_invalid_key_version_qs;
        reg_rdata_next[5] = debug_invalid_key_qs;
        reg_rdata_next[6] = debug_invalid_digest_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  logic rst_done;
  logic shadow_rst_done;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rst_done <= '0;
    end else begin
      rst_done <= 1'b1;
    end
  end

  always_ff @(posedge clk_i or negedge rst_shadowed_ni) begin
    if (!rst_shadowed_ni) begin
      shadow_rst_done <= '0;
    end else begin
      shadow_rst_done <= 1'b1;
    end
  end

  // both shadow and normal resets have been released
  assign shadow_busy = ~(rst_done & shadow_rst_done);

  // Collect up storage and update errors
  assign shadowed_storage_err_o = |{
    control_shadowed_operation_storage_err,
    control_shadowed_cdi_sel_storage_err,
    control_shadowed_dest_sel_storage_err,
    reseed_interval_shadowed_storage_err,
    max_creator_key_ver_shadowed_storage_err,
    max_owner_int_key_ver_shadowed_storage_err,
    max_owner_key_ver_shadowed_storage_err
  };
  assign shadowed_update_err_o = |{
    control_shadowed_operation_update_err,
    control_shadowed_cdi_sel_update_err,
    control_shadowed_dest_sel_update_err,
    reseed_interval_shadowed_update_err,
    max_creator_key_ver_shadowed_update_err,
    max_owner_int_key_ver_shadowed_update_err,
    max_owner_key_ver_shadowed_update_err
  };

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager entropy reseed controls
//

`include "prim_assert.sv"

module keymgr_reseed_ctrl import keymgr_pkg::*; (
  input clk_i,
  input rst_ni,
  input clk_edn_i,
  input rst_edn_ni,

  // interface to keymgr_ctrl
  input reseed_req_i,
  output logic reseed_ack_o,

  // interface to software
  input [15:0] reseed_interval_i,

  // interface to edn
  output edn_pkg::edn_req_t edn_o,
  input edn_pkg::edn_rsp_t edn_i,

  // interface to lfsr
  output logic seed_en_o,
  output logic [LfsrWidth-1:0] seed_o,

  // error condition
  output logic cnt_err_o
);

  logic local_req;
  logic edn_req;
  logic edn_ack;
  logic [15:0] reseed_cnt;
  logic edn_done;

  assign edn_done = edn_req & edn_ack;

  // An edn request can either come from counter or from external
  assign local_req = reseed_cnt >= reseed_interval_i;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      edn_req <= '0;
    end else if (edn_done) begin
      edn_req <= '0;
    end else if (!edn_req && (reseed_req_i || local_req)) begin
      // if edn request is not going, make a new request
      edn_req <= 1'b1;
    end
  end

  assign seed_en_o = edn_ack;
  assign reseed_ack_o = reseed_req_i & edn_ack;

  prim_edn_req #(
    .OutWidth(LfsrWidth)
  ) u_edn_req (
    .clk_i,
    .rst_ni,
    .req_chk_i(1'b1),
    .req_i(edn_req),
    .ack_o(edn_ack),
    .data_o(seed_o),
    .fips_o(),
    .err_o(),
    .clk_edn_i,
    .rst_edn_ni,
    .edn_o,
    .edn_i
  );


  // suppress first reseed count until the first transaction has gone through.
  // This ensures the first entropy fetch is controlled by software timing and
  // there is no chance to accidentally pick-up boot time entropy unless intended by software.
  logic cnt_en;
  always_ff @(posedge clk_i or negedge rst_ni) begin
     if (!rst_ni) begin
       cnt_en <= '0;
     end else if (edn_done) begin
       cnt_en <= 1'b1;
     end
  end

  // whenever reseed count reaches reseed_interval, issue a request and wait for ack
  // SEC_CM: RESEED.CTR.REDUN
  prim_count #(
    .Width(16)
  ) u_reseed_cnt (
    .clk_i,
    .rst_ni,
    .clr_i(edn_done),
    .set_i('0),
    .set_cnt_i('0),
    .incr_en_i(cnt_en),
    .decr_en_i(1'b0),
    .step_i(16'h1),
    .cnt_o(reseed_cnt),
    .cnt_next_o(),
    .err_o(cnt_err_o)
  );

endmodule // keymgr_reseed_ctrl


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Key manager sideload key

`include "prim_assert.sv"

module keymgr_sideload_key import keymgr_pkg::*; #(
  parameter int Width = KeyWidth
) (
  input clk_i,
  input rst_ni,
  input en_i,
  input set_en_i,
  input set_i,
  input clr_i,
  input [Shares-1:0][RandWidth-1:0] entropy_i,
  input [Shares-1:0][Width-1:0] key_i,
  output logic valid_o,
  output logic [Shares-1:0][Width-1:0] key_o
);

  localparam int EntropyCopies = Width / RandWidth;

  logic valid_q;
  logic [Shares-1:0][Width-1:0] key_q;

  assign valid_o = valid_q & en_i;
  assign key_o = key_q;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      valid_q <= 1'b0;
    end else if (!en_i || clr_i) begin
      valid_q <= 1'b0;
    end else if (set_i) begin
      valid_q <= 1'b1;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      key_q <= '0;
    end else if (clr_i) begin
      for (int i = 0; i < Shares; i++) begin
        key_q[i] <= {EntropyCopies{entropy_i[i]}};
      end
    end else if (set_i) begin
      for (int i = 0; i < Shares; i++) begin
        key_q[i] <= set_en_i ? key_i[i] : {EntropyCopies{entropy_i[i]}};
      end
    end
  end

endmodule // keymgr_sideload_key


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Manage all sideload keys

`include "prim_assert.sv"

module keymgr_sideload_key_ctrl import keymgr_pkg::*;(
  input clk_i,
  input rst_ni,
  input init_i,
  input keymgr_sideload_clr_e clr_key_i, // clear key just deletes the key
  input wipe_key_i,  // wipe key deletes and renders sideloads useless until reboot
  input [Shares-1:0][RandWidth-1:0] entropy_i,
  input keymgr_key_dest_e dest_sel_i,
  input prim_mubi_pkg::mubi4_t hw_key_sel_i,
  input data_en_i,
  input data_valid_i,
  input hw_key_req_t key_i,
  input [Shares-1:0][kmac_pkg::AppDigestW-1:0] data_i,
  output logic prng_en_o,
  output hw_key_req_t aes_key_o,
  output hw_key_req_t kmac_key_o,
  output otbn_key_req_t otbn_key_o,
  output logic sideload_sel_err_o,
  output logic fsm_err_o
);

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 5 -m 4 -n 10 \
  //      -s 1700801647 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: --
  //  4: --
  //  5: |||||||||||||||||||| (33.33%)
  //  6: |||||||||| (16.67%)
  //  7: |||||||||||||||||||| (33.33%)
  //  8: |||||||||| (16.67%)
  //  9: --
  // 10: --
  //
  // Minimum Hamming distance: 5
  // Maximum Hamming distance: 8
  // Minimum Hamming weight: 3
  // Maximum Hamming weight: 7
  //
  localparam int StateWidth = 10;
  typedef enum logic [StateWidth-1:0] {
    StSideloadReset = 10'b0011111011,
    StSideloadIdle  = 10'b0101000101,
    StSideloadWipe  = 10'b1110110010,
    StSideloadStop  = 10'b1000001010
  } keymgr_sideload_e;

  keymgr_sideload_e state_q, state_d;

  // This primitive is used to place a size-only constraint on the
  // flops in order to prevent FSM state encoding optimizations.
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, keymgr_sideload_e, StSideloadReset)

  logic keys_en;
  logic [Shares-1:0][KeyWidth-1:0] data_truncated;
  for(genvar i = 0; i < Shares; i++) begin : gen_truncate_data
    assign data_truncated[i] = data_i[i][KeyWidth-1:0];
  end

  // clear all keys when selected by software, or when
  // wipe command is received
  logic clr_all_keys;
  logic [LastIdx-1:0] slot_clr;
  assign clr_all_keys = wipe_key_i |
                        !(clr_key_i inside {SideLoadClrIdle,
                                            SideLoadClrAes,
                                            SideLoadClrKmac,
                                            SideLoadClrOtbn});

  assign slot_clr[AesIdx]  = clr_all_keys | (clr_key_i == SideLoadClrAes);
  assign slot_clr[KmacIdx] = clr_all_keys | (clr_key_i == SideLoadClrKmac);
  assign slot_clr[OtbnIdx] = clr_all_keys | (clr_key_i == SideLoadClrOtbn);

  logic clr;
  assign clr = |slot_clr;

  always_comb begin
    keys_en = 1'b0;
    state_d = state_q;
    fsm_err_o = 1'b0;

    unique case (state_q)
      StSideloadReset: begin
        if (init_i) begin
          state_d = StSideloadIdle;
        end
      end

      // when clear is received, delete the selected key
      // when wipe is received, delete the key and disable sideload until reboot.
      StSideloadIdle: begin
        keys_en = 1'b1;
        if (wipe_key_i) begin
          state_d = StSideloadWipe;
        end
      end

      StSideloadWipe: begin
        keys_en = 1'b0;
        if (!wipe_key_i) begin
          state_d = StSideloadStop;
        end
      end

      // intentional terminal state
      StSideloadStop: begin
        keys_en = 1'b0;
      end

      default: begin
        fsm_err_o = 1'b1;
      end

    endcase // unique case (state_q)
  end

  import prim_mubi_pkg::mubi4_test_true_strict;
  prim_mubi_pkg::mubi4_t [LastIdx-1:0] hw_key_sel;
  prim_mubi4_sync #(
    .NumCopies(int'(LastIdx)),
    .AsyncOn(0) // clock/reset below is only used for SVAs.
  ) u_mubi_buf (
    .clk_i,
    .rst_ni,
    .mubi_i(hw_key_sel_i),
    .mubi_o(hw_key_sel)
  );

  logic [LastIdx-1:0] slot_sel;
  assign slot_sel[AesIdx] = (dest_sel_i == Aes) & mubi4_test_true_strict(hw_key_sel[AesIdx]);
  assign slot_sel[KmacIdx] = (dest_sel_i == Kmac) & mubi4_test_true_strict(hw_key_sel[KmacIdx]);
  assign slot_sel[OtbnIdx] = (dest_sel_i == Otbn) & mubi4_test_true_strict(hw_key_sel[OtbnIdx]);

  keymgr_sideload_key u_aes_key (
    .clk_i,
    .rst_ni,
    .en_i(keys_en),
    .set_en_i(data_en_i),
    .set_i(data_valid_i & slot_sel[AesIdx]),
    .clr_i(slot_clr[AesIdx]),
    .entropy_i(entropy_i),
    .key_i(data_truncated),
    .valid_o(aes_key_o.valid),
    .key_o(aes_key_o.key)
  );

  keymgr_sideload_key #(
    .Width(OtbnKeyWidth)
  ) u_otbn_key (
    .clk_i,
    .rst_ni,
    .en_i(keys_en),
    .set_en_i(data_en_i),
    .set_i(data_valid_i & slot_sel[OtbnIdx]),
    .clr_i(slot_clr[OtbnIdx]),
    .entropy_i(entropy_i),
    .key_i(data_i),
    .valid_o(otbn_key_o.valid),
    .key_o(otbn_key_o.key)
  );

  hw_key_req_t kmac_sideload_key;
  keymgr_sideload_key u_kmac_key (
    .clk_i,
    .rst_ni,
    .en_i(keys_en),
    .set_en_i(data_en_i),
    .set_i(data_valid_i & slot_sel[KmacIdx]),
    .clr_i(slot_clr[KmacIdx]),
    .entropy_i(entropy_i),
    .key_i(data_truncated),
    .valid_o(kmac_sideload_key.valid),
    .key_o(kmac_sideload_key.key)
  );

  logic [LastIdx-1:0] valid_tracking_q;
  for (genvar i = int'(AesIdx); i < LastIdx; i++) begin : gen_tracking_valid
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        valid_tracking_q[i] <= '0;
      end else if (slot_clr[i]) begin
        valid_tracking_q[i] <= '0;
      end else if (slot_sel[i])begin
        valid_tracking_q[i] <= 1'b1;
      end
    end
  end

  // SEC_CM: SIDE_LOAD_SEL.CTRL.CONSISTENCY
  logic [LastIdx-1:0] valids;
  assign valids[AesIdx] = aes_key_o.valid;
  assign valids[KmacIdx] = kmac_sideload_key.valid;
  assign valids[OtbnIdx] = otbn_key_o.valid;

  // If valid tracking claims a valid should be 0 but 1 is observed, it is
  // an error.
  // Note the sideload error is not a direct constant comparision. Instead
  // it provides hint when valids is allowed to be valid.  If valid becomes
  // 1 outside that window, then an error is triggered.
  assign sideload_sel_err_o = |(~valid_tracking_q & valids);

  // when directed by keymgr_ctrl, switch over to internal key and feed to kmac
  assign kmac_key_o = key_i.valid ? key_i : kmac_sideload_key;

  // when clearing, request prng
  assign prng_en_o = clr;


  /////////////////////////////////////
  //  Assertions
  /////////////////////////////////////

  // When updating a sideload key, the secret key state must always be used as the source
  `ASSERT(KmacKeySource_a, data_valid_i |-> key_i.valid)

endmodule // keymgr_sideload_key_ctrl


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package kmac_reg_pkg;

  // Param list
  parameter int NumWordsKey = 16;
  parameter int NumWordsPrefix = 11;
  parameter int NumEntriesMsgFifo = 10;
  parameter int NumBytesMsgFifoEntry = 8;
  parameter int unsigned HashCntW = 10;
  parameter int NumSeedsEntropyLfsr = 5;
  parameter int NumAlerts = 2;

  // Address widths within the block
  parameter int BlockAw = 12;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
    } kmac_done;
    struct packed {
      logic        q;
    } fifo_empty;
    struct packed {
      logic        q;
    } kmac_err;
  } kmac_reg2hw_intr_state_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } kmac_done;
    struct packed {
      logic        q;
    } fifo_empty;
    struct packed {
      logic        q;
    } kmac_err;
  } kmac_reg2hw_intr_enable_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } kmac_done;
    struct packed {
      logic        q;
      logic        qe;
    } fifo_empty;
    struct packed {
      logic        q;
      logic        qe;
    } kmac_err;
  } kmac_reg2hw_intr_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } recov_operation_err;
    struct packed {
      logic        q;
      logic        qe;
    } fatal_fault_err;
  } kmac_reg2hw_alert_test_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } kmac_en;
    struct packed {
      logic [2:0]  q;
      logic        qe;
    } kstrength;
    struct packed {
      logic [1:0]  q;
      logic        qe;
    } mode;
    struct packed {
      logic        q;
      logic        qe;
    } msg_endianness;
    struct packed {
      logic        q;
      logic        qe;
    } state_endianness;
    struct packed {
      logic        q;
      logic        qe;
    } sideload;
    struct packed {
      logic [1:0]  q;
      logic        qe;
    } entropy_mode;
    struct packed {
      logic        q;
      logic        qe;
    } entropy_fast_process;
    struct packed {
      logic        q;
      logic        qe;
    } msg_mask;
    struct packed {
      logic        q;
      logic        qe;
    } entropy_ready;
    struct packed {
      logic        q;
      logic        qe;
    } err_processed;
    struct packed {
      logic        q;
      logic        qe;
    } en_unsupported_modestrength;
  } kmac_reg2hw_cfg_shadowed_reg_t;

  typedef struct packed {
    struct packed {
      logic [5:0]  q;
      logic        qe;
    } cmd;
    struct packed {
      logic        q;
      logic        qe;
    } entropy_req;
    struct packed {
      logic        q;
      logic        qe;
    } hash_cnt_clr;
  } kmac_reg2hw_cmd_reg_t;

  typedef struct packed {
    struct packed {
      logic [9:0] q;
    } prescaler;
    struct packed {
      logic [15:0] q;
    } wait_timer;
  } kmac_reg2hw_entropy_period_reg_t;

  typedef struct packed {
    logic [9:0] q;
  } kmac_reg2hw_entropy_refresh_threshold_shadowed_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } kmac_reg2hw_entropy_seed_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } kmac_reg2hw_key_share0_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } kmac_reg2hw_key_share1_mreg_t;

  typedef struct packed {
    logic [2:0]  q;
  } kmac_reg2hw_key_len_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } kmac_reg2hw_prefix_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } kmac_done;
    struct packed {
      logic        d;
      logic        de;
    } fifo_empty;
    struct packed {
      logic        d;
      logic        de;
    } kmac_err;
  } kmac_hw2reg_intr_state_reg_t;

  typedef struct packed {
    logic        d;
  } kmac_hw2reg_cfg_regwen_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
    } sha3_idle;
    struct packed {
      logic        d;
    } sha3_absorb;
    struct packed {
      logic        d;
    } sha3_squeeze;
    struct packed {
      logic [4:0]  d;
    } fifo_depth;
    struct packed {
      logic        d;
    } fifo_empty;
    struct packed {
      logic        d;
    } fifo_full;
    struct packed {
      logic        d;
    } alert_fatal_fault;
    struct packed {
      logic        d;
    } alert_recov_ctrl_update_err;
  } kmac_hw2reg_status_reg_t;

  typedef struct packed {
    logic [9:0] d;
    logic        de;
  } kmac_hw2reg_entropy_refresh_hash_cnt_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } kmac_hw2reg_err_code_reg_t;

  // Register -> HW type
  typedef struct packed {
    kmac_reg2hw_intr_state_reg_t intr_state; // [1666:1664]
    kmac_reg2hw_intr_enable_reg_t intr_enable; // [1663:1661]
    kmac_reg2hw_intr_test_reg_t intr_test; // [1660:1655]
    kmac_reg2hw_alert_test_reg_t alert_test; // [1654:1651]
    kmac_reg2hw_cfg_shadowed_reg_t cfg_shadowed; // [1650:1623]
    kmac_reg2hw_cmd_reg_t cmd; // [1622:1612]
    kmac_reg2hw_entropy_period_reg_t entropy_period; // [1611:1586]
    kmac_reg2hw_entropy_refresh_threshold_shadowed_reg_t
        entropy_refresh_threshold_shadowed; // [1585:1576]
    kmac_reg2hw_entropy_seed_mreg_t [4:0] entropy_seed; // [1575:1411]
    kmac_reg2hw_key_share0_mreg_t [15:0] key_share0; // [1410:883]
    kmac_reg2hw_key_share1_mreg_t [15:0] key_share1; // [882:355]
    kmac_reg2hw_key_len_reg_t key_len; // [354:352]
    kmac_reg2hw_prefix_mreg_t [10:0] prefix; // [351:0]
  } kmac_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    kmac_hw2reg_intr_state_reg_t intr_state; // [62:57]
    kmac_hw2reg_cfg_regwen_reg_t cfg_regwen; // [56:56]
    kmac_hw2reg_status_reg_t status; // [55:44]
    kmac_hw2reg_entropy_refresh_hash_cnt_reg_t entropy_refresh_hash_cnt; // [43:33]
    kmac_hw2reg_err_code_reg_t err_code; // [32:0]
  } kmac_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] KMAC_INTR_STATE_OFFSET = 12'h 0;
  parameter logic [BlockAw-1:0] KMAC_INTR_ENABLE_OFFSET = 12'h 4;
  parameter logic [BlockAw-1:0] KMAC_INTR_TEST_OFFSET = 12'h 8;
  parameter logic [BlockAw-1:0] KMAC_ALERT_TEST_OFFSET = 12'h c;
  parameter logic [BlockAw-1:0] KMAC_CFG_REGWEN_OFFSET = 12'h 10;
  parameter logic [BlockAw-1:0] KMAC_CFG_SHADOWED_OFFSET = 12'h 14;
  parameter logic [BlockAw-1:0] KMAC_CMD_OFFSET = 12'h 18;
  parameter logic [BlockAw-1:0] KMAC_STATUS_OFFSET = 12'h 1c;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_PERIOD_OFFSET = 12'h 20;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_REFRESH_HASH_CNT_OFFSET = 12'h 24;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_REFRESH_THRESHOLD_SHADOWED_OFFSET = 12'h 28;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_SEED_0_OFFSET = 12'h 2c;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_SEED_1_OFFSET = 12'h 30;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_SEED_2_OFFSET = 12'h 34;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_SEED_3_OFFSET = 12'h 38;
  parameter logic [BlockAw-1:0] KMAC_ENTROPY_SEED_4_OFFSET = 12'h 3c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_0_OFFSET = 12'h 40;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_1_OFFSET = 12'h 44;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_2_OFFSET = 12'h 48;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_3_OFFSET = 12'h 4c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_4_OFFSET = 12'h 50;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_5_OFFSET = 12'h 54;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_6_OFFSET = 12'h 58;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_7_OFFSET = 12'h 5c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_8_OFFSET = 12'h 60;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_9_OFFSET = 12'h 64;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_10_OFFSET = 12'h 68;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_11_OFFSET = 12'h 6c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_12_OFFSET = 12'h 70;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_13_OFFSET = 12'h 74;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_14_OFFSET = 12'h 78;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE0_15_OFFSET = 12'h 7c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_0_OFFSET = 12'h 80;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_1_OFFSET = 12'h 84;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_2_OFFSET = 12'h 88;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_3_OFFSET = 12'h 8c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_4_OFFSET = 12'h 90;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_5_OFFSET = 12'h 94;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_6_OFFSET = 12'h 98;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_7_OFFSET = 12'h 9c;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_8_OFFSET = 12'h a0;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_9_OFFSET = 12'h a4;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_10_OFFSET = 12'h a8;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_11_OFFSET = 12'h ac;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_12_OFFSET = 12'h b0;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_13_OFFSET = 12'h b4;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_14_OFFSET = 12'h b8;
  parameter logic [BlockAw-1:0] KMAC_KEY_SHARE1_15_OFFSET = 12'h bc;
  parameter logic [BlockAw-1:0] KMAC_KEY_LEN_OFFSET = 12'h c0;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_0_OFFSET = 12'h c4;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_1_OFFSET = 12'h c8;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_2_OFFSET = 12'h cc;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_3_OFFSET = 12'h d0;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_4_OFFSET = 12'h d4;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_5_OFFSET = 12'h d8;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_6_OFFSET = 12'h dc;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_7_OFFSET = 12'h e0;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_8_OFFSET = 12'h e4;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_9_OFFSET = 12'h e8;
  parameter logic [BlockAw-1:0] KMAC_PREFIX_10_OFFSET = 12'h ec;
  parameter logic [BlockAw-1:0] KMAC_ERR_CODE_OFFSET = 12'h f0;

  // Reset values for hwext registers and their fields
  parameter logic [2:0] KMAC_INTR_TEST_RESVAL = 3'h 0;
  parameter logic [0:0] KMAC_INTR_TEST_KMAC_DONE_RESVAL = 1'h 0;
  parameter logic [0:0] KMAC_INTR_TEST_FIFO_EMPTY_RESVAL = 1'h 0;
  parameter logic [0:0] KMAC_INTR_TEST_KMAC_ERR_RESVAL = 1'h 0;
  parameter logic [1:0] KMAC_ALERT_TEST_RESVAL = 2'h 0;
  parameter logic [0:0] KMAC_ALERT_TEST_RECOV_OPERATION_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] KMAC_ALERT_TEST_FATAL_FAULT_ERR_RESVAL = 1'h 0;
  parameter logic [0:0] KMAC_CFG_REGWEN_RESVAL = 1'h 1;
  parameter logic [0:0] KMAC_CFG_REGWEN_EN_RESVAL = 1'h 1;
  parameter logic [9:0] KMAC_CMD_RESVAL = 10'h 0;
  parameter logic [17:0] KMAC_STATUS_RESVAL = 18'h 4001;
  parameter logic [0:0] KMAC_STATUS_SHA3_IDLE_RESVAL = 1'h 1;
  parameter logic [0:0] KMAC_STATUS_FIFO_EMPTY_RESVAL = 1'h 1;
  parameter logic [0:0] KMAC_STATUS_ALERT_FATAL_FAULT_RESVAL = 1'h 0;
  parameter logic [0:0] KMAC_STATUS_ALERT_RECOV_CTRL_UPDATE_ERR_RESVAL = 1'h 0;
  parameter logic [31:0] KMAC_ENTROPY_SEED_0_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_ENTROPY_SEED_1_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_ENTROPY_SEED_2_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_ENTROPY_SEED_3_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_ENTROPY_SEED_4_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_0_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_1_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_2_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_3_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_4_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_5_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_6_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_7_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_8_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_9_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_10_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_11_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_12_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_13_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_14_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE0_15_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_0_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_1_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_2_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_3_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_4_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_5_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_6_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_7_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_8_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_9_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_10_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_11_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_12_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_13_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_14_RESVAL = 32'h 0;
  parameter logic [31:0] KMAC_KEY_SHARE1_15_RESVAL = 32'h 0;

  // Window parameters
  parameter logic [BlockAw-1:0] KMAC_STATE_OFFSET = 12'h 400;
  parameter int unsigned        KMAC_STATE_SIZE   = 'h 200;
  parameter logic [BlockAw-1:0] KMAC_MSG_FIFO_OFFSET = 12'h 800;
  parameter int unsigned        KMAC_MSG_FIFO_SIZE   = 'h 800;

  // Register index
  typedef enum int {
    KMAC_INTR_STATE,
    KMAC_INTR_ENABLE,
    KMAC_INTR_TEST,
    KMAC_ALERT_TEST,
    KMAC_CFG_REGWEN,
    KMAC_CFG_SHADOWED,
    KMAC_CMD,
    KMAC_STATUS,
    KMAC_ENTROPY_PERIOD,
    KMAC_ENTROPY_REFRESH_HASH_CNT,
    KMAC_ENTROPY_REFRESH_THRESHOLD_SHADOWED,
    KMAC_ENTROPY_SEED_0,
    KMAC_ENTROPY_SEED_1,
    KMAC_ENTROPY_SEED_2,
    KMAC_ENTROPY_SEED_3,
    KMAC_ENTROPY_SEED_4,
    KMAC_KEY_SHARE0_0,
    KMAC_KEY_SHARE0_1,
    KMAC_KEY_SHARE0_2,
    KMAC_KEY_SHARE0_3,
    KMAC_KEY_SHARE0_4,
    KMAC_KEY_SHARE0_5,
    KMAC_KEY_SHARE0_6,
    KMAC_KEY_SHARE0_7,
    KMAC_KEY_SHARE0_8,
    KMAC_KEY_SHARE0_9,
    KMAC_KEY_SHARE0_10,
    KMAC_KEY_SHARE0_11,
    KMAC_KEY_SHARE0_12,
    KMAC_KEY_SHARE0_13,
    KMAC_KEY_SHARE0_14,
    KMAC_KEY_SHARE0_15,
    KMAC_KEY_SHARE1_0,
    KMAC_KEY_SHARE1_1,
    KMAC_KEY_SHARE1_2,
    KMAC_KEY_SHARE1_3,
    KMAC_KEY_SHARE1_4,
    KMAC_KEY_SHARE1_5,
    KMAC_KEY_SHARE1_6,
    KMAC_KEY_SHARE1_7,
    KMAC_KEY_SHARE1_8,
    KMAC_KEY_SHARE1_9,
    KMAC_KEY_SHARE1_10,
    KMAC_KEY_SHARE1_11,
    KMAC_KEY_SHARE1_12,
    KMAC_KEY_SHARE1_13,
    KMAC_KEY_SHARE1_14,
    KMAC_KEY_SHARE1_15,
    KMAC_KEY_LEN,
    KMAC_PREFIX_0,
    KMAC_PREFIX_1,
    KMAC_PREFIX_2,
    KMAC_PREFIX_3,
    KMAC_PREFIX_4,
    KMAC_PREFIX_5,
    KMAC_PREFIX_6,
    KMAC_PREFIX_7,
    KMAC_PREFIX_8,
    KMAC_PREFIX_9,
    KMAC_PREFIX_10,
    KMAC_ERR_CODE
  } kmac_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] KMAC_PERMIT [61] = '{
    4'b 0001, // index[ 0] KMAC_INTR_STATE
    4'b 0001, // index[ 1] KMAC_INTR_ENABLE
    4'b 0001, // index[ 2] KMAC_INTR_TEST
    4'b 0001, // index[ 3] KMAC_ALERT_TEST
    4'b 0001, // index[ 4] KMAC_CFG_REGWEN
    4'b 1111, // index[ 5] KMAC_CFG_SHADOWED
    4'b 0011, // index[ 6] KMAC_CMD
    4'b 0111, // index[ 7] KMAC_STATUS
    4'b 1111, // index[ 8] KMAC_ENTROPY_PERIOD
    4'b 0011, // index[ 9] KMAC_ENTROPY_REFRESH_HASH_CNT
    4'b 0011, // index[10] KMAC_ENTROPY_REFRESH_THRESHOLD_SHADOWED
    4'b 1111, // index[11] KMAC_ENTROPY_SEED_0
    4'b 1111, // index[12] KMAC_ENTROPY_SEED_1
    4'b 1111, // index[13] KMAC_ENTROPY_SEED_2
    4'b 1111, // index[14] KMAC_ENTROPY_SEED_3
    4'b 1111, // index[15] KMAC_ENTROPY_SEED_4
    4'b 1111, // index[16] KMAC_KEY_SHARE0_0
    4'b 1111, // index[17] KMAC_KEY_SHARE0_1
    4'b 1111, // index[18] KMAC_KEY_SHARE0_2
    4'b 1111, // index[19] KMAC_KEY_SHARE0_3
    4'b 1111, // index[20] KMAC_KEY_SHARE0_4
    4'b 1111, // index[21] KMAC_KEY_SHARE0_5
    4'b 1111, // index[22] KMAC_KEY_SHARE0_6
    4'b 1111, // index[23] KMAC_KEY_SHARE0_7
    4'b 1111, // index[24] KMAC_KEY_SHARE0_8
    4'b 1111, // index[25] KMAC_KEY_SHARE0_9
    4'b 1111, // index[26] KMAC_KEY_SHARE0_10
    4'b 1111, // index[27] KMAC_KEY_SHARE0_11
    4'b 1111, // index[28] KMAC_KEY_SHARE0_12
    4'b 1111, // index[29] KMAC_KEY_SHARE0_13
    4'b 1111, // index[30] KMAC_KEY_SHARE0_14
    4'b 1111, // index[31] KMAC_KEY_SHARE0_15
    4'b 1111, // index[32] KMAC_KEY_SHARE1_0
    4'b 1111, // index[33] KMAC_KEY_SHARE1_1
    4'b 1111, // index[34] KMAC_KEY_SHARE1_2
    4'b 1111, // index[35] KMAC_KEY_SHARE1_3
    4'b 1111, // index[36] KMAC_KEY_SHARE1_4
    4'b 1111, // index[37] KMAC_KEY_SHARE1_5
    4'b 1111, // index[38] KMAC_KEY_SHARE1_6
    4'b 1111, // index[39] KMAC_KEY_SHARE1_7
    4'b 1111, // index[40] KMAC_KEY_SHARE1_8
    4'b 1111, // index[41] KMAC_KEY_SHARE1_9
    4'b 1111, // index[42] KMAC_KEY_SHARE1_10
    4'b 1111, // index[43] KMAC_KEY_SHARE1_11
    4'b 1111, // index[44] KMAC_KEY_SHARE1_12
    4'b 1111, // index[45] KMAC_KEY_SHARE1_13
    4'b 1111, // index[46] KMAC_KEY_SHARE1_14
    4'b 1111, // index[47] KMAC_KEY_SHARE1_15
    4'b 0001, // index[48] KMAC_KEY_LEN
    4'b 1111, // index[49] KMAC_PREFIX_0
    4'b 1111, // index[50] KMAC_PREFIX_1
    4'b 1111, // index[51] KMAC_PREFIX_2
    4'b 1111, // index[52] KMAC_PREFIX_3
    4'b 1111, // index[53] KMAC_PREFIX_4
    4'b 1111, // index[54] KMAC_PREFIX_5
    4'b 1111, // index[55] KMAC_PREFIX_6
    4'b 1111, // index[56] KMAC_PREFIX_7
    4'b 1111, // index[57] KMAC_PREFIX_8
    4'b 1111, // index[58] KMAC_PREFIX_9
    4'b 1111, // index[59] KMAC_PREFIX_10
    4'b 1111  // index[60] KMAC_ERR_CODE
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module kmac_reg_top (
  input clk_i,
  input rst_ni,
  input rst_shadowed_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // Output port for window
  output tlul_pkg::tl_h2d_t tl_win_o  [2],
  input  tlul_pkg::tl_d2h_t tl_win_i  [2],

  // To HW
  output kmac_reg_pkg::kmac_reg2hw_t reg2hw, // Write
  input  kmac_reg_pkg::kmac_hw2reg_t hw2reg, // Read

  output logic shadowed_storage_err_o,
  output logic shadowed_update_err_o,

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import kmac_reg_pkg::* ;

  localparam int AW = 12;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [60:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(61)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  tlul_pkg::tl_h2d_t tl_socket_h2d [3];
  tlul_pkg::tl_d2h_t tl_socket_d2h [3];

  logic [1:0] reg_steer;

  // socket_1n connection
  assign tl_reg_h2d = tl_socket_h2d[2];
  assign tl_socket_d2h[2] = tl_reg_d2h;

  assign tl_win_o[0] = tl_socket_h2d[0];
  assign tl_socket_d2h[0] = tl_win_i[0];
  assign tl_win_o[1] = tl_socket_h2d[1];
  assign tl_socket_d2h[1] = tl_win_i[1];

  // Create Socket_1n
  tlul_socket_1n #(
    .N            (3),
    .HReqPass     (1'b1),
    .HRspPass     (1'b1),
    .DReqPass     ({3{1'b1}}),
    .DRspPass     ({3{1'b1}}),
    .HReqDepth    (4'h0),
    .HRspDepth    (4'h0),
    .DReqDepth    ({3{4'h0}}),
    .DRspDepth    ({3{4'h0}}),
    .ExplicitErrs (1'b0)
  ) u_socket (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),
    .tl_h_i (tl_i),
    .tl_h_o (tl_o_pre),
    .tl_d_o (tl_socket_h2d),
    .tl_d_i (tl_socket_d2h),
    .dev_select_i (reg_steer)
  );

  // Create steering logic
  always_comb begin
    reg_steer =
        tl_i.a_address[AW-1:0] inside {[1024:1535]} ? 2'd0 :
        tl_i.a_address[AW-1:0] inside {[2048:4095]} ? 2'd1 :
        // Default set to register
        2'd2;

    // Override this in case of an integrity error
    if (intg_err) begin
      reg_steer = 2'd2;
    end
  end

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic intr_state_we;
  logic intr_state_kmac_done_qs;
  logic intr_state_kmac_done_wd;
  logic intr_state_fifo_empty_qs;
  logic intr_state_fifo_empty_wd;
  logic intr_state_kmac_err_qs;
  logic intr_state_kmac_err_wd;
  logic intr_enable_we;
  logic intr_enable_kmac_done_qs;
  logic intr_enable_kmac_done_wd;
  logic intr_enable_fifo_empty_qs;
  logic intr_enable_fifo_empty_wd;
  logic intr_enable_kmac_err_qs;
  logic intr_enable_kmac_err_wd;
  logic intr_test_we;
  logic intr_test_kmac_done_wd;
  logic intr_test_fifo_empty_wd;
  logic intr_test_kmac_err_wd;
  logic alert_test_we;
  logic alert_test_recov_operation_err_wd;
  logic alert_test_fatal_fault_err_wd;
  logic cfg_regwen_re;
  logic cfg_regwen_qs;
  logic cfg_shadowed_re;
  logic cfg_shadowed_we;
  logic cfg_shadowed_kmac_en_qs;
  logic cfg_shadowed_kmac_en_wd;
  logic cfg_shadowed_kmac_en_storage_err;
  logic cfg_shadowed_kmac_en_update_err;
  logic [2:0] cfg_shadowed_kstrength_qs;
  logic [2:0] cfg_shadowed_kstrength_wd;
  logic cfg_shadowed_kstrength_storage_err;
  logic cfg_shadowed_kstrength_update_err;
  logic [1:0] cfg_shadowed_mode_qs;
  logic [1:0] cfg_shadowed_mode_wd;
  logic cfg_shadowed_mode_storage_err;
  logic cfg_shadowed_mode_update_err;
  logic cfg_shadowed_msg_endianness_qs;
  logic cfg_shadowed_msg_endianness_wd;
  logic cfg_shadowed_msg_endianness_storage_err;
  logic cfg_shadowed_msg_endianness_update_err;
  logic cfg_shadowed_state_endianness_qs;
  logic cfg_shadowed_state_endianness_wd;
  logic cfg_shadowed_state_endianness_storage_err;
  logic cfg_shadowed_state_endianness_update_err;
  logic cfg_shadowed_sideload_qs;
  logic cfg_shadowed_sideload_wd;
  logic cfg_shadowed_sideload_storage_err;
  logic cfg_shadowed_sideload_update_err;
  logic [1:0] cfg_shadowed_entropy_mode_qs;
  logic [1:0] cfg_shadowed_entropy_mode_wd;
  logic cfg_shadowed_entropy_mode_storage_err;
  logic cfg_shadowed_entropy_mode_update_err;
  logic cfg_shadowed_entropy_fast_process_qs;
  logic cfg_shadowed_entropy_fast_process_wd;
  logic cfg_shadowed_entropy_fast_process_storage_err;
  logic cfg_shadowed_entropy_fast_process_update_err;
  logic cfg_shadowed_msg_mask_qs;
  logic cfg_shadowed_msg_mask_wd;
  logic cfg_shadowed_msg_mask_storage_err;
  logic cfg_shadowed_msg_mask_update_err;
  logic cfg_shadowed_entropy_ready_qs;
  logic cfg_shadowed_entropy_ready_wd;
  logic cfg_shadowed_entropy_ready_storage_err;
  logic cfg_shadowed_entropy_ready_update_err;
  logic cfg_shadowed_err_processed_qs;
  logic cfg_shadowed_err_processed_wd;
  logic cfg_shadowed_err_processed_storage_err;
  logic cfg_shadowed_err_processed_update_err;
  logic cfg_shadowed_en_unsupported_modestrength_qs;
  logic cfg_shadowed_en_unsupported_modestrength_wd;
  logic cfg_shadowed_en_unsupported_modestrength_storage_err;
  logic cfg_shadowed_en_unsupported_modestrength_update_err;
  logic cmd_we;
  logic [5:0] cmd_cmd_wd;
  logic cmd_entropy_req_wd;
  logic cmd_hash_cnt_clr_wd;
  logic status_re;
  logic status_sha3_idle_qs;
  logic status_sha3_absorb_qs;
  logic status_sha3_squeeze_qs;
  logic [4:0] status_fifo_depth_qs;
  logic status_fifo_empty_qs;
  logic status_fifo_full_qs;
  logic status_alert_fatal_fault_qs;
  logic status_alert_recov_ctrl_update_err_qs;
  logic entropy_period_we;
  logic [9:0] entropy_period_prescaler_qs;
  logic [9:0] entropy_period_prescaler_wd;
  logic [15:0] entropy_period_wait_timer_qs;
  logic [15:0] entropy_period_wait_timer_wd;
  logic [9:0] entropy_refresh_hash_cnt_qs;
  logic entropy_refresh_threshold_shadowed_re;
  logic entropy_refresh_threshold_shadowed_we;
  logic [9:0] entropy_refresh_threshold_shadowed_qs;
  logic [9:0] entropy_refresh_threshold_shadowed_wd;
  logic entropy_refresh_threshold_shadowed_storage_err;
  logic entropy_refresh_threshold_shadowed_update_err;
  logic entropy_seed_0_we;
  logic [31:0] entropy_seed_0_wd;
  logic entropy_seed_1_we;
  logic [31:0] entropy_seed_1_wd;
  logic entropy_seed_2_we;
  logic [31:0] entropy_seed_2_wd;
  logic entropy_seed_3_we;
  logic [31:0] entropy_seed_3_wd;
  logic entropy_seed_4_we;
  logic [31:0] entropy_seed_4_wd;
  logic key_share0_0_we;
  logic [31:0] key_share0_0_wd;
  logic key_share0_1_we;
  logic [31:0] key_share0_1_wd;
  logic key_share0_2_we;
  logic [31:0] key_share0_2_wd;
  logic key_share0_3_we;
  logic [31:0] key_share0_3_wd;
  logic key_share0_4_we;
  logic [31:0] key_share0_4_wd;
  logic key_share0_5_we;
  logic [31:0] key_share0_5_wd;
  logic key_share0_6_we;
  logic [31:0] key_share0_6_wd;
  logic key_share0_7_we;
  logic [31:0] key_share0_7_wd;
  logic key_share0_8_we;
  logic [31:0] key_share0_8_wd;
  logic key_share0_9_we;
  logic [31:0] key_share0_9_wd;
  logic key_share0_10_we;
  logic [31:0] key_share0_10_wd;
  logic key_share0_11_we;
  logic [31:0] key_share0_11_wd;
  logic key_share0_12_we;
  logic [31:0] key_share0_12_wd;
  logic key_share0_13_we;
  logic [31:0] key_share0_13_wd;
  logic key_share0_14_we;
  logic [31:0] key_share0_14_wd;
  logic key_share0_15_we;
  logic [31:0] key_share0_15_wd;
  logic key_share1_0_we;
  logic [31:0] key_share1_0_wd;
  logic key_share1_1_we;
  logic [31:0] key_share1_1_wd;
  logic key_share1_2_we;
  logic [31:0] key_share1_2_wd;
  logic key_share1_3_we;
  logic [31:0] key_share1_3_wd;
  logic key_share1_4_we;
  logic [31:0] key_share1_4_wd;
  logic key_share1_5_we;
  logic [31:0] key_share1_5_wd;
  logic key_share1_6_we;
  logic [31:0] key_share1_6_wd;
  logic key_share1_7_we;
  logic [31:0] key_share1_7_wd;
  logic key_share1_8_we;
  logic [31:0] key_share1_8_wd;
  logic key_share1_9_we;
  logic [31:0] key_share1_9_wd;
  logic key_share1_10_we;
  logic [31:0] key_share1_10_wd;
  logic key_share1_11_we;
  logic [31:0] key_share1_11_wd;
  logic key_share1_12_we;
  logic [31:0] key_share1_12_wd;
  logic key_share1_13_we;
  logic [31:0] key_share1_13_wd;
  logic key_share1_14_we;
  logic [31:0] key_share1_14_wd;
  logic key_share1_15_we;
  logic [31:0] key_share1_15_wd;
  logic key_len_we;
  logic [2:0] key_len_wd;
  logic prefix_0_we;
  logic [31:0] prefix_0_qs;
  logic [31:0] prefix_0_wd;
  logic prefix_1_we;
  logic [31:0] prefix_1_qs;
  logic [31:0] prefix_1_wd;
  logic prefix_2_we;
  logic [31:0] prefix_2_qs;
  logic [31:0] prefix_2_wd;
  logic prefix_3_we;
  logic [31:0] prefix_3_qs;
  logic [31:0] prefix_3_wd;
  logic prefix_4_we;
  logic [31:0] prefix_4_qs;
  logic [31:0] prefix_4_wd;
  logic prefix_5_we;
  logic [31:0] prefix_5_qs;
  logic [31:0] prefix_5_wd;
  logic prefix_6_we;
  logic [31:0] prefix_6_qs;
  logic [31:0] prefix_6_wd;
  logic prefix_7_we;
  logic [31:0] prefix_7_qs;
  logic [31:0] prefix_7_wd;
  logic prefix_8_we;
  logic [31:0] prefix_8_qs;
  logic [31:0] prefix_8_wd;
  logic prefix_9_we;
  logic [31:0] prefix_9_qs;
  logic [31:0] prefix_9_wd;
  logic prefix_10_we;
  logic [31:0] prefix_10_qs;
  logic [31:0] prefix_10_wd;
  logic [31:0] err_code_qs;

  // Register instances
  // R[intr_state]: V(False)
  //   F[kmac_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_kmac_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_kmac_done_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.kmac_done.de),
    .d      (hw2reg.intr_state.kmac_done.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.kmac_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_kmac_done_qs)
  );

  //   F[fifo_empty]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_fifo_empty (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_fifo_empty_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.fifo_empty.de),
    .d      (hw2reg.intr_state.fifo_empty.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.fifo_empty.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_fifo_empty_qs)
  );

  //   F[kmac_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessW1C),
    .RESVAL  (1'h0)
  ) u_intr_state_kmac_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_state_we),
    .wd     (intr_state_kmac_err_wd),

    // from internal hardware
    .de     (hw2reg.intr_state.kmac_err.de),
    .d      (hw2reg.intr_state.kmac_err.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_state.kmac_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_state_kmac_err_qs)
  );


  // R[intr_enable]: V(False)
  //   F[kmac_done]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_kmac_done (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_kmac_done_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.kmac_done.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_kmac_done_qs)
  );

  //   F[fifo_empty]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_fifo_empty (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_fifo_empty_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.fifo_empty.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_fifo_empty_qs)
  );

  //   F[kmac_err]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_intr_enable_kmac_err (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (intr_enable_we),
    .wd     (intr_enable_kmac_err_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.intr_enable.kmac_err.q),
    .ds     (),

    // to register interface (read)
    .qs     (intr_enable_kmac_err_qs)
  );


  // R[intr_test]: V(True)
  logic intr_test_qe;
  logic [2:0] intr_test_flds_we;
  assign intr_test_qe = &intr_test_flds_we;
  //   F[kmac_done]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_kmac_done (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_kmac_done_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[0]),
    .q      (reg2hw.intr_test.kmac_done.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.kmac_done.qe = intr_test_qe;

  //   F[fifo_empty]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_fifo_empty (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_fifo_empty_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[1]),
    .q      (reg2hw.intr_test.fifo_empty.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.fifo_empty.qe = intr_test_qe;

  //   F[kmac_err]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_intr_test_kmac_err (
    .re     (1'b0),
    .we     (intr_test_we),
    .wd     (intr_test_kmac_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (intr_test_flds_we[2]),
    .q      (reg2hw.intr_test.kmac_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.intr_test.kmac_err.qe = intr_test_qe;


  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [1:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  //   F[recov_operation_err]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_recov_operation_err (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_recov_operation_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.recov_operation_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.recov_operation_err.qe = alert_test_qe;

  //   F[fatal_fault_err]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test_fatal_fault_err (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_fatal_fault_err_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[1]),
    .q      (reg2hw.alert_test.fatal_fault_err.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.fatal_fault_err.qe = alert_test_qe;


  // R[cfg_regwen]: V(True)
  prim_subreg_ext #(
    .DW    (1)
  ) u_cfg_regwen (
    .re     (cfg_regwen_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.cfg_regwen.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (cfg_regwen_qs)
  );


  // R[cfg_shadowed]: V(False)
  logic cfg_shadowed_qe;
  logic [11:0] cfg_shadowed_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_cfg_shadowed0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&cfg_shadowed_flds_we),
    .q_o(cfg_shadowed_qe)
  );
  // Create REGWEN-gated WE signal
  logic cfg_shadowed_gated_we;
  assign cfg_shadowed_gated_we = cfg_shadowed_we & cfg_regwen_qs;
  //   F[kmac_en]: 0:0
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_kmac_en (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_kmac_en_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[0]),
    .q      (reg2hw.cfg_shadowed.kmac_en.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_kmac_en_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_kmac_en_update_err),
    .err_storage (cfg_shadowed_kmac_en_storage_err)
  );
  assign reg2hw.cfg_shadowed.kmac_en.qe = cfg_shadowed_qe;

  //   F[kstrength]: 3:1
  prim_subreg_shadow #(
    .DW      (3),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (3'h0)
  ) u_cfg_shadowed_kstrength (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_kstrength_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[1]),
    .q      (reg2hw.cfg_shadowed.kstrength.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_kstrength_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_kstrength_update_err),
    .err_storage (cfg_shadowed_kstrength_storage_err)
  );
  assign reg2hw.cfg_shadowed.kstrength.qe = cfg_shadowed_qe;

  //   F[mode]: 5:4
  prim_subreg_shadow #(
    .DW      (2),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (2'h0)
  ) u_cfg_shadowed_mode (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_mode_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[2]),
    .q      (reg2hw.cfg_shadowed.mode.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_mode_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_mode_update_err),
    .err_storage (cfg_shadowed_mode_storage_err)
  );
  assign reg2hw.cfg_shadowed.mode.qe = cfg_shadowed_qe;

  //   F[msg_endianness]: 8:8
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_msg_endianness (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_msg_endianness_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[3]),
    .q      (reg2hw.cfg_shadowed.msg_endianness.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_msg_endianness_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_msg_endianness_update_err),
    .err_storage (cfg_shadowed_msg_endianness_storage_err)
  );
  assign reg2hw.cfg_shadowed.msg_endianness.qe = cfg_shadowed_qe;

  //   F[state_endianness]: 9:9
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_state_endianness (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_state_endianness_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[4]),
    .q      (reg2hw.cfg_shadowed.state_endianness.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_state_endianness_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_state_endianness_update_err),
    .err_storage (cfg_shadowed_state_endianness_storage_err)
  );
  assign reg2hw.cfg_shadowed.state_endianness.qe = cfg_shadowed_qe;

  //   F[sideload]: 12:12
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_sideload (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_sideload_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[5]),
    .q      (reg2hw.cfg_shadowed.sideload.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_sideload_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_sideload_update_err),
    .err_storage (cfg_shadowed_sideload_storage_err)
  );
  assign reg2hw.cfg_shadowed.sideload.qe = cfg_shadowed_qe;

  //   F[entropy_mode]: 17:16
  prim_subreg_shadow #(
    .DW      (2),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (2'h0)
  ) u_cfg_shadowed_entropy_mode (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_entropy_mode_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[6]),
    .q      (reg2hw.cfg_shadowed.entropy_mode.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_entropy_mode_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_entropy_mode_update_err),
    .err_storage (cfg_shadowed_entropy_mode_storage_err)
  );
  assign reg2hw.cfg_shadowed.entropy_mode.qe = cfg_shadowed_qe;

  //   F[entropy_fast_process]: 19:19
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_entropy_fast_process (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_entropy_fast_process_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[7]),
    .q      (reg2hw.cfg_shadowed.entropy_fast_process.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_entropy_fast_process_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_entropy_fast_process_update_err),
    .err_storage (cfg_shadowed_entropy_fast_process_storage_err)
  );
  assign reg2hw.cfg_shadowed.entropy_fast_process.qe = cfg_shadowed_qe;

  //   F[msg_mask]: 20:20
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_msg_mask (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_msg_mask_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[8]),
    .q      (reg2hw.cfg_shadowed.msg_mask.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_msg_mask_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_msg_mask_update_err),
    .err_storage (cfg_shadowed_msg_mask_storage_err)
  );
  assign reg2hw.cfg_shadowed.msg_mask.qe = cfg_shadowed_qe;

  //   F[entropy_ready]: 24:24
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_entropy_ready (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_entropy_ready_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[9]),
    .q      (reg2hw.cfg_shadowed.entropy_ready.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_entropy_ready_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_entropy_ready_update_err),
    .err_storage (cfg_shadowed_entropy_ready_storage_err)
  );
  assign reg2hw.cfg_shadowed.entropy_ready.qe = cfg_shadowed_qe;

  //   F[err_processed]: 25:25
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_err_processed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_err_processed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[10]),
    .q      (reg2hw.cfg_shadowed.err_processed.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_err_processed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_err_processed_update_err),
    .err_storage (cfg_shadowed_err_processed_storage_err)
  );
  assign reg2hw.cfg_shadowed.err_processed.qe = cfg_shadowed_qe;

  //   F[en_unsupported_modestrength]: 26:26
  prim_subreg_shadow #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_cfg_shadowed_en_unsupported_modestrength (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (cfg_shadowed_re),
    .we     (cfg_shadowed_gated_we),
    .wd     (cfg_shadowed_en_unsupported_modestrength_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (cfg_shadowed_flds_we[11]),
    .q      (reg2hw.cfg_shadowed.en_unsupported_modestrength.q),
    .ds     (),

    // to register interface (read)
    .qs     (cfg_shadowed_en_unsupported_modestrength_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (cfg_shadowed_en_unsupported_modestrength_update_err),
    .err_storage (cfg_shadowed_en_unsupported_modestrength_storage_err)
  );
  assign reg2hw.cfg_shadowed.en_unsupported_modestrength.qe = cfg_shadowed_qe;


  // R[cmd]: V(True)
  logic cmd_qe;
  logic [2:0] cmd_flds_we;
  assign cmd_qe = &cmd_flds_we;
  //   F[cmd]: 5:0
  prim_subreg_ext #(
    .DW    (6)
  ) u_cmd_cmd (
    .re     (1'b0),
    .we     (cmd_we),
    .wd     (cmd_cmd_wd),
    .d      ('0),
    .qre    (),
    .qe     (cmd_flds_we[0]),
    .q      (reg2hw.cmd.cmd.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.cmd.cmd.qe = cmd_qe;

  //   F[entropy_req]: 8:8
  prim_subreg_ext #(
    .DW    (1)
  ) u_cmd_entropy_req (
    .re     (1'b0),
    .we     (cmd_we),
    .wd     (cmd_entropy_req_wd),
    .d      ('0),
    .qre    (),
    .qe     (cmd_flds_we[1]),
    .q      (reg2hw.cmd.entropy_req.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.cmd.entropy_req.qe = cmd_qe;

  //   F[hash_cnt_clr]: 9:9
  prim_subreg_ext #(
    .DW    (1)
  ) u_cmd_hash_cnt_clr (
    .re     (1'b0),
    .we     (cmd_we),
    .wd     (cmd_hash_cnt_clr_wd),
    .d      ('0),
    .qre    (),
    .qe     (cmd_flds_we[2]),
    .q      (reg2hw.cmd.hash_cnt_clr.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.cmd.hash_cnt_clr.qe = cmd_qe;


  // R[status]: V(True)
  //   F[sha3_idle]: 0:0
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_sha3_idle (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.sha3_idle.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_sha3_idle_qs)
  );

  //   F[sha3_absorb]: 1:1
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_sha3_absorb (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.sha3_absorb.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_sha3_absorb_qs)
  );

  //   F[sha3_squeeze]: 2:2
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_sha3_squeeze (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.sha3_squeeze.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_sha3_squeeze_qs)
  );

  //   F[fifo_depth]: 12:8
  prim_subreg_ext #(
    .DW    (5)
  ) u_status_fifo_depth (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.fifo_depth.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_fifo_depth_qs)
  );

  //   F[fifo_empty]: 14:14
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_fifo_empty (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.fifo_empty.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_fifo_empty_qs)
  );

  //   F[fifo_full]: 15:15
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_fifo_full (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.fifo_full.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_fifo_full_qs)
  );

  //   F[alert_fatal_fault]: 16:16
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_alert_fatal_fault (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.alert_fatal_fault.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_alert_fatal_fault_qs)
  );

  //   F[alert_recov_ctrl_update_err]: 17:17
  prim_subreg_ext #(
    .DW    (1)
  ) u_status_alert_recov_ctrl_update_err (
    .re     (status_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.status.alert_recov_ctrl_update_err.d),
    .qre    (),
    .qe     (),
    .q      (),
    .ds     (),
    .qs     (status_alert_recov_ctrl_update_err_qs)
  );


  // R[entropy_period]: V(False)
  // Create REGWEN-gated WE signal
  logic entropy_period_gated_we;
  assign entropy_period_gated_we = entropy_period_we & cfg_regwen_qs;
  //   F[prescaler]: 9:0
  prim_subreg #(
    .DW      (10),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (10'h0)
  ) u_entropy_period_prescaler (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (entropy_period_gated_we),
    .wd     (entropy_period_prescaler_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.entropy_period.prescaler.q),
    .ds     (),

    // to register interface (read)
    .qs     (entropy_period_prescaler_qs)
  );

  //   F[wait_timer]: 31:16
  prim_subreg #(
    .DW      (16),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (16'h0)
  ) u_entropy_period_wait_timer (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (entropy_period_gated_we),
    .wd     (entropy_period_wait_timer_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.entropy_period.wait_timer.q),
    .ds     (),

    // to register interface (read)
    .qs     (entropy_period_wait_timer_qs)
  );


  // R[entropy_refresh_hash_cnt]: V(False)
  prim_subreg #(
    .DW      (10),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (10'h0)
  ) u_entropy_refresh_hash_cnt (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.entropy_refresh_hash_cnt.de),
    .d      (hw2reg.entropy_refresh_hash_cnt.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (entropy_refresh_hash_cnt_qs)
  );


  // R[entropy_refresh_threshold_shadowed]: V(False)
  // Create REGWEN-gated WE signal
  logic entropy_refresh_threshold_shadowed_gated_we;
  assign entropy_refresh_threshold_shadowed_gated_we =
    entropy_refresh_threshold_shadowed_we & cfg_regwen_qs;
  prim_subreg_shadow #(
    .DW      (10),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (10'h0)
  ) u_entropy_refresh_threshold_shadowed (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .rst_shadowed_ni (rst_shadowed_ni),

    // from register interface
    .re     (entropy_refresh_threshold_shadowed_re),
    .we     (entropy_refresh_threshold_shadowed_gated_we),
    .wd     (entropy_refresh_threshold_shadowed_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.entropy_refresh_threshold_shadowed.q),
    .ds     (),

    // to register interface (read)
    .qs     (entropy_refresh_threshold_shadowed_qs),

    // Shadow register phase. Relevant for hwext only.
    .phase  (),

    // Shadow register error conditions
    .err_update  (entropy_refresh_threshold_shadowed_update_err),
    .err_storage (entropy_refresh_threshold_shadowed_storage_err)
  );


  // Subregister 0 of Multireg entropy_seed
  // R[entropy_seed_0]: V(True)
  logic entropy_seed_0_qe;
  logic [0:0] entropy_seed_0_flds_we;
  assign entropy_seed_0_qe = &entropy_seed_0_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_entropy_seed_0 (
    .re     (1'b0),
    .we     (entropy_seed_0_we),
    .wd     (entropy_seed_0_wd),
    .d      ('0),
    .qre    (),
    .qe     (entropy_seed_0_flds_we[0]),
    .q      (reg2hw.entropy_seed[0].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.entropy_seed[0].qe = entropy_seed_0_qe;


  // Subregister 1 of Multireg entropy_seed
  // R[entropy_seed_1]: V(True)
  logic entropy_seed_1_qe;
  logic [0:0] entropy_seed_1_flds_we;
  assign entropy_seed_1_qe = &entropy_seed_1_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_entropy_seed_1 (
    .re     (1'b0),
    .we     (entropy_seed_1_we),
    .wd     (entropy_seed_1_wd),
    .d      ('0),
    .qre    (),
    .qe     (entropy_seed_1_flds_we[0]),
    .q      (reg2hw.entropy_seed[1].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.entropy_seed[1].qe = entropy_seed_1_qe;


  // Subregister 2 of Multireg entropy_seed
  // R[entropy_seed_2]: V(True)
  logic entropy_seed_2_qe;
  logic [0:0] entropy_seed_2_flds_we;
  assign entropy_seed_2_qe = &entropy_seed_2_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_entropy_seed_2 (
    .re     (1'b0),
    .we     (entropy_seed_2_we),
    .wd     (entropy_seed_2_wd),
    .d      ('0),
    .qre    (),
    .qe     (entropy_seed_2_flds_we[0]),
    .q      (reg2hw.entropy_seed[2].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.entropy_seed[2].qe = entropy_seed_2_qe;


  // Subregister 3 of Multireg entropy_seed
  // R[entropy_seed_3]: V(True)
  logic entropy_seed_3_qe;
  logic [0:0] entropy_seed_3_flds_we;
  assign entropy_seed_3_qe = &entropy_seed_3_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_entropy_seed_3 (
    .re     (1'b0),
    .we     (entropy_seed_3_we),
    .wd     (entropy_seed_3_wd),
    .d      ('0),
    .qre    (),
    .qe     (entropy_seed_3_flds_we[0]),
    .q      (reg2hw.entropy_seed[3].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.entropy_seed[3].qe = entropy_seed_3_qe;


  // Subregister 4 of Multireg entropy_seed
  // R[entropy_seed_4]: V(True)
  logic entropy_seed_4_qe;
  logic [0:0] entropy_seed_4_flds_we;
  assign entropy_seed_4_qe = &entropy_seed_4_flds_we;
  prim_subreg_ext #(
    .DW    (32)
  ) u_entropy_seed_4 (
    .re     (1'b0),
    .we     (entropy_seed_4_we),
    .wd     (entropy_seed_4_wd),
    .d      ('0),
    .qre    (),
    .qe     (entropy_seed_4_flds_we[0]),
    .q      (reg2hw.entropy_seed[4].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.entropy_seed[4].qe = entropy_seed_4_qe;


  // Subregister 0 of Multireg key_share0
  // R[key_share0_0]: V(True)
  logic key_share0_0_qe;
  logic [0:0] key_share0_0_flds_we;
  assign key_share0_0_qe = &key_share0_0_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_0_gated_we;
  assign key_share0_0_gated_we = key_share0_0_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_0 (
    .re     (1'b0),
    .we     (key_share0_0_gated_we),
    .wd     (key_share0_0_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_0_flds_we[0]),
    .q      (reg2hw.key_share0[0].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[0].qe = key_share0_0_qe;


  // Subregister 1 of Multireg key_share0
  // R[key_share0_1]: V(True)
  logic key_share0_1_qe;
  logic [0:0] key_share0_1_flds_we;
  assign key_share0_1_qe = &key_share0_1_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_1_gated_we;
  assign key_share0_1_gated_we = key_share0_1_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_1 (
    .re     (1'b0),
    .we     (key_share0_1_gated_we),
    .wd     (key_share0_1_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_1_flds_we[0]),
    .q      (reg2hw.key_share0[1].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[1].qe = key_share0_1_qe;


  // Subregister 2 of Multireg key_share0
  // R[key_share0_2]: V(True)
  logic key_share0_2_qe;
  logic [0:0] key_share0_2_flds_we;
  assign key_share0_2_qe = &key_share0_2_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_2_gated_we;
  assign key_share0_2_gated_we = key_share0_2_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_2 (
    .re     (1'b0),
    .we     (key_share0_2_gated_we),
    .wd     (key_share0_2_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_2_flds_we[0]),
    .q      (reg2hw.key_share0[2].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[2].qe = key_share0_2_qe;


  // Subregister 3 of Multireg key_share0
  // R[key_share0_3]: V(True)
  logic key_share0_3_qe;
  logic [0:0] key_share0_3_flds_we;
  assign key_share0_3_qe = &key_share0_3_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_3_gated_we;
  assign key_share0_3_gated_we = key_share0_3_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_3 (
    .re     (1'b0),
    .we     (key_share0_3_gated_we),
    .wd     (key_share0_3_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_3_flds_we[0]),
    .q      (reg2hw.key_share0[3].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[3].qe = key_share0_3_qe;


  // Subregister 4 of Multireg key_share0
  // R[key_share0_4]: V(True)
  logic key_share0_4_qe;
  logic [0:0] key_share0_4_flds_we;
  assign key_share0_4_qe = &key_share0_4_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_4_gated_we;
  assign key_share0_4_gated_we = key_share0_4_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_4 (
    .re     (1'b0),
    .we     (key_share0_4_gated_we),
    .wd     (key_share0_4_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_4_flds_we[0]),
    .q      (reg2hw.key_share0[4].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[4].qe = key_share0_4_qe;


  // Subregister 5 of Multireg key_share0
  // R[key_share0_5]: V(True)
  logic key_share0_5_qe;
  logic [0:0] key_share0_5_flds_we;
  assign key_share0_5_qe = &key_share0_5_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_5_gated_we;
  assign key_share0_5_gated_we = key_share0_5_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_5 (
    .re     (1'b0),
    .we     (key_share0_5_gated_we),
    .wd     (key_share0_5_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_5_flds_we[0]),
    .q      (reg2hw.key_share0[5].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[5].qe = key_share0_5_qe;


  // Subregister 6 of Multireg key_share0
  // R[key_share0_6]: V(True)
  logic key_share0_6_qe;
  logic [0:0] key_share0_6_flds_we;
  assign key_share0_6_qe = &key_share0_6_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_6_gated_we;
  assign key_share0_6_gated_we = key_share0_6_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_6 (
    .re     (1'b0),
    .we     (key_share0_6_gated_we),
    .wd     (key_share0_6_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_6_flds_we[0]),
    .q      (reg2hw.key_share0[6].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[6].qe = key_share0_6_qe;


  // Subregister 7 of Multireg key_share0
  // R[key_share0_7]: V(True)
  logic key_share0_7_qe;
  logic [0:0] key_share0_7_flds_we;
  assign key_share0_7_qe = &key_share0_7_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_7_gated_we;
  assign key_share0_7_gated_we = key_share0_7_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_7 (
    .re     (1'b0),
    .we     (key_share0_7_gated_we),
    .wd     (key_share0_7_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_7_flds_we[0]),
    .q      (reg2hw.key_share0[7].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[7].qe = key_share0_7_qe;


  // Subregister 8 of Multireg key_share0
  // R[key_share0_8]: V(True)
  logic key_share0_8_qe;
  logic [0:0] key_share0_8_flds_we;
  assign key_share0_8_qe = &key_share0_8_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_8_gated_we;
  assign key_share0_8_gated_we = key_share0_8_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_8 (
    .re     (1'b0),
    .we     (key_share0_8_gated_we),
    .wd     (key_share0_8_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_8_flds_we[0]),
    .q      (reg2hw.key_share0[8].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[8].qe = key_share0_8_qe;


  // Subregister 9 of Multireg key_share0
  // R[key_share0_9]: V(True)
  logic key_share0_9_qe;
  logic [0:0] key_share0_9_flds_we;
  assign key_share0_9_qe = &key_share0_9_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_9_gated_we;
  assign key_share0_9_gated_we = key_share0_9_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_9 (
    .re     (1'b0),
    .we     (key_share0_9_gated_we),
    .wd     (key_share0_9_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_9_flds_we[0]),
    .q      (reg2hw.key_share0[9].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[9].qe = key_share0_9_qe;


  // Subregister 10 of Multireg key_share0
  // R[key_share0_10]: V(True)
  logic key_share0_10_qe;
  logic [0:0] key_share0_10_flds_we;
  assign key_share0_10_qe = &key_share0_10_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_10_gated_we;
  assign key_share0_10_gated_we = key_share0_10_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_10 (
    .re     (1'b0),
    .we     (key_share0_10_gated_we),
    .wd     (key_share0_10_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_10_flds_we[0]),
    .q      (reg2hw.key_share0[10].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[10].qe = key_share0_10_qe;


  // Subregister 11 of Multireg key_share0
  // R[key_share0_11]: V(True)
  logic key_share0_11_qe;
  logic [0:0] key_share0_11_flds_we;
  assign key_share0_11_qe = &key_share0_11_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_11_gated_we;
  assign key_share0_11_gated_we = key_share0_11_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_11 (
    .re     (1'b0),
    .we     (key_share0_11_gated_we),
    .wd     (key_share0_11_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_11_flds_we[0]),
    .q      (reg2hw.key_share0[11].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[11].qe = key_share0_11_qe;


  // Subregister 12 of Multireg key_share0
  // R[key_share0_12]: V(True)
  logic key_share0_12_qe;
  logic [0:0] key_share0_12_flds_we;
  assign key_share0_12_qe = &key_share0_12_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_12_gated_we;
  assign key_share0_12_gated_we = key_share0_12_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_12 (
    .re     (1'b0),
    .we     (key_share0_12_gated_we),
    .wd     (key_share0_12_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_12_flds_we[0]),
    .q      (reg2hw.key_share0[12].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[12].qe = key_share0_12_qe;


  // Subregister 13 of Multireg key_share0
  // R[key_share0_13]: V(True)
  logic key_share0_13_qe;
  logic [0:0] key_share0_13_flds_we;
  assign key_share0_13_qe = &key_share0_13_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_13_gated_we;
  assign key_share0_13_gated_we = key_share0_13_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_13 (
    .re     (1'b0),
    .we     (key_share0_13_gated_we),
    .wd     (key_share0_13_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_13_flds_we[0]),
    .q      (reg2hw.key_share0[13].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[13].qe = key_share0_13_qe;


  // Subregister 14 of Multireg key_share0
  // R[key_share0_14]: V(True)
  logic key_share0_14_qe;
  logic [0:0] key_share0_14_flds_we;
  assign key_share0_14_qe = &key_share0_14_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_14_gated_we;
  assign key_share0_14_gated_we = key_share0_14_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_14 (
    .re     (1'b0),
    .we     (key_share0_14_gated_we),
    .wd     (key_share0_14_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_14_flds_we[0]),
    .q      (reg2hw.key_share0[14].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[14].qe = key_share0_14_qe;


  // Subregister 15 of Multireg key_share0
  // R[key_share0_15]: V(True)
  logic key_share0_15_qe;
  logic [0:0] key_share0_15_flds_we;
  assign key_share0_15_qe = &key_share0_15_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share0_15_gated_we;
  assign key_share0_15_gated_we = key_share0_15_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share0_15 (
    .re     (1'b0),
    .we     (key_share0_15_gated_we),
    .wd     (key_share0_15_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share0_15_flds_we[0]),
    .q      (reg2hw.key_share0[15].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share0[15].qe = key_share0_15_qe;


  // Subregister 0 of Multireg key_share1
  // R[key_share1_0]: V(True)
  logic key_share1_0_qe;
  logic [0:0] key_share1_0_flds_we;
  assign key_share1_0_qe = &key_share1_0_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_0_gated_we;
  assign key_share1_0_gated_we = key_share1_0_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_0 (
    .re     (1'b0),
    .we     (key_share1_0_gated_we),
    .wd     (key_share1_0_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_0_flds_we[0]),
    .q      (reg2hw.key_share1[0].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[0].qe = key_share1_0_qe;


  // Subregister 1 of Multireg key_share1
  // R[key_share1_1]: V(True)
  logic key_share1_1_qe;
  logic [0:0] key_share1_1_flds_we;
  assign key_share1_1_qe = &key_share1_1_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_1_gated_we;
  assign key_share1_1_gated_we = key_share1_1_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_1 (
    .re     (1'b0),
    .we     (key_share1_1_gated_we),
    .wd     (key_share1_1_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_1_flds_we[0]),
    .q      (reg2hw.key_share1[1].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[1].qe = key_share1_1_qe;


  // Subregister 2 of Multireg key_share1
  // R[key_share1_2]: V(True)
  logic key_share1_2_qe;
  logic [0:0] key_share1_2_flds_we;
  assign key_share1_2_qe = &key_share1_2_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_2_gated_we;
  assign key_share1_2_gated_we = key_share1_2_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_2 (
    .re     (1'b0),
    .we     (key_share1_2_gated_we),
    .wd     (key_share1_2_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_2_flds_we[0]),
    .q      (reg2hw.key_share1[2].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[2].qe = key_share1_2_qe;


  // Subregister 3 of Multireg key_share1
  // R[key_share1_3]: V(True)
  logic key_share1_3_qe;
  logic [0:0] key_share1_3_flds_we;
  assign key_share1_3_qe = &key_share1_3_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_3_gated_we;
  assign key_share1_3_gated_we = key_share1_3_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_3 (
    .re     (1'b0),
    .we     (key_share1_3_gated_we),
    .wd     (key_share1_3_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_3_flds_we[0]),
    .q      (reg2hw.key_share1[3].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[3].qe = key_share1_3_qe;


  // Subregister 4 of Multireg key_share1
  // R[key_share1_4]: V(True)
  logic key_share1_4_qe;
  logic [0:0] key_share1_4_flds_we;
  assign key_share1_4_qe = &key_share1_4_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_4_gated_we;
  assign key_share1_4_gated_we = key_share1_4_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_4 (
    .re     (1'b0),
    .we     (key_share1_4_gated_we),
    .wd     (key_share1_4_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_4_flds_we[0]),
    .q      (reg2hw.key_share1[4].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[4].qe = key_share1_4_qe;


  // Subregister 5 of Multireg key_share1
  // R[key_share1_5]: V(True)
  logic key_share1_5_qe;
  logic [0:0] key_share1_5_flds_we;
  assign key_share1_5_qe = &key_share1_5_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_5_gated_we;
  assign key_share1_5_gated_we = key_share1_5_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_5 (
    .re     (1'b0),
    .we     (key_share1_5_gated_we),
    .wd     (key_share1_5_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_5_flds_we[0]),
    .q      (reg2hw.key_share1[5].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[5].qe = key_share1_5_qe;


  // Subregister 6 of Multireg key_share1
  // R[key_share1_6]: V(True)
  logic key_share1_6_qe;
  logic [0:0] key_share1_6_flds_we;
  assign key_share1_6_qe = &key_share1_6_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_6_gated_we;
  assign key_share1_6_gated_we = key_share1_6_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_6 (
    .re     (1'b0),
    .we     (key_share1_6_gated_we),
    .wd     (key_share1_6_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_6_flds_we[0]),
    .q      (reg2hw.key_share1[6].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[6].qe = key_share1_6_qe;


  // Subregister 7 of Multireg key_share1
  // R[key_share1_7]: V(True)
  logic key_share1_7_qe;
  logic [0:0] key_share1_7_flds_we;
  assign key_share1_7_qe = &key_share1_7_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_7_gated_we;
  assign key_share1_7_gated_we = key_share1_7_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_7 (
    .re     (1'b0),
    .we     (key_share1_7_gated_we),
    .wd     (key_share1_7_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_7_flds_we[0]),
    .q      (reg2hw.key_share1[7].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[7].qe = key_share1_7_qe;


  // Subregister 8 of Multireg key_share1
  // R[key_share1_8]: V(True)
  logic key_share1_8_qe;
  logic [0:0] key_share1_8_flds_we;
  assign key_share1_8_qe = &key_share1_8_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_8_gated_we;
  assign key_share1_8_gated_we = key_share1_8_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_8 (
    .re     (1'b0),
    .we     (key_share1_8_gated_we),
    .wd     (key_share1_8_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_8_flds_we[0]),
    .q      (reg2hw.key_share1[8].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[8].qe = key_share1_8_qe;


  // Subregister 9 of Multireg key_share1
  // R[key_share1_9]: V(True)
  logic key_share1_9_qe;
  logic [0:0] key_share1_9_flds_we;
  assign key_share1_9_qe = &key_share1_9_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_9_gated_we;
  assign key_share1_9_gated_we = key_share1_9_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_9 (
    .re     (1'b0),
    .we     (key_share1_9_gated_we),
    .wd     (key_share1_9_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_9_flds_we[0]),
    .q      (reg2hw.key_share1[9].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[9].qe = key_share1_9_qe;


  // Subregister 10 of Multireg key_share1
  // R[key_share1_10]: V(True)
  logic key_share1_10_qe;
  logic [0:0] key_share1_10_flds_we;
  assign key_share1_10_qe = &key_share1_10_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_10_gated_we;
  assign key_share1_10_gated_we = key_share1_10_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_10 (
    .re     (1'b0),
    .we     (key_share1_10_gated_we),
    .wd     (key_share1_10_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_10_flds_we[0]),
    .q      (reg2hw.key_share1[10].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[10].qe = key_share1_10_qe;


  // Subregister 11 of Multireg key_share1
  // R[key_share1_11]: V(True)
  logic key_share1_11_qe;
  logic [0:0] key_share1_11_flds_we;
  assign key_share1_11_qe = &key_share1_11_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_11_gated_we;
  assign key_share1_11_gated_we = key_share1_11_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_11 (
    .re     (1'b0),
    .we     (key_share1_11_gated_we),
    .wd     (key_share1_11_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_11_flds_we[0]),
    .q      (reg2hw.key_share1[11].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[11].qe = key_share1_11_qe;


  // Subregister 12 of Multireg key_share1
  // R[key_share1_12]: V(True)
  logic key_share1_12_qe;
  logic [0:0] key_share1_12_flds_we;
  assign key_share1_12_qe = &key_share1_12_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_12_gated_we;
  assign key_share1_12_gated_we = key_share1_12_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_12 (
    .re     (1'b0),
    .we     (key_share1_12_gated_we),
    .wd     (key_share1_12_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_12_flds_we[0]),
    .q      (reg2hw.key_share1[12].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[12].qe = key_share1_12_qe;


  // Subregister 13 of Multireg key_share1
  // R[key_share1_13]: V(True)
  logic key_share1_13_qe;
  logic [0:0] key_share1_13_flds_we;
  assign key_share1_13_qe = &key_share1_13_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_13_gated_we;
  assign key_share1_13_gated_we = key_share1_13_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_13 (
    .re     (1'b0),
    .we     (key_share1_13_gated_we),
    .wd     (key_share1_13_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_13_flds_we[0]),
    .q      (reg2hw.key_share1[13].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[13].qe = key_share1_13_qe;


  // Subregister 14 of Multireg key_share1
  // R[key_share1_14]: V(True)
  logic key_share1_14_qe;
  logic [0:0] key_share1_14_flds_we;
  assign key_share1_14_qe = &key_share1_14_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_14_gated_we;
  assign key_share1_14_gated_we = key_share1_14_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_14 (
    .re     (1'b0),
    .we     (key_share1_14_gated_we),
    .wd     (key_share1_14_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_14_flds_we[0]),
    .q      (reg2hw.key_share1[14].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[14].qe = key_share1_14_qe;


  // Subregister 15 of Multireg key_share1
  // R[key_share1_15]: V(True)
  logic key_share1_15_qe;
  logic [0:0] key_share1_15_flds_we;
  assign key_share1_15_qe = &key_share1_15_flds_we;
  // Create REGWEN-gated WE signal
  logic key_share1_15_gated_we;
  assign key_share1_15_gated_we = key_share1_15_we & cfg_regwen_qs;
  prim_subreg_ext #(
    .DW    (32)
  ) u_key_share1_15 (
    .re     (1'b0),
    .we     (key_share1_15_gated_we),
    .wd     (key_share1_15_wd),
    .d      ('0),
    .qre    (),
    .qe     (key_share1_15_flds_we[0]),
    .q      (reg2hw.key_share1[15].q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.key_share1[15].qe = key_share1_15_qe;


  // R[key_len]: V(False)
  // Create REGWEN-gated WE signal
  logic key_len_gated_we;
  assign key_len_gated_we = key_len_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (3),
    .SwAccess(prim_subreg_pkg::SwAccessWO),
    .RESVAL  (3'h0)
  ) u_key_len (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (key_len_gated_we),
    .wd     (key_len_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.key_len.q),
    .ds     (),

    // to register interface (read)
    .qs     ()
  );


  // Subregister 0 of Multireg prefix
  // R[prefix_0]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_0_gated_we;
  assign prefix_0_gated_we = prefix_0_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_0_gated_we),
    .wd     (prefix_0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_0_qs)
  );


  // Subregister 1 of Multireg prefix
  // R[prefix_1]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_1_gated_we;
  assign prefix_1_gated_we = prefix_1_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_1_gated_we),
    .wd     (prefix_1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_1_qs)
  );


  // Subregister 2 of Multireg prefix
  // R[prefix_2]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_2_gated_we;
  assign prefix_2_gated_we = prefix_2_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_2_gated_we),
    .wd     (prefix_2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_2_qs)
  );


  // Subregister 3 of Multireg prefix
  // R[prefix_3]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_3_gated_we;
  assign prefix_3_gated_we = prefix_3_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_3_gated_we),
    .wd     (prefix_3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_3_qs)
  );


  // Subregister 4 of Multireg prefix
  // R[prefix_4]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_4_gated_we;
  assign prefix_4_gated_we = prefix_4_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_4_gated_we),
    .wd     (prefix_4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_4_qs)
  );


  // Subregister 5 of Multireg prefix
  // R[prefix_5]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_5_gated_we;
  assign prefix_5_gated_we = prefix_5_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_5_gated_we),
    .wd     (prefix_5_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_5_qs)
  );


  // Subregister 6 of Multireg prefix
  // R[prefix_6]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_6_gated_we;
  assign prefix_6_gated_we = prefix_6_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_6_gated_we),
    .wd     (prefix_6_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_6_qs)
  );


  // Subregister 7 of Multireg prefix
  // R[prefix_7]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_7_gated_we;
  assign prefix_7_gated_we = prefix_7_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_7_gated_we),
    .wd     (prefix_7_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_7_qs)
  );


  // Subregister 8 of Multireg prefix
  // R[prefix_8]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_8_gated_we;
  assign prefix_8_gated_we = prefix_8_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_8 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_8_gated_we),
    .wd     (prefix_8_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[8].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_8_qs)
  );


  // Subregister 9 of Multireg prefix
  // R[prefix_9]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_9_gated_we;
  assign prefix_9_gated_we = prefix_9_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_9 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_9_gated_we),
    .wd     (prefix_9_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[9].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_9_qs)
  );


  // Subregister 10 of Multireg prefix
  // R[prefix_10]: V(False)
  // Create REGWEN-gated WE signal
  logic prefix_10_gated_we;
  assign prefix_10_gated_we = prefix_10_we & cfg_regwen_qs;
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_prefix_10 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (prefix_10_gated_we),
    .wd     (prefix_10_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.prefix[10].q),
    .ds     (),

    // to register interface (read)
    .qs     (prefix_10_qs)
  );


  // R[err_code]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_err_code (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.err_code.de),
    .d      (hw2reg.err_code.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (err_code_qs)
  );



  logic [60:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == KMAC_INTR_STATE_OFFSET);
    addr_hit[ 1] = (reg_addr == KMAC_INTR_ENABLE_OFFSET);
    addr_hit[ 2] = (reg_addr == KMAC_INTR_TEST_OFFSET);
    addr_hit[ 3] = (reg_addr == KMAC_ALERT_TEST_OFFSET);
    addr_hit[ 4] = (reg_addr == KMAC_CFG_REGWEN_OFFSET);
    addr_hit[ 5] = (reg_addr == KMAC_CFG_SHADOWED_OFFSET);
    addr_hit[ 6] = (reg_addr == KMAC_CMD_OFFSET);
    addr_hit[ 7] = (reg_addr == KMAC_STATUS_OFFSET);
    addr_hit[ 8] = (reg_addr == KMAC_ENTROPY_PERIOD_OFFSET);
    addr_hit[ 9] = (reg_addr == KMAC_ENTROPY_REFRESH_HASH_CNT_OFFSET);
    addr_hit[10] = (reg_addr == KMAC_ENTROPY_REFRESH_THRESHOLD_SHADOWED_OFFSET);
    addr_hit[11] = (reg_addr == KMAC_ENTROPY_SEED_0_OFFSET);
    addr_hit[12] = (reg_addr == KMAC_ENTROPY_SEED_1_OFFSET);
    addr_hit[13] = (reg_addr == KMAC_ENTROPY_SEED_2_OFFSET);
    addr_hit[14] = (reg_addr == KMAC_ENTROPY_SEED_3_OFFSET);
    addr_hit[15] = (reg_addr == KMAC_ENTROPY_SEED_4_OFFSET);
    addr_hit[16] = (reg_addr == KMAC_KEY_SHARE0_0_OFFSET);
    addr_hit[17] = (reg_addr == KMAC_KEY_SHARE0_1_OFFSET);
    addr_hit[18] = (reg_addr == KMAC_KEY_SHARE0_2_OFFSET);
    addr_hit[19] = (reg_addr == KMAC_KEY_SHARE0_3_OFFSET);
    addr_hit[20] = (reg_addr == KMAC_KEY_SHARE0_4_OFFSET);
    addr_hit[21] = (reg_addr == KMAC_KEY_SHARE0_5_OFFSET);
    addr_hit[22] = (reg_addr == KMAC_KEY_SHARE0_6_OFFSET);
    addr_hit[23] = (reg_addr == KMAC_KEY_SHARE0_7_OFFSET);
    addr_hit[24] = (reg_addr == KMAC_KEY_SHARE0_8_OFFSET);
    addr_hit[25] = (reg_addr == KMAC_KEY_SHARE0_9_OFFSET);
    addr_hit[26] = (reg_addr == KMAC_KEY_SHARE0_10_OFFSET);
    addr_hit[27] = (reg_addr == KMAC_KEY_SHARE0_11_OFFSET);
    addr_hit[28] = (reg_addr == KMAC_KEY_SHARE0_12_OFFSET);
    addr_hit[29] = (reg_addr == KMAC_KEY_SHARE0_13_OFFSET);
    addr_hit[30] = (reg_addr == KMAC_KEY_SHARE0_14_OFFSET);
    addr_hit[31] = (reg_addr == KMAC_KEY_SHARE0_15_OFFSET);
    addr_hit[32] = (reg_addr == KMAC_KEY_SHARE1_0_OFFSET);
    addr_hit[33] = (reg_addr == KMAC_KEY_SHARE1_1_OFFSET);
    addr_hit[34] = (reg_addr == KMAC_KEY_SHARE1_2_OFFSET);
    addr_hit[35] = (reg_addr == KMAC_KEY_SHARE1_3_OFFSET);
    addr_hit[36] = (reg_addr == KMAC_KEY_SHARE1_4_OFFSET);
    addr_hit[37] = (reg_addr == KMAC_KEY_SHARE1_5_OFFSET);
    addr_hit[38] = (reg_addr == KMAC_KEY_SHARE1_6_OFFSET);
    addr_hit[39] = (reg_addr == KMAC_KEY_SHARE1_7_OFFSET);
    addr_hit[40] = (reg_addr == KMAC_KEY_SHARE1_8_OFFSET);
    addr_hit[41] = (reg_addr == KMAC_KEY_SHARE1_9_OFFSET);
    addr_hit[42] = (reg_addr == KMAC_KEY_SHARE1_10_OFFSET);
    addr_hit[43] = (reg_addr == KMAC_KEY_SHARE1_11_OFFSET);
    addr_hit[44] = (reg_addr == KMAC_KEY_SHARE1_12_OFFSET);
    addr_hit[45] = (reg_addr == KMAC_KEY_SHARE1_13_OFFSET);
    addr_hit[46] = (reg_addr == KMAC_KEY_SHARE1_14_OFFSET);
    addr_hit[47] = (reg_addr == KMAC_KEY_SHARE1_15_OFFSET);
    addr_hit[48] = (reg_addr == KMAC_KEY_LEN_OFFSET);
    addr_hit[49] = (reg_addr == KMAC_PREFIX_0_OFFSET);
    addr_hit[50] = (reg_addr == KMAC_PREFIX_1_OFFSET);
    addr_hit[51] = (reg_addr == KMAC_PREFIX_2_OFFSET);
    addr_hit[52] = (reg_addr == KMAC_PREFIX_3_OFFSET);
    addr_hit[53] = (reg_addr == KMAC_PREFIX_4_OFFSET);
    addr_hit[54] = (reg_addr == KMAC_PREFIX_5_OFFSET);
    addr_hit[55] = (reg_addr == KMAC_PREFIX_6_OFFSET);
    addr_hit[56] = (reg_addr == KMAC_PREFIX_7_OFFSET);
    addr_hit[57] = (reg_addr == KMAC_PREFIX_8_OFFSET);
    addr_hit[58] = (reg_addr == KMAC_PREFIX_9_OFFSET);
    addr_hit[59] = (reg_addr == KMAC_PREFIX_10_OFFSET);
    addr_hit[60] = (reg_addr == KMAC_ERR_CODE_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(KMAC_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(KMAC_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(KMAC_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(KMAC_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(KMAC_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(KMAC_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(KMAC_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(KMAC_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(KMAC_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(KMAC_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(KMAC_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(KMAC_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(KMAC_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(KMAC_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(KMAC_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(KMAC_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(KMAC_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(KMAC_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(KMAC_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(KMAC_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(KMAC_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(KMAC_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(KMAC_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(KMAC_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(KMAC_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(KMAC_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(KMAC_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(KMAC_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(KMAC_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(KMAC_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(KMAC_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(KMAC_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(KMAC_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(KMAC_PERMIT[33] & ~reg_be))) |
               (addr_hit[34] & (|(KMAC_PERMIT[34] & ~reg_be))) |
               (addr_hit[35] & (|(KMAC_PERMIT[35] & ~reg_be))) |
               (addr_hit[36] & (|(KMAC_PERMIT[36] & ~reg_be))) |
               (addr_hit[37] & (|(KMAC_PERMIT[37] & ~reg_be))) |
               (addr_hit[38] & (|(KMAC_PERMIT[38] & ~reg_be))) |
               (addr_hit[39] & (|(KMAC_PERMIT[39] & ~reg_be))) |
               (addr_hit[40] & (|(KMAC_PERMIT[40] & ~reg_be))) |
               (addr_hit[41] & (|(KMAC_PERMIT[41] & ~reg_be))) |
               (addr_hit[42] & (|(KMAC_PERMIT[42] & ~reg_be))) |
               (addr_hit[43] & (|(KMAC_PERMIT[43] & ~reg_be))) |
               (addr_hit[44] & (|(KMAC_PERMIT[44] & ~reg_be))) |
               (addr_hit[45] & (|(KMAC_PERMIT[45] & ~reg_be))) |
               (addr_hit[46] & (|(KMAC_PERMIT[46] & ~reg_be))) |
               (addr_hit[47] & (|(KMAC_PERMIT[47] & ~reg_be))) |
               (addr_hit[48] & (|(KMAC_PERMIT[48] & ~reg_be))) |
               (addr_hit[49] & (|(KMAC_PERMIT[49] & ~reg_be))) |
               (addr_hit[50] & (|(KMAC_PERMIT[50] & ~reg_be))) |
               (addr_hit[51] & (|(KMAC_PERMIT[51] & ~reg_be))) |
               (addr_hit[52] & (|(KMAC_PERMIT[52] & ~reg_be))) |
               (addr_hit[53] & (|(KMAC_PERMIT[53] & ~reg_be))) |
               (addr_hit[54] & (|(KMAC_PERMIT[54] & ~reg_be))) |
               (addr_hit[55] & (|(KMAC_PERMIT[55] & ~reg_be))) |
               (addr_hit[56] & (|(KMAC_PERMIT[56] & ~reg_be))) |
               (addr_hit[57] & (|(KMAC_PERMIT[57] & ~reg_be))) |
               (addr_hit[58] & (|(KMAC_PERMIT[58] & ~reg_be))) |
               (addr_hit[59] & (|(KMAC_PERMIT[59] & ~reg_be))) |
               (addr_hit[60] & (|(KMAC_PERMIT[60] & ~reg_be)))));
  end

  // Generate write-enables
  assign intr_state_we = addr_hit[0] & reg_we & !reg_error;

  assign intr_state_kmac_done_wd = reg_wdata[0];

  assign intr_state_fifo_empty_wd = reg_wdata[1];

  assign intr_state_kmac_err_wd = reg_wdata[2];
  assign intr_enable_we = addr_hit[1] & reg_we & !reg_error;

  assign intr_enable_kmac_done_wd = reg_wdata[0];

  assign intr_enable_fifo_empty_wd = reg_wdata[1];

  assign intr_enable_kmac_err_wd = reg_wdata[2];
  assign intr_test_we = addr_hit[2] & reg_we & !reg_error;

  assign intr_test_kmac_done_wd = reg_wdata[0];

  assign intr_test_fifo_empty_wd = reg_wdata[1];

  assign intr_test_kmac_err_wd = reg_wdata[2];
  assign alert_test_we = addr_hit[3] & reg_we & !reg_error;

  assign alert_test_recov_operation_err_wd = reg_wdata[0];

  assign alert_test_fatal_fault_err_wd = reg_wdata[1];
  assign cfg_regwen_re = addr_hit[4] & reg_re & !reg_error;
  assign cfg_shadowed_re = addr_hit[5] & reg_re & !reg_error;
  assign cfg_shadowed_we = addr_hit[5] & reg_we & !reg_error;

  assign cfg_shadowed_kmac_en_wd = reg_wdata[0];

  assign cfg_shadowed_kstrength_wd = reg_wdata[3:1];

  assign cfg_shadowed_mode_wd = reg_wdata[5:4];

  assign cfg_shadowed_msg_endianness_wd = reg_wdata[8];

  assign cfg_shadowed_state_endianness_wd = reg_wdata[9];

  assign cfg_shadowed_sideload_wd = reg_wdata[12];

  assign cfg_shadowed_entropy_mode_wd = reg_wdata[17:16];

  assign cfg_shadowed_entropy_fast_process_wd = reg_wdata[19];

  assign cfg_shadowed_msg_mask_wd = reg_wdata[20];

  assign cfg_shadowed_entropy_ready_wd = reg_wdata[24];

  assign cfg_shadowed_err_processed_wd = reg_wdata[25];

  assign cfg_shadowed_en_unsupported_modestrength_wd = reg_wdata[26];
  assign cmd_we = addr_hit[6] & reg_we & !reg_error;

  assign cmd_cmd_wd = reg_wdata[5:0];

  assign cmd_entropy_req_wd = reg_wdata[8];

  assign cmd_hash_cnt_clr_wd = reg_wdata[9];
  assign status_re = addr_hit[7] & reg_re & !reg_error;
  assign entropy_period_we = addr_hit[8] & reg_we & !reg_error;

  assign entropy_period_prescaler_wd = reg_wdata[9:0];

  assign entropy_period_wait_timer_wd = reg_wdata[31:16];
  assign entropy_refresh_threshold_shadowed_re = addr_hit[10] & reg_re & !reg_error;
  assign entropy_refresh_threshold_shadowed_we = addr_hit[10] & reg_we & !reg_error;

  assign entropy_refresh_threshold_shadowed_wd = reg_wdata[9:0];
  assign entropy_seed_0_we = addr_hit[11] & reg_we & !reg_error;

  assign entropy_seed_0_wd = reg_wdata[31:0];
  assign entropy_seed_1_we = addr_hit[12] & reg_we & !reg_error;

  assign entropy_seed_1_wd = reg_wdata[31:0];
  assign entropy_seed_2_we = addr_hit[13] & reg_we & !reg_error;

  assign entropy_seed_2_wd = reg_wdata[31:0];
  assign entropy_seed_3_we = addr_hit[14] & reg_we & !reg_error;

  assign entropy_seed_3_wd = reg_wdata[31:0];
  assign entropy_seed_4_we = addr_hit[15] & reg_we & !reg_error;

  assign entropy_seed_4_wd = reg_wdata[31:0];
  assign key_share0_0_we = addr_hit[16] & reg_we & !reg_error;

  assign key_share0_0_wd = reg_wdata[31:0];
  assign key_share0_1_we = addr_hit[17] & reg_we & !reg_error;

  assign key_share0_1_wd = reg_wdata[31:0];
  assign key_share0_2_we = addr_hit[18] & reg_we & !reg_error;

  assign key_share0_2_wd = reg_wdata[31:0];
  assign key_share0_3_we = addr_hit[19] & reg_we & !reg_error;

  assign key_share0_3_wd = reg_wdata[31:0];
  assign key_share0_4_we = addr_hit[20] & reg_we & !reg_error;

  assign key_share0_4_wd = reg_wdata[31:0];
  assign key_share0_5_we = addr_hit[21] & reg_we & !reg_error;

  assign key_share0_5_wd = reg_wdata[31:0];
  assign key_share0_6_we = addr_hit[22] & reg_we & !reg_error;

  assign key_share0_6_wd = reg_wdata[31:0];
  assign key_share0_7_we = addr_hit[23] & reg_we & !reg_error;

  assign key_share0_7_wd = reg_wdata[31:0];
  assign key_share0_8_we = addr_hit[24] & reg_we & !reg_error;

  assign key_share0_8_wd = reg_wdata[31:0];
  assign key_share0_9_we = addr_hit[25] & reg_we & !reg_error;

  assign key_share0_9_wd = reg_wdata[31:0];
  assign key_share0_10_we = addr_hit[26] & reg_we & !reg_error;

  assign key_share0_10_wd = reg_wdata[31:0];
  assign key_share0_11_we = addr_hit[27] & reg_we & !reg_error;

  assign key_share0_11_wd = reg_wdata[31:0];
  assign key_share0_12_we = addr_hit[28] & reg_we & !reg_error;

  assign key_share0_12_wd = reg_wdata[31:0];
  assign key_share0_13_we = addr_hit[29] & reg_we & !reg_error;

  assign key_share0_13_wd = reg_wdata[31:0];
  assign key_share0_14_we = addr_hit[30] & reg_we & !reg_error;

  assign key_share0_14_wd = reg_wdata[31:0];
  assign key_share0_15_we = addr_hit[31] & reg_we & !reg_error;

  assign key_share0_15_wd = reg_wdata[31:0];
  assign key_share1_0_we = addr_hit[32] & reg_we & !reg_error;

  assign key_share1_0_wd = reg_wdata[31:0];
  assign key_share1_1_we = addr_hit[33] & reg_we & !reg_error;

  assign key_share1_1_wd = reg_wdata[31:0];
  assign key_share1_2_we = addr_hit[34] & reg_we & !reg_error;

  assign key_share1_2_wd = reg_wdata[31:0];
  assign key_share1_3_we = addr_hit[35] & reg_we & !reg_error;

  assign key_share1_3_wd = reg_wdata[31:0];
  assign key_share1_4_we = addr_hit[36] & reg_we & !reg_error;

  assign key_share1_4_wd = reg_wdata[31:0];
  assign key_share1_5_we = addr_hit[37] & reg_we & !reg_error;

  assign key_share1_5_wd = reg_wdata[31:0];
  assign key_share1_6_we = addr_hit[38] & reg_we & !reg_error;

  assign key_share1_6_wd = reg_wdata[31:0];
  assign key_share1_7_we = addr_hit[39] & reg_we & !reg_error;

  assign key_share1_7_wd = reg_wdata[31:0];
  assign key_share1_8_we = addr_hit[40] & reg_we & !reg_error;

  assign key_share1_8_wd = reg_wdata[31:0];
  assign key_share1_9_we = addr_hit[41] & reg_we & !reg_error;

  assign key_share1_9_wd = reg_wdata[31:0];
  assign key_share1_10_we = addr_hit[42] & reg_we & !reg_error;

  assign key_share1_10_wd = reg_wdata[31:0];
  assign key_share1_11_we = addr_hit[43] & reg_we & !reg_error;

  assign key_share1_11_wd = reg_wdata[31:0];
  assign key_share1_12_we = addr_hit[44] & reg_we & !reg_error;

  assign key_share1_12_wd = reg_wdata[31:0];
  assign key_share1_13_we = addr_hit[45] & reg_we & !reg_error;

  assign key_share1_13_wd = reg_wdata[31:0];
  assign key_share1_14_we = addr_hit[46] & reg_we & !reg_error;

  assign key_share1_14_wd = reg_wdata[31:0];
  assign key_share1_15_we = addr_hit[47] & reg_we & !reg_error;

  assign key_share1_15_wd = reg_wdata[31:0];
  assign key_len_we = addr_hit[48] & reg_we & !reg_error;

  assign key_len_wd = reg_wdata[2:0];
  assign prefix_0_we = addr_hit[49] & reg_we & !reg_error;

  assign prefix_0_wd = reg_wdata[31:0];
  assign prefix_1_we = addr_hit[50] & reg_we & !reg_error;

  assign prefix_1_wd = reg_wdata[31:0];
  assign prefix_2_we = addr_hit[51] & reg_we & !reg_error;

  assign prefix_2_wd = reg_wdata[31:0];
  assign prefix_3_we = addr_hit[52] & reg_we & !reg_error;

  assign prefix_3_wd = reg_wdata[31:0];
  assign prefix_4_we = addr_hit[53] & reg_we & !reg_error;

  assign prefix_4_wd = reg_wdata[31:0];
  assign prefix_5_we = addr_hit[54] & reg_we & !reg_error;

  assign prefix_5_wd = reg_wdata[31:0];
  assign prefix_6_we = addr_hit[55] & reg_we & !reg_error;

  assign prefix_6_wd = reg_wdata[31:0];
  assign prefix_7_we = addr_hit[56] & reg_we & !reg_error;

  assign prefix_7_wd = reg_wdata[31:0];
  assign prefix_8_we = addr_hit[57] & reg_we & !reg_error;

  assign prefix_8_wd = reg_wdata[31:0];
  assign prefix_9_we = addr_hit[58] & reg_we & !reg_error;

  assign prefix_9_wd = reg_wdata[31:0];
  assign prefix_10_we = addr_hit[59] & reg_we & !reg_error;

  assign prefix_10_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = intr_state_we;
    reg_we_check[1] = intr_enable_we;
    reg_we_check[2] = intr_test_we;
    reg_we_check[3] = alert_test_we;
    reg_we_check[4] = 1'b0;
    reg_we_check[5] = cfg_shadowed_gated_we;
    reg_we_check[6] = cmd_we;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = entropy_period_gated_we;
    reg_we_check[9] = 1'b0;
    reg_we_check[10] = entropy_refresh_threshold_shadowed_gated_we;
    reg_we_check[11] = entropy_seed_0_we;
    reg_we_check[12] = entropy_seed_1_we;
    reg_we_check[13] = entropy_seed_2_we;
    reg_we_check[14] = entropy_seed_3_we;
    reg_we_check[15] = entropy_seed_4_we;
    reg_we_check[16] = key_share0_0_gated_we;
    reg_we_check[17] = key_share0_1_gated_we;
    reg_we_check[18] = key_share0_2_gated_we;
    reg_we_check[19] = key_share0_3_gated_we;
    reg_we_check[20] = key_share0_4_gated_we;
    reg_we_check[21] = key_share0_5_gated_we;
    reg_we_check[22] = key_share0_6_gated_we;
    reg_we_check[23] = key_share0_7_gated_we;
    reg_we_check[24] = key_share0_8_gated_we;
    reg_we_check[25] = key_share0_9_gated_we;
    reg_we_check[26] = key_share0_10_gated_we;
    reg_we_check[27] = key_share0_11_gated_we;
    reg_we_check[28] = key_share0_12_gated_we;
    reg_we_check[29] = key_share0_13_gated_we;
    reg_we_check[30] = key_share0_14_gated_we;
    reg_we_check[31] = key_share0_15_gated_we;
    reg_we_check[32] = key_share1_0_gated_we;
    reg_we_check[33] = key_share1_1_gated_we;
    reg_we_check[34] = key_share1_2_gated_we;
    reg_we_check[35] = key_share1_3_gated_we;
    reg_we_check[36] = key_share1_4_gated_we;
    reg_we_check[37] = key_share1_5_gated_we;
    reg_we_check[38] = key_share1_6_gated_we;
    reg_we_check[39] = key_share1_7_gated_we;
    reg_we_check[40] = key_share1_8_gated_we;
    reg_we_check[41] = key_share1_9_gated_we;
    reg_we_check[42] = key_share1_10_gated_we;
    reg_we_check[43] = key_share1_11_gated_we;
    reg_we_check[44] = key_share1_12_gated_we;
    reg_we_check[45] = key_share1_13_gated_we;
    reg_we_check[46] = key_share1_14_gated_we;
    reg_we_check[47] = key_share1_15_gated_we;
    reg_we_check[48] = key_len_gated_we;
    reg_we_check[49] = prefix_0_gated_we;
    reg_we_check[50] = prefix_1_gated_we;
    reg_we_check[51] = prefix_2_gated_we;
    reg_we_check[52] = prefix_3_gated_we;
    reg_we_check[53] = prefix_4_gated_we;
    reg_we_check[54] = prefix_5_gated_we;
    reg_we_check[55] = prefix_6_gated_we;
    reg_we_check[56] = prefix_7_gated_we;
    reg_we_check[57] = prefix_8_gated_we;
    reg_we_check[58] = prefix_9_gated_we;
    reg_we_check[59] = prefix_10_gated_we;
    reg_we_check[60] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = intr_state_kmac_done_qs;
        reg_rdata_next[1] = intr_state_fifo_empty_qs;
        reg_rdata_next[2] = intr_state_kmac_err_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = intr_enable_kmac_done_qs;
        reg_rdata_next[1] = intr_enable_fifo_empty_qs;
        reg_rdata_next[2] = intr_enable_kmac_err_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
        reg_rdata_next[2] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[0] = '0;
        reg_rdata_next[1] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[0] = cfg_regwen_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[0] = cfg_shadowed_kmac_en_qs;
        reg_rdata_next[3:1] = cfg_shadowed_kstrength_qs;
        reg_rdata_next[5:4] = cfg_shadowed_mode_qs;
        reg_rdata_next[8] = cfg_shadowed_msg_endianness_qs;
        reg_rdata_next[9] = cfg_shadowed_state_endianness_qs;
        reg_rdata_next[12] = cfg_shadowed_sideload_qs;
        reg_rdata_next[17:16] = cfg_shadowed_entropy_mode_qs;
        reg_rdata_next[19] = cfg_shadowed_entropy_fast_process_qs;
        reg_rdata_next[20] = cfg_shadowed_msg_mask_qs;
        reg_rdata_next[24] = cfg_shadowed_entropy_ready_qs;
        reg_rdata_next[25] = cfg_shadowed_err_processed_qs;
        reg_rdata_next[26] = cfg_shadowed_en_unsupported_modestrength_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[5:0] = '0;
        reg_rdata_next[8] = '0;
        reg_rdata_next[9] = '0;
      end

      addr_hit[7]: begin
        reg_rdata_next[0] = status_sha3_idle_qs;
        reg_rdata_next[1] = status_sha3_absorb_qs;
        reg_rdata_next[2] = status_sha3_squeeze_qs;
        reg_rdata_next[12:8] = status_fifo_depth_qs;
        reg_rdata_next[14] = status_fifo_empty_qs;
        reg_rdata_next[15] = status_fifo_full_qs;
        reg_rdata_next[16] = status_alert_fatal_fault_qs;
        reg_rdata_next[17] = status_alert_recov_ctrl_update_err_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[9:0] = entropy_period_prescaler_qs;
        reg_rdata_next[31:16] = entropy_period_wait_timer_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[9:0] = entropy_refresh_hash_cnt_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[9:0] = entropy_refresh_threshold_shadowed_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[29]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[30]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[36]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[38]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[40]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[41]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[42]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[43]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[44]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[45]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[46]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[47]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[48]: begin
        reg_rdata_next[2:0] = '0;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = prefix_0_qs;
      end

      addr_hit[50]: begin
        reg_rdata_next[31:0] = prefix_1_qs;
      end

      addr_hit[51]: begin
        reg_rdata_next[31:0] = prefix_2_qs;
      end

      addr_hit[52]: begin
        reg_rdata_next[31:0] = prefix_3_qs;
      end

      addr_hit[53]: begin
        reg_rdata_next[31:0] = prefix_4_qs;
      end

      addr_hit[54]: begin
        reg_rdata_next[31:0] = prefix_5_qs;
      end

      addr_hit[55]: begin
        reg_rdata_next[31:0] = prefix_6_qs;
      end

      addr_hit[56]: begin
        reg_rdata_next[31:0] = prefix_7_qs;
      end

      addr_hit[57]: begin
        reg_rdata_next[31:0] = prefix_8_qs;
      end

      addr_hit[58]: begin
        reg_rdata_next[31:0] = prefix_9_qs;
      end

      addr_hit[59]: begin
        reg_rdata_next[31:0] = prefix_10_qs;
      end

      addr_hit[60]: begin
        reg_rdata_next[31:0] = err_code_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  logic rst_done;
  logic shadow_rst_done;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rst_done <= '0;
    end else begin
      rst_done <= 1'b1;
    end
  end

  always_ff @(posedge clk_i or negedge rst_shadowed_ni) begin
    if (!rst_shadowed_ni) begin
      shadow_rst_done <= '0;
    end else begin
      shadow_rst_done <= 1'b1;
    end
  end

  // both shadow and normal resets have been released
  assign shadow_busy = ~(rst_done & shadow_rst_done);

  // Collect up storage and update errors
  assign shadowed_storage_err_o = |{
    cfg_shadowed_kmac_en_storage_err,
    cfg_shadowed_kstrength_storage_err,
    cfg_shadowed_mode_storage_err,
    cfg_shadowed_msg_endianness_storage_err,
    cfg_shadowed_state_endianness_storage_err,
    cfg_shadowed_sideload_storage_err,
    cfg_shadowed_entropy_mode_storage_err,
    cfg_shadowed_entropy_fast_process_storage_err,
    cfg_shadowed_msg_mask_storage_err,
    cfg_shadowed_entropy_ready_storage_err,
    cfg_shadowed_err_processed_storage_err,
    cfg_shadowed_en_unsupported_modestrength_storage_err,
    entropy_refresh_threshold_shadowed_storage_err
  };
  assign shadowed_update_err_o = |{
    cfg_shadowed_kmac_en_update_err,
    cfg_shadowed_kstrength_update_err,
    cfg_shadowed_mode_update_err,
    cfg_shadowed_msg_endianness_update_err,
    cfg_shadowed_state_endianness_update_err,
    cfg_shadowed_sideload_update_err,
    cfg_shadowed_entropy_mode_update_err,
    cfg_shadowed_entropy_fast_process_update_err,
    cfg_shadowed_msg_mask_update_err,
    cfg_shadowed_entropy_ready_update_err,
    cfg_shadowed_err_processed_update_err,
    cfg_shadowed_en_unsupported_modestrength_update_err,
    entropy_refresh_threshold_shadowed_update_err
  };

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// KMAC control and padding logic

`include "prim_assert.sv"

module kmac_core
  import kmac_pkg::*;
#(
  // EnMasking: Enable masking security hardening inside keccak_round
  // If it is enabled, the result digest will be two set of 1600bit.
  parameter  bit EnMasking = 0,
  localparam int Share = (EnMasking) ? 2 : 1 // derived parameter
) (
  input clk_i,
  input rst_ni,

  // From Message FIFO
  input                fifo_valid_i,
  input [MsgWidth-1:0] fifo_data_i [Share],
  input [MsgStrbW-1:0] fifo_strb_i,
  output logic         fifo_ready_o,

  // to SHA3 Core
  output logic                msg_valid_o,
  output logic [MsgWidth-1:0] msg_data_o  [Share],
  output logic [MsgStrbW-1:0] msg_strb_o,
  input                       msg_ready_i,

  // Configurations

  // If kmac_en is cleared, Core logic doesn't function but forward incoming
  // message to SHA3 core
  input                             kmac_en_i,
  input sha3_pkg::sha3_mode_e       mode_i,
  input sha3_pkg::keccak_strength_e strength_i,

  // Key input from CSR
  input [MaxKeyLen-1:0] key_data_i [Share],
  input key_len_e       key_len_i,

  // Controls : same to SHA3 core
  input start_i,
  input process_i,
  input prim_mubi_pkg::mubi4_t done_i,

  // Control to SHA3 core
  output logic process_o,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  output logic sparse_fsm_error_o,
  output logic key_index_error_o
);

  import sha3_pkg::KeccakMsgAddrW;
  import sha3_pkg::KeccakCountW;
  import sha3_pkg::KeccakRate;
  import sha3_pkg::L128;
  import sha3_pkg::L224;
  import sha3_pkg::L256;
  import sha3_pkg::L384;
  import sha3_pkg::L512;

  /////////////////
  // Definitions //
  /////////////////

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 5 -n 6 \
  //      -s 401658243 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (50.00%)
  //  4: |||||||||||||||| (40.00%)
  //  5: |||| (10.00%)
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 5
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 4
  //
  localparam int StateWidth = 6;
  typedef enum logic [StateWidth-1:0] {
    StKmacIdle = 6'b011000,

    // Secret Key pushing stage
    // The key is sliced by prim_slicer. This state pushes the sliced data into
    // SHA3 hashing engine. When it hits the block size limit,
    // (same as in sha3pad) the state machine moves to Message.
    StKey = 6'b010111,

    // Incoming Message
    // The core does nothing but forwarding the incoming message to SHA3 hashing
    // engine by turning off `en_kmac_datapath`.
    StKmacMsg = 6'b001110,

    // Wait till done signal
    StKmacFlush = 6'b101011,

    // Terminal Error
    StTerminalError = 6'b100000
  } kmac_st_e ;

  /////////////
  // Signals //
  /////////////

  // represents encode_string(K)
  logic [MaxEncodedKeyW-1:0] encoded_key [Share];

  // Key slice address
  // This signal controls the 64 bit output of the sliced secret_key.
  logic [sha3_pkg::KeccakMsgAddrW-1:0] key_index;
  logic inc_keyidx, clr_keyidx;

  // `sent_blocksize` indicates that the encoded key is sent to sha3 hashing
  // engine. If this hits at StKey stage, the state moves to message state.
  logic [sha3_pkg::KeccakCountW-1:0] block_addr_limit;
  logic sent_blocksize;

  // Internal message signals
  logic                kmac_valid       ;
  logic [MsgWidth-1:0] kmac_data [Share];
  logic [MsgStrbW-1:0] kmac_strb        ;

  // Control SHA3 core
  // `kmac_process` is to forward the process signal to SHA3 core only after
  // the KMAC core writes the key block in case of the message is empty.
  // If the incoming message is empty, there's chance that the `process_i`
  // signal can be asserted while KMAC core processing the key block.
  logic kmac_process, process_latched;

  // Indication of Secret key write stage. Only in this stage, the internal
  // message interface is active.
  logic en_key_write;
  logic en_kmac_datapath;

  // Encoded key has wider bits. `key_sliced` is the data to send to sha3
  logic [MsgWidth-1:0] key_sliced [Share];

  sha3_pkg::sha3_mode_e unused_mode;
  assign unused_mode = mode_i;

  /////////
  // FSM //
  /////////
  kmac_st_e st, st_d;

  // State register
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, st_d, st, kmac_st_e, StKmacIdle)

  // Next state and output logic
  // SEC_CM: FSM.SPARSE
  always_comb begin
    st_d = st;

    en_kmac_datapath = 1'b 0;
    en_key_write = 1'b 0;

    clr_keyidx = 1'b 0;

    kmac_valid = 1'b 0;
    kmac_process = 1'b 0;

    sparse_fsm_error_o = 1'b 0;

    unique case (st)
      StKmacIdle: begin
        if (kmac_en_i && start_i) begin
          st_d = StKey;
        end else begin
          st_d = StKmacIdle;
        end
      end

      // If State enters here, regardless of the `process_i`, the state writes
      // full block size of the key into SHA3 hashing engine.
      StKey: begin
        en_kmac_datapath = 1'b 1;
        en_key_write = 1'b 1;

        if (sent_blocksize) begin
          st_d = StKmacMsg;

          kmac_valid = 1'b 0;
          clr_keyidx = 1'b 1;
        end else begin
          st_d = StKey;

          kmac_valid = 1'b 1;
        end
      end

      StKmacMsg: begin
        // If process is previously latched, it is sent to SHA3 here.
        if (process_i || process_latched) begin
          st_d = StKmacFlush;

          kmac_process = 1'b 1;
        end else begin
          st_d = StKmacMsg;
        end
      end

      StKmacFlush: begin
        if (prim_mubi_pkg::mubi4_test_true_strict(done_i)) begin
          st_d = StKmacIdle;
        end else begin
          st_d = StKmacFlush;
        end
      end

      StTerminalError: begin
        // this state is terminal
        st_d = st;
        sparse_fsm_error_o = 1'b 1;
      end

      default: begin
        // this state is terminal
        st_d = StTerminalError;
        sparse_fsm_error_o = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      st_d = StTerminalError;
    end
  end

  //////////////
  // Datapath //
  //////////////

  // DATA Mux depending on kmac_en
  // When Key write happens, hold the FIFO request. so fifo_ready_o is tied to 0
  assign msg_valid_o  = (en_kmac_datapath) ? kmac_valid : fifo_valid_i;
  assign msg_data_o   = (en_kmac_datapath) ? kmac_data  : fifo_data_i ;
  assign msg_strb_o   = (en_kmac_datapath) ? kmac_strb  : fifo_strb_i ;
  assign fifo_ready_o = (en_kmac_datapath) ? 1'b 0      : msg_ready_i ;

  // secret key write request to SHA3 hashing engine is always full width write.
  // KeyMgr is fixed 256 bit output. So `right_encode(256)` is 0x020100 --> strb 3
  assign kmac_strb = (en_key_write ) ? '1 : '0;

  assign kmac_data = (en_key_write) ? key_sliced : '{default:'0};

  // Process is controlled by the KMAC core always.
  // This is mainly to prevent process_i asserted while KMAC core is writing
  // the secret key to SHA3 hashing engine (the empty message case)
  assign process_o = (kmac_en_i) ? kmac_process : process_i ;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      process_latched <= 1'b 0;
    end else if (process_i && !process_o) begin
      process_latched <= 1'b 1;
    end else if (process_o ||
      prim_mubi_pkg::mubi4_test_true_strict(done_i)) begin
      process_latched <= 1'b 0;
    end
  end

  // bytepad(encode_string(K), 168 or 136) =====================================
  // 1. Prepare left_encode(w)
  // 2. Prepare left_encode(len(secret_key))
  // 3. Concatenate left_encode(len(secret_key)) || secret_key
  // 4. Concaatenate left_encode(w) || encode_string(secret_key)
  // 5. Based on the address, slice out the data into MsgWidth bits

  // left_encode(w): Same as used in sha3pad logic.
  logic [15:0] encode_bytepad;
  assign encode_bytepad = sha3_pkg::encode_bytepad_len(strength_i);

  // left_encode(len(secret_key))
  // encoded length is always byte size. Use MaxEncodedKeyLenByte parameter
  // from kmac_pkg and add one more byte to indicate how many bytes used to
  // represent len(secret_key)
  // Note that if the secret_key is 128 bit, only lower 16 bits of
  // `encode_keylen` are valid. Refer `encoded_key` concatenation logic below.
  // As the encoded string in the spec big-endian, The endian swap is a must.
  logic [MaxEncodedKeyLenSize + 8 - 1:0] encode_keylen [Share];

  always_comb begin
    // the spec mentioned the key length is encoded in left_encode()
    // The number is represented in big-endian. For example:
    // 384 ==> 0x02 0x01 0x80
    // The first byte is the number of bytes to represent 384
    // The second byte represents 2**8 number, which is 256 here.
    // The third byte represents 2**0 number, which is 128.
    // The data put into MsgFIFO is little-endian and SHA3(Keccak) processes in
    // little-endian. So, below keylen swaps the byte order
    unique case (key_len_i)
      //                           endian-swapped key_length          num_bytes
      // Key128: encode_keylen[0] = {{<<8{MaxEncodedKeyLenSize'(128)}}, 8'h 01};
      // Key192: encode_keylen[0] = {{<<8{MaxEncodedKeyLenSize'(192)}}, 8'h 01};
      // Key256: encode_keylen[0] = {{<<8{MaxEncodedKeyLenSize'(256)}}, 8'h 02};
      // Key384: encode_keylen[0] = {{<<8{MaxEncodedKeyLenSize'(384)}}, 8'h 02};
      // Key512: encode_keylen[0] = {{<<8{MaxEncodedKeyLenSize'(512)}}, 8'h 02};

      // Vivado does not support stream swap for non context value. So assign
      // the value directly.
      Key128: encode_keylen[0] = (MaxEncodedKeyLenSize+8)'('h 0080_01);
      Key192: encode_keylen[0] = (MaxEncodedKeyLenSize+8)'('h 00C0_01);
      Key256: encode_keylen[0] = (MaxEncodedKeyLenSize+8)'('h 0001_02);
      Key384: encode_keylen[0] = (MaxEncodedKeyLenSize+8)'('h 8001_02);
      Key512: encode_keylen[0] = (MaxEncodedKeyLenSize+8)'('h 0002_02);
      default: encode_keylen[0] = '0;
    endcase
  end

  if (EnMasking) begin: gen_encode_keylen_masked
    assign encode_keylen[1] = '0;
  end

  // encode_string(secret_key): Concatenate key
  // Based on the left_encode(len(secret_key)) size, the concatenation logic
  // should be changed. If key length is 128 bit, only lower 16 bits of the
  // encoded length are used so that the upper 8 bits are padded with 0 as
  // defined in bytepad() function.

  for (genvar i = 0 ; i < Share; i++) begin : gen_encoded_key
    always_comb begin
      unique case (key_len_i)
        // In Key 128, 192 case, only lower parts of encode_keylen signal is
        // used. So upper padding requires 8 more bits than MaxKeyLen - keylen
        Key128: encoded_key[i] = {(8 + MaxKeyLen - 128)'(0),
                                  key_data_i[i][0+:128],
                                  encode_keylen[i][0+:MaxEncodedKeyLenSize]};

        Key192: encoded_key[i] = {(8 + MaxKeyLen - 192)'(0),
                                  key_data_i[i][0+:192],
                                  encode_keylen[i][0+:MaxEncodedKeyLenSize]};

        Key256: encoded_key[i] = {(MaxKeyLen - 256)'(0),
                                  key_data_i[i][0+:256],
                                  encode_keylen[i]};

        Key384: encoded_key[i] = {(MaxKeyLen - 384)'(0),
                                  key_data_i[i][0+:384],
                                  encode_keylen[i]};

        // Assume 512bit is the MaxKeyLen
        Key512: encoded_key[i] = {key_data_i[i][0+:512],
                                  encode_keylen[i]};

        default: encoded_key[i] = '0;
      endcase
    end
  end : gen_encoded_key

  // Above logic assumes MaxKeyLen as 512 bits. Revise if it is not.
  `ASSERT_INIT(MaxKeyLenMatchToKey512_A, kmac_pkg::MaxKeyLen == 512)

  // Combine the bytepad `left_encode(w)` and the `encode_string(secret_key)`
  logic [MaxEncodedKeyW + 16 -1 :0] encoded_key_block [Share];

  assign encoded_key_block[0] = {encoded_key[0], encode_bytepad};

  if (EnMasking) begin : gen_encoded_key_block_masked
    assign encoded_key_block[1] = {encoded_key[1], 16'h 0};
  end

  // Slicer to slice out 64 bits
  for (genvar i = 0 ; i < Share ; i++) begin : gen_key_slicer
    prim_slicer #(
      .InW (MaxEncodedKeyW+16),
      .IndexW(KeccakMsgAddrW),
      .OutW(MsgWidth)
    ) u_key_slicer (
      .sel_i  (key_index),
      .data_i (encoded_key_block[i]),
      .data_o (key_sliced[i])
    );
  end

  // `key_index` logic
  // key_index is used to select MsgWidth data from long `encoded_key_block`
  // It behaves same as `keccak_addr` or `prefix_index` in sha3pad module.
  assign inc_keyidx = kmac_valid & msg_ready_i ;

  // This primitive is used to place a hardened counter
  // SEC_CM: CTR.REDUN
  prim_count #(
    .Width(sha3_pkg::KeccakMsgAddrW)
  ) u_key_index_count (
    .clk_i,
    .rst_ni,
    .clr_i(clr_keyidx),
    .set_i(1'b0),
    .set_cnt_i('0),
    .incr_en_i(inc_keyidx),
    .decr_en_i(1'b0),
    .step_i(sha3_pkg::KeccakMsgAddrW'(1)),
    .cnt_o(key_index),
    .cnt_next_o(),
    .err_o(key_index_error_o)
  );

  // Block size based on the address.
  // This is used for bytepad() and also pad10*1()
  // assign block_addr_limit = KeccakRate[strength_i];
  // but below is easier to understand
  always_comb begin
    unique case (strength_i)
      L128: block_addr_limit = KeccakCountW'(KeccakRate[L128]);
      L224: block_addr_limit = KeccakCountW'(KeccakRate[L224]);
      L256: block_addr_limit = KeccakCountW'(KeccakRate[L256]);
      L384: block_addr_limit = KeccakCountW'(KeccakRate[L384]);
      L512: block_addr_limit = KeccakCountW'(KeccakRate[L512]);

      default: block_addr_limit = '0;
    endcase
  end

  assign sent_blocksize = (key_index == block_addr_limit);


  // Encoded Output Length =====================================================
  //
  // KMAC(K,X,L,S) := cSHAKE(newX,L,"KMAC",S)
  //   K : Secret Key
  //   X : Input Message
  //   L : Output Length
  //   S : Customization input string
  //   newX = bytepad(encode_string(key), 168or136) || X || right_encode(L)
  //
  // Software writes desired output length as encoded value into the message
  // FIFO at the end of the message prior to set !!CMD.process.


  ////////////////
  // Assertions //
  ////////////////

  // If process_latched is set, then at Message state, it should be cleared

  `ASSERT(ProcessLatchedCleared_A,
          st == StKmacMsg && process_latched |=> !process_latched)

  // Assume configuration is stable during the operation
  `ASSUME(KmacEnStable_M, $changed(kmac_en_i) |-> st inside {StKmacIdle, StTerminalError})
  `ASSUME(ModeStable_M, $changed(mode_i) |-> st inside {StKmacIdle, StTerminalError})
  `ASSUME(StrengthStable_M,
          $changed(strength_i) |->
          (st inside {StKmacIdle, StTerminalError}) ||
          ($past(st) == StKmacIdle))
  `ASSUME(KeyLengthStable_M,
          $changed(key_len_i) |->
          (st inside {StKmacIdle, StTerminalError}) ||
          ($past(st) == StKmacIdle))
  `ASSUME(KeyDataStable_M,
          $changed(key_data_i) |->
          (st inside {StKmacIdle, StTerminalError}) ||
          ($past(st) == StKmacIdle))

  // no acked to MsgFIFO in StKmacMsg
  `ASSERT(AckOnlyInMessageState_A,
          fifo_valid_i && fifo_ready_o && kmac_en_i |-> st == StKmacMsg)

endmodule : kmac_core


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// KMAC MSG_FIFO
//
// This module converts TL-UL interface into MSG_FIFO interface used in KMAC.

`include "prim_assert.sv"

module kmac_msgfifo
  import kmac_pkg::*;
#(
  // OutWidth is MsgFIFO data width. prim_packer converts InW to OutW prior to
  // pushing to MsgFIFO
  parameter int OutWidth = 64,

  parameter bit EnMasking = 1'b 1,

  // Internal MsgFIFO Entry count
  parameter  int MsgDepth = 9,
  localparam int MsgDepthW = $clog2(MsgDepth+1) // derived parameter
) (
  input clk_i,
  input rst_ni,

  // from REG or KeyMgr Intf input
  input                fifo_valid_i,
  input [OutWidth-1:0] fifo_data_i,
  input [OutWidth-1:0] fifo_mask_i,
  output               fifo_ready_o,

  // MSG interface
  output logic                  msg_valid_o,
  output logic [OutWidth-1:0]   msg_data_o,
  output logic [OutWidth/8-1:0] msg_strb_o,
  input                         msg_ready_i,

  output logic                 fifo_empty_o,
  output logic                 fifo_full_o,
  output logic [MsgDepthW-1:0] fifo_depth_o,

  // Control
  input prim_mubi_pkg::mubi4_t clear_i,

  // process_i --> process_o
  // process_o asserted after all internal messages are flushed out to MSG interface
  input        process_i,
  output logic process_o,

  err_t err_o
);

  /////////////////
  // Definitions //
  /////////////////
  typedef struct packed {
    logic [OutWidth-1:0]   data;
    logic [OutWidth/8-1:0] strb; // one bit per byte
  } fifo_t;

  typedef enum logic [1:0] {
    // In Idle, it checks if process input received or not.
    // If received, the signal goes to packer and flush internal pending data
    FlushIdle,

    // In Packer state, it waits the packer flush operation completes.
    // The flush_done signal do nothing but after this, it is assumed that
    // MSG FIFO received the request.
    FlushPacker,

    // In Fifo, it waits until MsgFifo is empty. Then asserts process_o
    FlushFifo,

    // After flushing, it waits the done (clear) signal. It is assumed that
    // no incoming messages are transmitted between `process_i` and `clear_i`
    FlushClear
  } flush_st_e;

  /////////////
  // Signals //
  /////////////

  // Packer write path
  logic                packer_wvalid;
  logic [OutWidth-1:0] packer_wdata;
  logic [OutWidth-1:0] packer_wmask;
  logic                packer_wready;

  // Message FIFO signals
  logic  fifo_wvalid;
  fifo_t fifo_wdata;
  logic  fifo_wready;
  logic  fifo_rvalid;
  fifo_t fifo_rdata;
  logic  fifo_rready;

  logic fifo_err; // FIFO dup. counter error

  // packer flush to msg_fifo, then msg_fifo empty out the internals
  // then assert msgfifo_flush_done
  logic packer_flush_done;
  logic msgfifo_flush_done;

  logic packer_err;

  // SEC_CM: PACKER.CTR.REDUN
  prim_packer #(
    .InW          (OutWidth),
    .OutW         (OutWidth),
    .HintByteData (1),

    // Turn on dup counter when EnMasking is set
    .EnProtection (EnMasking)
  ) u_packer (
    .clk_i,
    .rst_ni,

    .valid_i      (fifo_valid_i),
    .data_i       (fifo_data_i),
    .mask_i       (fifo_mask_i),
    .ready_o      (fifo_ready_o),

    .valid_o      (packer_wvalid),
    .data_o       (packer_wdata),
    .mask_o       (packer_wmask),
    .ready_i      (packer_wready),

    .flush_i      (process_i),
    .flush_done_o (packer_flush_done),

    .err_o (packer_err)
  );

  // Assign packer wdata and wmask to FIFO struct
  // In contrast to HMAC case, KMAC SHA3 operates in little-endian. MSG fifo is
  // converted into 3-D form so the endianess here is not a problem.
  assign fifo_wdata.data = packer_wdata;
  always_comb begin
    fifo_wdata.strb = '0;
    for (int i = 0 ; i < OutWidth/8 ; i++) begin
      fifo_wdata.strb[i] = packer_wmask[8*i];
    end
  end

  // MsgFIFO
  prim_fifo_sync #(
    .Width  ($bits(fifo_t)),
    .Pass   (1'b 1),
    .Depth  (MsgDepth),
    .Secure (EnMasking)
  ) u_msgfifo (
    .clk_i,
    .rst_ni,
    .clr_i   (prim_mubi_pkg::mubi4_test_true_strict(clear_i)),

    .wvalid_i(fifo_wvalid),
    .wready_o(fifo_wready),
    .wdata_i (fifo_wdata),

    .rvalid_o (fifo_rvalid),
    .rready_i (fifo_rready),
    .rdata_o  (fifo_rdata),

    .full_o  (fifo_full_o),
    .depth_o (fifo_depth_o),
    .err_o   (fifo_err)

  );

  assign fifo_wvalid = packer_wvalid;
  assign packer_wready = fifo_wready;

  assign msg_valid_o = fifo_rvalid;
  assign fifo_rready = msg_ready_i;
  assign msg_data_o  = fifo_rdata.data;
  assign msg_strb_o  = fifo_rdata.strb;

  assign fifo_empty_o = !fifo_rvalid;

  // Flush (process from outside) handling
  flush_st_e flush_st, flush_st_d;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      flush_st <= FlushIdle;
    end else begin
      flush_st <= flush_st_d;
    end
  end

  always_comb begin
    flush_st_d = flush_st;

    msgfifo_flush_done = 1'b 0;

    unique case (flush_st)
      FlushIdle: begin
        if (process_i) begin
          flush_st_d = FlushPacker;
        end else begin
          flush_st_d = FlushIdle;
        end
      end

      FlushPacker: begin
        if (packer_flush_done) begin
          flush_st_d = FlushFifo;
        end else begin
          flush_st_d = FlushPacker;
        end
      end

      FlushFifo: begin
        if (fifo_empty_o) begin
          flush_st_d = FlushClear;

          msgfifo_flush_done = 1'b 1;
        end else begin
          flush_st_d = FlushFifo;
        end
      end

      FlushClear: begin
        if (prim_mubi_pkg::mubi4_test_true_strict(clear_i)) begin
          flush_st_d = FlushIdle;
        end else begin
          flush_st_d = FlushClear;
        end
      end

      default: begin
        flush_st_d = FlushIdle;
      end
    endcase
  end

  assign process_o = msgfifo_flush_done;

  // Error assign
  always_comb begin : error_logic
    err_o = '{
      valid: 1'b 0,
      code: kmac_pkg::ErrNone,
      info: '0
    };

    // Priority case -> if .. else if
    if (packer_err) begin
      err_o = '{
        // If EnProtection is 0, packer_err is tied to 0
        valid: 1'b 1,
        code:  kmac_pkg::ErrPackerIntegrity,
        info:  kmac_pkg::ErrInfoW'(flush_st)
      };
    end else if (fifo_err) begin
      err_o = '{
        valid: 1'b 1,
        code:  kmac_pkg::ErrMsgFifoIntegrity,
        info:  kmac_pkg::ErrInfoW'(flush_st)
      };
    end
  end : error_logic

  ////////////////
  // Assertions //
  ////////////////

  // Flush state known checker
  `ASSERT(FlushStInValid_A, flush_st inside {FlushIdle, FlushPacker, FlushFifo, FlushClear})

  // Packer done signal is asserted at least one cycle later
  `ASSERT(PackerDoneDelay_A, $onehot0({process_i, packer_flush_done}))

  // process_i not asserted during the flush operation
  `ASSUME(PackerDoneValid_a, process_i |-> flush_st == FlushIdle)

  // No messages in between `process_i` and `clear_i`
  `ASSUME(MessageValid_a, fifo_valid_i |-> flush_st == FlushIdle)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Keccak state read

`include "prim_assert.sv"

module kmac_staterd
  import kmac_pkg::*;
#(
  // TL-UL Address Width. Should be bigger than
  // $clog2(kmac_pkg::StateW) * Share
  parameter int AddrW = 9,

  // EnMasking: Enable masking security hardening inside keccak_round
  // If it is enabled, the result digest will be two set of 1600bit.
  parameter  bit EnMasking = 1'b0,
  localparam int Share = (EnMasking) ? 2 : 1  // derived parameter
) (
  input clk_i,
  input rst_ni,

  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // State in
  input [sha3_pkg::StateW-1:0] state_i [Share],

  // Config
  input endian_swap_i
);

  localparam int StateAddrW = $clog2(sha3_pkg::StateW/32);
  localparam int SelAddrW   = AddrW-2-StateAddrW;

  /////////////
  // Signals //
  /////////////

  // TL-UL Adapter signals
  logic             tlram_req;
  logic             tlram_gnt;
  logic             tlram_we;
  logic [AddrW-3:0] tlram_addr;   // Word base
  logic [31:0]      unused_tlram_wdata;
  logic [31:0]      unused_tlram_wmask;
  logic [31:0]      tlram_rdata;
  logic             tlram_rvalid;
  logic [1:0]       tlram_rerror;
  logic [31:0]      tlram_rdata_endian;

  // TL Adapter
  tlul_adapter_sram #(
    .SramAw (AddrW-2),
    .SramDw (32),
    .Outstanding (1),
    .ByteAccess  (1),
    .ErrOnWrite  (1),
    .ErrOnRead   (0)
  ) u_tlul_adapter (
    .clk_i,
    .rst_ni,

    .tl_i,
    .tl_o,
    .en_ifetch_i (prim_mubi_pkg::MuBi4False),
    .req_o       (tlram_req),
    .req_type_o  (),
    .gnt_i       (tlram_gnt),
    .we_o        (tlram_we ),
    .addr_o      (tlram_addr),
    .wdata_o     (unused_tlram_wdata),
    .wmask_o     (unused_tlram_wmask),
    .intg_error_o(),
    .rdata_i     (tlram_rdata),
    .rvalid_i    (tlram_rvalid),
    .rerror_i    (tlram_rerror)
  );

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      tlram_rdata <= '0;
    end else if (tlram_req & ~tlram_we) begin
      tlram_rdata <= conv_endian32(tlram_rdata_endian, endian_swap_i);
    end
  end

  // Always grant
  assign tlram_gnt = tlram_req & ~tlram_we;

  // always no error on reading
  assign tlram_rerror = '0;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) tlram_rvalid <= 1'b0;
    else         tlram_rvalid <= tlram_req & !tlram_we;
  end

  logic [31:0] muxed_state [Share];


  for (genvar i = 0 ; i < Share ; i++) begin : gen_slicer
    prim_slicer #(
      .InW (sha3_pkg::StateW),
      .OutW (32),
      .IndexW (StateAddrW)
    ) u_state_slice (
      .sel_i (tlram_addr[StateAddrW-1:0]),
      .data_i (state_i[i]),
      .data_o (muxed_state[i])
    );
  end : gen_slicer

  logic [SelAddrW-1:0] addr_sel;
  assign addr_sel = tlram_addr[StateAddrW+:SelAddrW];

  assign tlram_rdata_endian = int'(addr_sel) < Share ? muxed_state[addr_sel] : 0;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// KMAC Application interface

`include "prim_assert.sv"

module kmac_app
  import kmac_pkg::*;
#(
  // App specific configs are defined in kmac_pkg
  parameter  bit EnMasking = 1'b0,
  localparam int Share = (EnMasking) ? 2 : 1, // derived parameter
  parameter  bit SecIdleAcceptSwMsg = 1'b0
) (
  input clk_i,
  input rst_ni,

  // Secret Key from register
  input [MaxKeyLen-1:0] reg_key_data_i [Share],
  input key_len_e       reg_key_len_i,

  // Prefix from register
  input [sha3_pkg::NSRegisterSize*8-1:0] reg_prefix_i,

  // mode, strength, kmac_en from register
  input                             reg_kmac_en_i,
  input sha3_pkg::sha3_mode_e       reg_sha3_mode_i,
  input sha3_pkg::keccak_strength_e reg_keccak_strength_i,

  // Data from Software
  input                sw_valid_i,
  input [MsgWidth-1:0] sw_data_i,
  input [MsgWidth-1:0] sw_mask_i,
  output logic         sw_ready_o,

  // KeyMgr Sideload Key interface
  input keymgr_pkg::hw_key_req_t keymgr_key_i,

  // Application Message in/ Digest out interface + control signals
  input  app_req_t [NumAppIntf-1:0] app_i,
  output app_rsp_t [NumAppIntf-1:0] app_o,

  // to KMAC Core: Secret key
  output logic [MaxKeyLen-1:0] key_data_o [Share],
  output key_len_e             key_len_o,

  // to MSG_FIFO
  output logic                kmac_valid_o,
  output logic [MsgWidth-1:0] kmac_data_o,
  output logic [MsgWidth-1:0] kmac_mask_o,
  input                       kmac_ready_i,

  // KMAC Core
  output logic kmac_en_o,

  // To Sha3 Core
  output logic [sha3_pkg::NSRegisterSize*8-1:0] sha3_prefix_o,
  output sha3_pkg::sha3_mode_e                  sha3_mode_o,
  output sha3_pkg::keccak_strength_e            keccak_strength_o,

  // STATE from SHA3 Core
  input                        keccak_state_valid_i,
  input [sha3_pkg::StateW-1:0] keccak_state_i [Share],

  // to STATE TL-window if Application is not active, the incoming state goes to
  // register if kdf_en is set, the state value goes to application and the
  // output to the register is all zero.
  output logic                        reg_state_valid_o,
  output logic [sha3_pkg::StateW-1:0] reg_state_o [Share],

  // Configurations If key_en is set, the logic uses KeyMgr's sideloaded key as
  // a secret key rather than register values. This only affects when software
  // initiates. If App initiates the hash operation and uses KMAC algorithm, it
  // always uses sideloaded key.
  input keymgr_key_en_i,

  // Commands
  // Command from software
  input kmac_cmd_e sw_cmd_i,

  // from SHA3
  input prim_mubi_pkg::mubi4_t absorbed_i,

  // to KMAC
  output kmac_cmd_e cmd_o,

  // to SW
  output prim_mubi_pkg::mubi4_t absorbed_o,

  // To status
  output logic app_active_o,

  // Status
  // - entropy_ready_i: Entropy configured by SW. It is used to check if App
  //                    is OK to request.
  input prim_mubi_pkg::mubi4_t entropy_ready_i,

  // Error input
  // This error comes from KMAC/SHA3 engine.
  // KeyMgr interface delivers the error signal to KeyMgr to drop the current op
  // and re-initiate.
  // If error happens, regardless of SW-initiated or KeyMgr-initiated, the error
  // is reported to the ERR_CODE so that SW can look into.
  input error_i,

  // SW sets err_processed bit in CTRL then the logic goes to Idle
  input err_processed_i,

  // error_o value is pushed to Error FIFO at KMAC/SHA3 top and reported to SW
  output kmac_pkg::err_t error_o,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  output logic sparse_fsm_error_o
);

  import sha3_pkg::KeccakBitCapacity;
  import sha3_pkg::L128;
  import sha3_pkg::L224;
  import sha3_pkg::L256;
  import sha3_pkg::L384;
  import sha3_pkg::L512;

  /////////////////
  // Definitions //
  /////////////////

  // Digest width is same to the key width `keymgr_pkg::KeyWidth`.
  localparam int KeyMgrKeyW = $bits(keymgr_key_i.key[0]);

  localparam key_len_e KeyLengths [5] = '{Key128, Key192, Key256, Key384, Key512};

  localparam int SelKeySize = (AppKeyW == 128) ? 0 :
                              (AppKeyW == 192) ? 1 :
                              (AppKeyW == 256) ? 2 :
                              (AppKeyW == 384) ? 3 :
                              (AppKeyW == 512) ? 4 : 0 ;
  localparam int SelDigSize = (AppDigestW == 128) ? 0 :
                              (AppDigestW == 192) ? 1 :
                              (AppDigestW == 256) ? 2 :
                              (AppDigestW == 384) ? 3 :
                              (AppDigestW == 512) ? 4 : 0 ;
  localparam key_len_e SideloadedKey = KeyLengths[SelKeySize];

  // Define right_encode(outlen) value here
  // Look at kmac_pkg::key_len_e for the kinds of key size
  //
  // These values should be exactly the same as the key length encodings
  // in kmac_core.sv, with the only difference being that the byte representing
  // the byte-length of the encoded value is in the MSB position due to right encoding
  // instead of in the LSB position (left encoding).
  localparam int OutLenW = 24;
  localparam logic [OutLenW-1:0] EncodedOutLen [5]= '{
    24'h 0001_80, // Key128
    24'h 0001_C0, // Key192
    24'h 02_0001, // Key256
    24'h 02_8001, // Key384
    24'h 02_0002  // Key512
  };

  localparam logic [OutLenW-1:0] EncodedOutLenMask [5] = '{
    24'h 00FFFF, // Key128,
    24'h 00FFFF, // Key192
    24'h FFFFFF, // Key256
    24'h FFFFFF, // Key384
    24'h FFFFFF  // Key512
  };

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 11 -n 10 \
  //      -s 155490773 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: ||||||||||||| (14.55%)
  //  4: |||||||||||||||||||| (21.82%)
  //  5: |||||||||||||||||| (20.00%)
  //  6: |||||||||||||||||||| (21.82%)
  //  7: |||||||||||||||||| (20.00%)
  //  8: | (1.82%)
  //  9: --
  // 10: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 8
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 9
  //
  localparam int StateWidth = 10;
  // States
  //  StIdle                  = 10'b0101110011,
  //  StAppCfg                = 10'b0001010000,
  //  StAppMsg                = 10'b0001011111,
  //  StAppOutLen             = 10'b1011001111,
  //  StAppProcess            = 10'b1000100110,
  //  StAppWait               = 10'b0010010110,
  //  StSw                    = 10'b0111111111,
  //  StKeyMgrErrKeyNotValid  = 10'b1001110100,
  //  StError                 = 10'b1101011101,
  //  StServiceRejectedError  = 10'b1110000110,
  //  StTerminalError         = 10'b0010001001
  typedef enum logic [StateWidth-1:0] {
    StIdle = 10'b0101110011,

    // Application operation.
    //
    // if start request comes from an App first, until the operation ends by the
    // requested App, all operations are granted to the specific App. SW
    // requests and other Apps requests will be ignored.
    //
    // App interface does not have control signals. When first data valid occurs
    // from an App, this logic asserts the start command to the downstream. When
    // last beat pulse comes, this logic asserts the process to downstream
    // (after the transaction is accepted regardless of partial writes or not)
    // When absorbed by SHA3 core, the logic sends digest to the requested App
    // and right next cycle, it triggers done command to downstream.

    // In StAppCfg state, it latches the cfg from AppCfg parameter to determine
    // the kmac_mode, sha3_mode, keccak strength.
    StAppCfg = 10'b0001010000,

    StAppMsg = 10'b0001011111,

    // In StKeyOutLen, this module pushes encoded outlen to the MSG_FIFO.
    // Assume the length is 256 bit, the data will be 48'h 02_0100
    StAppOutLen  = 10'b1011001111,
    StAppProcess = 10'b1000100110,
    StAppWait    = 10'b0010010110,

    // SW Controlled
    // If start request comes from SW first, until the operation ends, all
    // requests from KeyMgr will be discarded.
    StSw = 10'b0111111111,

    // Error KeyNotValid
    // When KeyMgr operates, the secret key is not ready yet.
    StKeyMgrErrKeyNotValid = 10'b1001110100,

    StError = 10'b1101011101,

    StServiceRejectedError = 10'b1110000110,

    // This state is used for terminal errors
    StTerminalError = 10'b0010001001
  } st_e;

  /////////////
  // Signals //
  /////////////

  st_e st, st_d;

  // app_rsp_t signals
  // The state machine controls mux selection, which controls the ready signal
  // the other responses are controled in separate logic. So define the signals
  // here and merge them to the response.
  logic app_data_ready, fsm_data_ready;
  logic app_digest_done, fsm_digest_done_q, fsm_digest_done_d;
  logic [AppDigestW-1:0] app_digest [2];

  // One more slot for value NumAppIntf. It is the value when no app intf is
  // chosen.
  localparam int unsigned AppIdxW = $clog2(NumAppIntf);

  // app_id indicates, which app interface was chosen. various logic use this
  // value to get the config or return the data.
  logic [AppIdxW-1:0] app_id, app_id_d;
  logic               clr_appid, set_appid;

  // Output length
  logic [OutLenW-1:0] encoded_outlen, encoded_outlen_mask;

  // state output
  // Mux selection signal
  app_mux_sel_e mux_sel;
  app_mux_sel_e mux_sel_buf_output;
  app_mux_sel_e mux_sel_buf_err_check;
  app_mux_sel_e mux_sel_buf_kmac;

  // Error checking logic

  kmac_pkg::err_t fsm_err, mux_err;

  logic service_rejected_error;
  logic service_rejected_error_set, service_rejected_error_clr;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)                         service_rejected_error <= 1'b 0;
    else if (service_rejected_error_set) service_rejected_error <= 1'b 1;
    else if (service_rejected_error_clr) service_rejected_error <= 1'b 0;
  end

  ////////////////////////////
  // Application Mux/ Demux //
  ////////////////////////////


  // Processing return data.
  // sends to only selected app intf.
  // clear digest right after done to not leak info to other interface
  always_comb begin
    for (int unsigned i = 0 ; i < NumAppIntf ; i++) begin
      if (i == app_id) begin
        app_o[i] = '{
          ready:         app_data_ready | fsm_data_ready,
          done:          app_digest_done | fsm_digest_done_q,
          digest_share0: app_digest[0],
          digest_share1: app_digest[1],
          // if fsm asserts done, should be an error case.
          error:         error_i | fsm_digest_done_q | sparse_fsm_error_o
                         | service_rejected_error
        };
      end else begin
        app_o[i] = '{
          ready: 1'b 0,
          done:  1'b 0,
          digest_share0: '0,
          digest_share1: '0,
          error: 1'b 0
        };
      end
    end // for {i, NumAppIntf, i++}
  end // aiways_comb

  // app_id latch
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) app_id <= AppIdxW'(0) ; // Do not select any
    else if (clr_appid) app_id <= AppIdxW'(0);
    else if (set_appid) app_id <= app_id_d;
  end

  // app_id selection as of now, app_id uses Priority. The assumption is that
  //  the request normally does not collide. (ROM_CTRL activates very early
  //  stage at the boot sequence)
  //
  //  If this assumption is not true, consider RR arbiter.

  // Prep for arbiter
  logic [NumAppIntf-1:0] app_reqs;
  logic [NumAppIntf-1:0] unused_app_gnts;
  logic [$clog2(NumAppIntf)-1:0] arb_idx;
  logic arb_valid;
  logic arb_ready;

  always_comb begin
    app_reqs = '0;
    for (int unsigned i = 0 ; i < NumAppIntf ; i++) begin
      app_reqs[i] = app_i[i].valid;
    end
  end

  prim_arbiter_fixed #(
    .N (NumAppIntf),
    .DW(1),
    .EnDataPort(1'b 0)
  ) u_appid_arb (
    .clk_i,
    .rst_ni,

    .req_i  (app_reqs),
    .data_i ('{default:'0}),
    .gnt_o  (unused_app_gnts),
    .idx_o  (arb_idx),

    .valid_o (arb_valid),
    .data_o  (), // not used
    .ready_i (arb_ready)
  );

  assign app_id_d = AppIdxW'(arb_idx);
  assign arb_ready = set_appid;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) fsm_digest_done_q <= 1'b 0;
    else         fsm_digest_done_q <= fsm_digest_done_d;
  end

  /////////
  // FSM //
  /////////

  // State register
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, st_d, st, st_e, StIdle)

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(KmacSecIdleAcceptSwMsgNonDefault, SecIdleAcceptSwMsg == 0)

  // Next State & output logic
  // SEC_CM: FSM.SPARSE
  always_comb begin
    st_d = st;

    mux_sel = SecIdleAcceptSwMsg ? SelSw : SelNone;

    // app_id control
    set_appid = 1'b 0;
    clr_appid = 1'b 0;

    // Commands
    cmd_o = CmdNone;

    // Software output
    absorbed_o = prim_mubi_pkg::MuBi4False;

    // Error
    fsm_err = '{valid: 1'b 0, code: ErrNone, info: '0};
    sparse_fsm_error_o = 1'b 0;

    service_rejected_error_set = 1'b 0;
    service_rejected_error_clr = 1'b 0;

    // If error happens, FSM asserts data ready but discard incoming msg
    fsm_data_ready = 1'b 0;
    fsm_digest_done_d = 1'b 0;

    unique case (st)
      StIdle: begin
        if (arb_valid) begin
          st_d = StAppCfg;

          // choose app_id
          set_appid = 1'b 1;
        end else if (sw_cmd_i == CmdStart) begin
          st_d = StSw;
          // Software initiates the sequence
          cmd_o = CmdStart;
        end else begin
          st_d = StIdle;
        end
      end

      StAppCfg: begin
        if (AppCfg[app_id].Mode == AppKMAC &&
          prim_mubi_pkg::mubi4_test_false_strict(entropy_ready_i)) begin
          // Check if the entropy is not configured but it is needed in
          // `AppCfg[app_id]` (KMAC mode).
          //
          // SW is not properly configured, report and not request Hashing
          // Return the app with errors
          st_d = StError;

          service_rejected_error_set = 1'b 1;

        end else if ((AppCfg[app_id].Mode == AppKMAC) &&
          !keymgr_key_i.valid) begin
          st_d = StKeyMgrErrKeyNotValid;

          // As mux_sel is not set to SelApp, app_data_ready is still 0.
          // This logic won't accept the requests from the selected App.

        end else begin
          // As Cfg is stable now, it sends cmd
          st_d = StAppMsg;

          // App initiates the data
          cmd_o = CmdStart;
        end
      end

      StAppMsg: begin
        mux_sel = SelApp;
        if (app_i[app_id].valid && app_o[app_id].ready && app_i[app_id].last) begin
          if (AppCfg[app_id].Mode == AppKMAC) begin
            st_d = StAppOutLen;
          end else begin
            st_d = StAppProcess;
          end
        end else begin
          st_d = StAppMsg;
        end
      end

      StAppOutLen: begin
        mux_sel = SelOutLen;

        if (kmac_valid_o && kmac_ready_i) begin
          st_d = StAppProcess;
        end else begin
          st_d = StAppOutLen;
        end
      end

      StAppProcess: begin
        cmd_o = CmdProcess;
        st_d = StAppWait;
      end

      StAppWait: begin
        if (prim_mubi_pkg::mubi4_test_true_strict(absorbed_i)) begin
          // Send digest to KeyMgr and complete the op
          st_d = StIdle;
          cmd_o = CmdDone;

          clr_appid = 1'b 1;
        end else begin
          st_d = StAppWait;
        end
      end

      StSw: begin
        mux_sel = SelSw;

        cmd_o = sw_cmd_i;
        absorbed_o = absorbed_i;

        if (sw_cmd_i == CmdDone) begin
          st_d = StIdle;
        end else begin
          st_d = StSw;
        end
      end

      StKeyMgrErrKeyNotValid: begin
        st_d = StError;

        // As mux_sel is not set to SelApp, app_data_ready is still 0.
        // This logic won't accept the requests from the selected App.
        fsm_err.valid = 1'b 1;
        fsm_err.code = ErrKeyNotValid;
        fsm_err.info = 24'(app_id);
      end

      StError: begin
        // In this state, the state machine flush out the request
        st_d = StError;

        fsm_data_ready = 1'b 1;

        if (err_processed_i) begin
          st_d = StIdle;

          // clear internal variables
          clr_appid = 1'b 1;
        end

        if (app_i[app_id].valid && app_i[app_id].last) begin
          // Send garbage digest to the app interface to complete transaction
          fsm_digest_done_d = 1'b 1;

          if (service_rejected_error) begin
            // If service was rejected, it is assumed the SW is not loaded
            // yet. In this case, return the request with error and keep
            // moving, hoping SW may handle the errors later
            st_d = StServiceRejectedError;
          end
        end

      end

      StServiceRejectedError: begin
        // Clear the error and move to Idle
        // At this state, the app responses the request with an error.
        st_d = StIdle;

        clr_appid = 1'b 1;
        service_rejected_error_clr = 1'b 1;
      end

      StTerminalError: begin
        // this state is terminal
        st_d = st;
        sparse_fsm_error_o = 1'b 1;
        fsm_err.valid = 1'b 1;
        fsm_err.code = ErrFatalError;
        fsm_err.info = 24'(app_id);
      end

      default: begin
        st_d = StTerminalError;
        sparse_fsm_error_o = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      st_d = StTerminalError;
    end
  end

  //////////////
  // Datapath //
  //////////////

  // Encoded output length
  assign encoded_outlen      = EncodedOutLen[SelDigSize];
  assign encoded_outlen_mask = EncodedOutLenMask[SelKeySize];

  // Data mux
  // This is the main part of the KeyMgr interface logic.
  // The FSM selects KeyMgr interface in a cycle after it receives the first
  // valid data from KeyMgr. The ready signal to the KeyMgr data interface
  // represents the MSG_FIFO ready, only when it is in StKeyMgrMsg state.
  // After KeyMgr sends last beat, the kmac interface (to MSG_FIFO) is switched
  // to OutLen. OutLen is pre-defined values. See `EncodeOutLen` parameter above.
  always_comb begin
    app_data_ready = 1'b 0;
    sw_ready_o = 1'b 1;

    kmac_valid_o = 1'b 0;
    kmac_data_o = '0;
    kmac_mask_o = '0;

    unique case (mux_sel_buf_kmac)
      SelApp: begin
        // app_id is valid at this time
        kmac_valid_o = app_i[app_id].valid;
        kmac_data_o  = app_i[app_id].data;
        // Expand strb to bits. prim_packer inside MSG_FIFO accepts the bit masks
        for (int i = 0 ; i < $bits(app_i[app_id].strb) ; i++) begin
          kmac_mask_o[8*i+:8] = {8{app_i[app_id].strb[i]}};
        end
        app_data_ready = kmac_ready_i;
      end

      SelOutLen: begin
        // Write encoded output length value
        kmac_valid_o = 1'b 1; // always write
        kmac_data_o  = MsgWidth'(encoded_outlen);
        kmac_mask_o  = MsgWidth'(encoded_outlen_mask);
      end

      SelSw: begin
        kmac_valid_o = sw_valid_i;
        kmac_data_o  = sw_data_i ;
        kmac_mask_o  = sw_mask_i ;
        sw_ready_o   = kmac_ready_i ;
      end

      default: begin // Incl. SelNone
        kmac_valid_o = 1'b 0;
        kmac_data_o = '0;
        kmac_mask_o = '0;
      end

    endcase
  end

  // Error checking for Mux
  always_comb begin
    mux_err = '{valid: 1'b 0, code: ErrNone, info: '0};

    if (mux_sel_buf_err_check != SelSw && sw_valid_i) begin
      // If SW writes message into FIFO
      mux_err = '{
        valid: 1'b 1,
        code: ErrSwPushedMsgFifo,
        info: 24'({8'h 00, 8'(st), 8'(mux_sel_buf_err_check)})
      };
    end else if (app_active_o && sw_cmd_i != CmdNone) begin
      // If SW issues command except start
      mux_err = '{
        valid: 1'b 1,
        code: ErrSwIssuedCmdInAppActive,
        info: 24'(sw_cmd_i)
      };
    end
  end

  logic [AppMuxWidth-1:0] mux_sel_buf_output_logic;
  assign mux_sel_buf_output = app_mux_sel_e'(mux_sel_buf_output_logic);

  // SEC_CM: LOGIC.INTEGRITY
  prim_sec_anchor_buf #(
   .Width(AppMuxWidth)
  ) u_prim_buf_state_output_sel (
    .in_i(mux_sel),
    .out_o(mux_sel_buf_output_logic)
  );

  logic [AppMuxWidth-1:0] mux_sel_buf_err_check_logic;
  assign mux_sel_buf_err_check = app_mux_sel_e'(mux_sel_buf_err_check_logic);

  // SEC_CM: LOGIC.INTEGRITY
  prim_sec_anchor_buf #(
   .Width(AppMuxWidth)
  ) u_prim_buf_state_err_check (
    .in_i(mux_sel),
    .out_o(mux_sel_buf_err_check_logic)
  );

  logic [AppMuxWidth-1:0] mux_sel_buf_kmac_logic;
  assign mux_sel_buf_kmac = app_mux_sel_e'(mux_sel_buf_kmac_logic);

  // SEC_CM: LOGIC.INTEGRITY
  prim_sec_anchor_buf #(
   .Width(AppMuxWidth)
  ) u_prim_buf_state_kmac_sel (
    .in_i(mux_sel),
    .out_o(mux_sel_buf_kmac_logic)
  );

  // SEC_CM: LOGIC.INTEGRITY
  logic reg_state_valid;
  prim_sec_anchor_buf #(
   .Width(1)
  ) u_prim_buf_state_output_valid (
    .in_i(reg_state_valid),
    .out_o(reg_state_valid_o)
  );

  // Keccak state Demux
  // Keccak state --> Register output is enabled when state is in StSw
  always_comb begin
    reg_state_valid = 1'b 0;
    reg_state_o = '{default:'0};
    if ((mux_sel_buf_output == SelSw) && (lc_escalate_en_i == lc_ctrl_pkg::Off)) begin
      reg_state_valid = keccak_state_valid_i;
      reg_state_o = keccak_state_i;
      // If key is sideloaded and KMAC is SW initiated
      // hide the capacity from SW by zeroing (see #17508)
      if (keymgr_key_en_i) begin
        for (int i = 0; i < Share; i++) begin
          unique case (reg_keccak_strength_i)
            L128: reg_state_o[i][sha3_pkg::StateW-1-:KeccakBitCapacity[L128]] = '0;
            L224: reg_state_o[i][sha3_pkg::StateW-1-:KeccakBitCapacity[L224]] = '0;
            L256: reg_state_o[i][sha3_pkg::StateW-1-:KeccakBitCapacity[L256]] = '0;
            L384: reg_state_o[i][sha3_pkg::StateW-1-:KeccakBitCapacity[L384]] = '0;
            L512: reg_state_o[i][sha3_pkg::StateW-1-:KeccakBitCapacity[L512]] = '0;
            default: reg_state_o[i] = '0;
          endcase
        end
      end
    end
  end

  // Keccak state --> KeyMgr
  always_comb begin
    app_digest_done = 1'b 0;
    app_digest = '{default:'0};
    if (st == StAppWait && prim_mubi_pkg::mubi4_test_true_strict(absorbed_i) &&
        lc_escalate_en_i == lc_ctrl_pkg::Off) begin
      // SHA3 engine has calculated the hash. Return the data to KeyMgr
      app_digest_done = 1'b 1;

      // digest has always 2 entries. If !EnMasking, second is tied to 0.
      for (int i = 0 ; i < Share ; i++) begin
        // Return the portion of state.
        app_digest[i] = keccak_state_i[i][AppDigestW-1:0];
      end
    end
  end


  // Secret Key Mux

  // Prepare merged key if EnMasking is not set.
  // Combine share keys into unpacked array for logic below to assign easily.
  // SEC_CM: KEY.SIDELOAD
  logic [MaxKeyLen-1:0] keymgr_key [Share];
  if (EnMasking == 1) begin : g_masked_key
    for (genvar i = 0; i < Share; i++) begin : gen_key_pad
      assign keymgr_key[i] =  {(MaxKeyLen-KeyMgrKeyW)'(0), keymgr_key_i.key[i]};
    end
  end else begin : g_unmasked_key
    always_comb begin
      keymgr_key[0] = '0;
      for (int i = 0; i < keymgr_pkg::Shares; i++) begin
        keymgr_key[0][KeyMgrKeyW-1:0] ^= keymgr_key_i.key[i];
      end
    end
  end

  // Sideloaded key manage: Keep use sideloaded key for KMAC AppIntf until the
  // hashing operation is finished.
  always_comb begin
    key_len_o  = reg_key_len_i;
    for (int i = 0 ; i < Share; i++) begin
      key_data_o[i] = reg_key_data_i[i];
    end

    unique case (st)
      StAppCfg, StAppMsg, StAppOutLen, StAppProcess, StAppWait: begin
        key_len_o = SideloadedKey;
        for (int i = 0 ; i < Share; i++) begin
          key_data_o[i] = keymgr_key[i];
        end
      end

      StSw: begin
        if (keymgr_key_en_i) begin
          key_len_o = SideloadedKey;
          for (int i = 0 ; i < Share; i++) begin
            key_data_o[i] = keymgr_key[i];
          end
        end
      end

      default: ;
    endcase
  end

  // Prefix Demux
  // For SW, always prefix register.
  // For App intf, check PrefixMode cfg and if 1, use Prefix cfg.
  always_comb begin
    sha3_prefix_o = '0;

    unique case (st)
      StAppCfg, StAppMsg, StAppOutLen, StAppProcess, StAppWait: begin
        // Check app intf cfg
        for (int unsigned i = 0 ; i < NumAppIntf ; i++) begin
          if (app_id == i) begin
            if (AppCfg[i].PrefixMode == 1'b 0) begin
              sha3_prefix_o = reg_prefix_i;
            end else begin
              sha3_prefix_o = AppCfg[i].Prefix;
            end
          end
        end
      end

      StSw: begin
        sha3_prefix_o = reg_prefix_i;
      end

      default: begin
        sha3_prefix_o = reg_prefix_i;
      end
    endcase
  end

  // KMAC en / SHA3 mode / Strength
  //  by default, it uses reg cfg. When app intf reqs come, it uses AppCfg.
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      kmac_en_o         <= 1'b 0;
      sha3_mode_o       <= sha3_pkg::Sha3;
      keccak_strength_o <= sha3_pkg::L256;
    end else if (clr_appid) begin
      // As App completed, latch reg value
      kmac_en_o         <= reg_kmac_en_i;
      sha3_mode_o       <= reg_sha3_mode_i;
      keccak_strength_o <= reg_keccak_strength_i;
    end else if (set_appid) begin
      kmac_en_o         <= AppCfg[arb_idx].Mode == AppKMAC ? 1'b 1 : 1'b 0;
      sha3_mode_o       <= AppCfg[arb_idx].Mode == AppSHA3
                           ? sha3_pkg::Sha3 : sha3_pkg::CShake;
      keccak_strength_o <= AppCfg[arb_idx].Strength ;
    end else if (st == StIdle) begin
      kmac_en_o         <= reg_kmac_en_i;
      sha3_mode_o       <= reg_sha3_mode_i;
      keccak_strength_o <= reg_keccak_strength_i;
    end
  end

  // Status
  assign app_active_o = (st inside {StAppCfg, StAppMsg, StAppOutLen,
                                    StAppProcess, StAppWait});

  // Error Reporting ==========================================================
  always_comb begin
    priority casez ({fsm_err.valid, mux_err.valid})
      2'b ?1: error_o = mux_err;
      2'b 10: error_o = fsm_err;
      default: error_o = '{valid: 1'b0, code: ErrNone, info: '0};
    endcase
  end

  ////////////////
  // Assertions //
  ////////////////

  // KeyMgr sideload key and the digest should be in the Key Length value
  `ASSERT_INIT(SideloadKeySameToDigest_A, KeyMgrKeyW <= AppDigestW)
  `ASSERT_INIT(AppIntfInRange_A, AppDigestW inside {128, 192, 256, 384, 512})

  // Issue(#13655): Having a coverage that sideload keylen and CSR keylen are
  // different.
  `COVER(AppIntfUseDifferentSizeKey_C,
    (st == StAppCfg && kmac_en_o) |-> reg_key_len_i != SideloadedKey)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// KMAC Entropy Generation module

`include "prim_assert.sv"

module kmac_entropy
  import kmac_pkg::*;
  import kmac_reg_pkg::*;
#(
  parameter lfsr_perm_t RndCnstLfsrPerm = RndCnstLfsrPermDefault,
  parameter lfsr_seed_t RndCnstLfsrSeed = RndCnstLfsrSeedDefault,
  parameter lfsr_fwd_perm_t RndCnstLfsrFwdPerm = RndCnstLfsrFwdPermDefault
) (
  input clk_i,
  input rst_ni,

  // EDN interface
  output logic                            entropy_req_o,
  input                                   entropy_ack_i,
  input [edn_pkg::ENDPOINT_BUS_WIDTH-1:0] entropy_data_i,

  // Entropy to internal
  output logic                          rand_valid_o,
  output logic                          rand_early_o,
  output logic [sha3_pkg::StateW/2-1:0] rand_data_o,
  output logic                          rand_aux_o,
  input                                 rand_consumed_i,

  // Status
  input in_keyblock_i,

  // Configurations
  input entropy_mode_e mode_i,
  //// SW sets ready bit when EDN is ready to accept requests through its app.
  //// interface.
  input entropy_ready_i,

  //// Garbage random value when not processing Keyblock, if this config is
  //// turned on, the logic sending garbage value and never de-assert
  //// rand_valid_o unless it is not processing KeyBlock.
  input fast_process_i,

  //// LFSR Enable for Message Masking
  //// If 1, LFSR advances to create 64-bit PRNG. This input is used to mask
  //// the message fed into SHA3 (Keccak).
  input                       msg_mask_en_i,
  output logic [MsgWidth-1:0] msg_mask_o,

  //// SW update of seed
  input [NumSeedsEntropyLfsr-1:0]       seed_update_i,
  input [NumSeedsEntropyLfsr-1:0][31:0] seed_data_i,

  //// SW may initiate manual EDN seed refresh
  input entropy_refresh_req_i,

  //// Timer limit value
  //// If value is 0, timer is disabled
  input [TimerPrescalerW-1:0] wait_timer_prescaler_i,
  input [EdnWaitTimerW-1:0]   wait_timer_limit_i,

  // Status out
  //// Hash Ops counter. Count how many hashing ops (KMAC) have run
  //// after the clear request from SW
  output logic [HashCntW-1:0] hash_cnt_o,
  input                       hash_cnt_clr_i,
  input        [HashCntW-1:0] hash_threshold_i,

  output prim_mubi_pkg::mubi4_t entropy_configured_o,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  // Error output
  output err_t err_o,
  output logic sparse_fsm_error_o,
  output logic count_error_o,
  input        err_processed_i
);

  /////////////////
  // Definitions //
  /////////////////

  // Timer Widths are defined in kmac_pkg

  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 9 -n 10 \
  //      -s 507672272 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: ||||||||||| (13.89%)
  //  4: ||||||||||||||| (19.44%)
  //  5: |||||||||||||||||||| (25.00%)
  //  6: ||||||||||||||| (19.44%)
  //  7: ||||||||||| (13.89%)
  //  8: |||| (5.56%)
  //  9: || (2.78%)
  // 10: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 9
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 7
  //
  localparam int StateWidth = 10;

  // States
  typedef enum logic [StateWidth-1:0] {
    // Reset: Reset state. The entropy is not ready. The state machine should
    // get new entropy from EDN or the seed should be feeded by the software.
    StRandReset = 10'b1001111000,

    // The seed is fed into LFSR and the entropy is ready. It means the
    // rand_valid is asserted with valid data. It takes a few steps to reach
    // this state from StRandReset.
    StRandReady = 10'b0110000100,

    // EDN interface: Send request and receive
    // RandEdnReq state can be transit from StRandReset or from StRandReady
    //
    // Reset --> EdnReq:
    //     If entropy source module is ready, the software sets a bit in CFG
    //     also sets the entropy mode to EdnMode. Then this FSM moves to EdnReq
    //     to initialize LFSR seed.
    //
    // Ready --> EdnReq:
    //     1. If a mode is configured as to update entropy everytime it is
    //        consumed, then the FSM moves from Ready to EdnReq to refresh seed
    //     2. If the software enabled EDN timer and the timer is expired and
    //        also the KMAC is processing the key block, the FSM moves to
    //        EdnReq to refresh seed
    //     3. If a KMAC operation is completed, the FSM also refreshes the LFSR
    //        seed to prepare next KMAC op or wipe out operation.
    StRandEdn = 10'b1100100111,

    // Sw Seed: If mode is set to manual mode, This entropy module needs initial
    // seed from the software. It waits the seed update signal to expand initial
    // entropy
    StSwSeedWait = 10'b1011110110,

    // Generate: In this state, the entropy generator advances the LFSRs to
    // generate the 800-bits of pseudo random data for the next evaluation.
    StRandGenerate = 10'b0000001100,

    // ErrWaitExpired: If Edn timer expires, FSM moves to this state and wait
    // the software response. Software should switch to manual mode then disable
    // the timer (to 0) and update the seed via register interface.
    StRandErrWaitExpired = 10'b0001100011,

    // ErrNoValidMode: If SW sets entropy ready but the mode is not either
    // Manual Mode nor EdnMode, this logic reports to SW with
    // NoValidEntropyMode.
    StRandErrIncorrectMode = 10'b1110010000,

    // Err: After the error is reported, FSM sits in Err state ignoring all the
    // requests. It does not generate new entropy and drops the entropy valid
    // signal.
    //
    // SW sets err_processed signal to clear the error. The software should
    // clear the entropy ready signal before clear the error interrupt so that
    // the FSM sits in StRandReset state not moving forward with incorrect
    // configurations.
    StRandErr = 10'b1000011110,

    StTerminalError = 10'b0010011000
  } rand_st_e;

  /////////////
  // Signals //
  /////////////

  // Timers
  // "Wait Timer": This timer is in active when FSM sends entropy request to EDN
  //   If EDN does not return the entropy data until the timer expired, FSM
  //   moves to error state and report the error to the system.

  localparam int unsigned TimerW = EdnWaitTimerW;
  logic timer_enable, timer_update, timer_expired, timer_pulse;
  logic [TimerW-1:0] timer_limit;
  logic [TimerW-1:0] timer_value;

  localparam int unsigned PrescalerW = TimerPrescalerW;
  logic [PrescalerW-1:0] prescaler_cnt;

  // LFSR
  // SW configures to use EDN or SEED register as a LFSR seed
  logic [NumSeedsEntropyLfsr-1:0]                            lfsr_seed_en_red;
  logic [NumChunksEntropyLfsr-1:0]                           lfsr_seed_en;
  logic [NumChunksEntropyLfsr-1:0][ChunkSizeEntropyLfsr-1:0] lfsr_seed;
  logic lfsr_seed_done;
  logic lfsr_en;
  logic [NumChunksEntropyLfsr-1:0][ChunkSizeEntropyLfsr-1:0] lfsr_data_chunked;
  logic [EntropyLfsrW-1:0] lfsr_data, lfsr_data_permuted;

  // Auxliliary randomness
  logic aux_rand_d, aux_rand_q;
  logic aux_update;

  // Randomness for controlling PRNG updates. This only matters for clock cycles
  // where the PRNG output is not actually used.
  logic [3:0] lfsr_en_rand_d, lfsr_en_rand_q;

  // Entropy valid signal
  // FSM set and clear the valid signal, rand_consume signal clear the valid
  // signal. Split the set, clear to make entropy valid while FSM is processing
  // other tasks.
  logic rand_valid_set, rand_valid_clear;

  // Signal to track whether the FSM should stay in the StRandReady state or
  // move to StRandGenerate upon getting the next rand_consumed_i.
  logic ready_phase_d, ready_phase_q;

  // FSM latches the mode and stores into mode_q when the FSM is out from
  // StReset. The following states, or internal datapath uses mode_q after that.
  // If the SW wants to change the mode, it requires resetting the IP.
  logic mode_latch;
  entropy_mode_e mode_q;

  // Status out: entropy configured
  prim_mubi_pkg::mubi4_t entropy_configured;

  //////////////
  // Datapath //
  //////////////

  // For latching (`wait_timer_limit_i` != 0) during last `timer_update`
  // See #16716
  logic non_zero_wait_timer_limit;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      non_zero_wait_timer_limit <= '0;
    end else if (timer_update) begin
      non_zero_wait_timer_limit <= |wait_timer_limit_i;
    end
  end

  logic [TimerPrescalerW-1:0] wait_timer_prescaler_d;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      wait_timer_prescaler_d <= '0;
    end else if (timer_update) begin
      wait_timer_prescaler_d <= wait_timer_prescaler_i;
    end
  end

  // Timers ===================================================================
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      timer_value <= '0;
    end else if (timer_update) begin
      timer_value <= timer_limit;
    end else if (timer_expired) begin
      timer_value <= '0; // keep the value
    end else if (timer_enable && timer_pulse && |timer_value) begin // if non-zero timer v
      timer_value <= timer_value - 1'b 1;
    end
  end

  assign timer_limit = TimerW'(wait_timer_limit_i);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      timer_expired <= 1'b 0;
    end else if (timer_update) begin
      timer_expired <= 1'b 0;
    end else if (timer_enable && (timer_value == '0)) begin
      timer_expired <= 1'b 1;
    end
  end

  // Prescaler
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      prescaler_cnt <= '0;
    end else if (timer_update) begin
      prescaler_cnt <= wait_timer_prescaler_i;
    end else if (timer_enable && prescaler_cnt == '0) begin
      prescaler_cnt <= wait_timer_prescaler_d;
    end else if (timer_enable) begin
      prescaler_cnt <= prescaler_cnt - 1'b 1;
    end
  end

  assign timer_pulse = (timer_enable && prescaler_cnt == '0);
  // Timers -------------------------------------------------------------------

  // Hash Counter
  logic threshold_hit;
  logic threshold_hit_q, threshold_hit_clr; // latched hit

  logic hash_progress_d, hash_progress_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) hash_progress_q <= 1'b 0;
    else         hash_progress_q <= hash_progress_d;
  end

  assign hash_progress_d = in_keyblock_i;

  logic hash_cnt_clr;
  assign hash_cnt_clr = hash_cnt_clr_i || threshold_hit || entropy_refresh_req_i;

  logic hash_cnt_en;
  assign hash_cnt_en = hash_progress_q && !hash_progress_d;

  logic hash_count_error;

  // SEC_CM CTR.REDUN
  // This primitive is used to place a hardened counter
  prim_count #(
    .Width(HashCntW)
  ) u_hash_count (
    .clk_i,
    .rst_ni,
    .clr_i(hash_cnt_clr),
    .set_i(1'b0),
    .set_cnt_i(HashCntW'(0)),
    .incr_en_i(hash_cnt_en),
    .decr_en_i(1'b0),
    .step_i(HashCntW'(1)),
    .cnt_o(hash_cnt_o),
    .cnt_next_o(),
    .err_o(hash_count_error)
  );

  assign threshold_hit = |hash_threshold_i && (hash_threshold_i <= hash_cnt_o);

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)                threshold_hit_q <= 1'b 0;
    else if (threshold_hit_clr) threshold_hit_q <= 1'b 0;
    else if (threshold_hit)     threshold_hit_q <= 1'b 1;
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)         mode_q <= EntropyModeNone;
    else if (mode_latch) mode_q <= mode_i;
  end

  // LFSRs ====================================================================

  // We use 25 32-bit LFSRs in parallel to generate the 800 bits of randomness
  // required by the DOM multipliers inside the Keccak core in a single clock
  // cycle. To reduce the entropy consumption for periodic reseeding, a cascaded
  // reseeding mechanism is used:
  //
  // - LFSR 0 (5/10/15/20) gets one 32-bit seed each from EDN/SW.
  // - LFSR 1 (6/11/16/21) gets the old state of LFSR 0 (5/10/15/20)
  // - ...
  // - LFSR 4 (9/14/19/24) gets the old state of LFSR 3 (8/13/18/23)
  //
  // In addition, the forwarded old states are permuted.
  //
  // This allows to reduce the entropy consumption. A full reseed of all 25
  // LFSRs is still possible by subsequently triggering 5 reseeding operations
  // though software.

  // Reseeding counter - We reseed one 32-bit chunk at a time and need to keep
  // track of which LFSR chunk to reseed next.
  localparam int unsigned SeedIdxWidth =
      prim_util_pkg::vbits(NumSeedsEntropyLfsr);
  logic [SeedIdxWidth-1:0] seed_idx;
  logic seed_idx_count_error;

  // SEC_CM CTR.REDUN
  // This primitive is used to place a hardened counter
  prim_count #(
    .Width(SeedIdxWidth)
  ) u_seed_idx_count (
    .clk_i,
    .rst_ni,
    .clr_i(lfsr_seed_done),
    .set_i(1'b0),
    .set_cnt_i(SeedIdxWidth'(0)),
    .incr_en_i(|lfsr_seed_en),
    .decr_en_i(1'b0),
    .step_i(SeedIdxWidth'(1)),
    .cnt_o(seed_idx),
    .cnt_next_o(),
    .err_o(seed_idx_count_error)
  );

  assign lfsr_seed_done =
      (seed_idx == SeedIdxWidth'(unsigned'(NumSeedsEntropyLfsr - 1))) &
      |lfsr_seed_en;

  // Seed selection - The reduced seed enable signal `lfsr_seed_en_red` is
  // controlled by the FSM. Here we just repliate it as we're always reseeding
  // 5 LFSRs together.
  for (genvar i = 0; i < 5; i++) begin : gen_lfsr_seed_en
    assign lfsr_seed_en[i * 5 +: 5] = {5{lfsr_seed_en_red[i]}};
  end

  // From software we get NumChunks 32-bit seeds but only one is valid. The
  // others may be zero.
  // From EDN we get a single 32-bit seed. This is the default value forwarded.
  for (genvar i = 0; i < NumSeedsEntropyLfsr; i++) begin : gen_lfsr_seed
    // LFSRs 0/5/10/15/20 get the fresh entropy.
    assign lfsr_seed[i * 5] =
        (mode_q == EntropyModeSw) ? seed_data_i[i] : entropy_data_i;

    // The other LFSRs get the permuted old states.
    for (genvar j = 0; j < 4; j++) begin : gen_fwd_seeds
      for (genvar k = 0; k < ChunkSizeEntropyLfsr; k++) begin : gen_fwd_perm
        assign lfsr_seed[i * 5 + j + 1][k] =
            lfsr_data_chunked[i * 5 + j][RndCnstLfsrFwdPerm[k]];
      end
    end
  end
  `ASSERT_KNOWN(ModeKnown_A, mode_i)

  // We employ five 32-bit LFSRs to generate 160 bits per clock cycle. Using
  // multiple 32-bit LFSRs with an additional permutation layer spanning across
  // all LFSRs has relevant advantages:
  // - Multiple simulateneous faults needs to be injected to get a fully
  //   deterministic output.
  // - No additional buffering is needed for reseeding. Both software and EDN
  //   provide 32 bits at a time meaning we can reseed the LFSRs directly as
  //   we get the entropy.
  // We use multiple LFSR instances each having a width of ChunkSize.
  for (genvar i = 0; i < NumChunksEntropyLfsr; i++) begin : gen_lfsrs
    prim_lfsr #(
      .LfsrType("GAL_XOR"),
      .LfsrDw(ChunkSizeEntropyLfsr),
      .StateOutDw(ChunkSizeEntropyLfsr),
      .DefaultSeed(RndCnstLfsrSeed[i * ChunkSizeEntropyLfsr +: ChunkSizeEntropyLfsr]),
      .StatePermEn(1'b0),
      .NonLinearOut(1'b1)
    ) u_lfsr_chunk (
      .clk_i,
      .rst_ni,
      .seed_en_i(lfsr_seed_en[i]),
      .seed_i   (lfsr_seed[i]),
      .lfsr_en_i(lfsr_en || msg_mask_en_i),
      .entropy_i('0),
      .state_o  (lfsr_data_chunked[i])
    );
  end

  // Add a permutation layer spanning across all LFSRs to break linear shift
  // patterns.
  assign lfsr_data = lfsr_data_chunked;
  for (genvar i = 0; i < EntropyLfsrW; i++) begin : gen_perm
    assign lfsr_data_permuted[i] = lfsr_data[RndCnstLfsrPerm[i]];
  end

  // Forwrad LSBs for masking the message.
  assign msg_mask_o = lfsr_data_permuted[MsgWidth-1:0];

  // LFSRs --------------------------------------------------------------------

  // Auxiliary randomness =====================================================
  assign aux_rand_d = aux_update ? lfsr_data_permuted[EntropyLfsrW - 1] :
                                   aux_rand_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      aux_rand_q <= '0;
    end else begin
      aux_rand_q <= aux_rand_d;
    end
  end

  // Auxiliary randomness -----------------------------------------------------

  // LFSR enable randomness ===================================================
  assign lfsr_en_rand_d =
      aux_update ? lfsr_data_permuted[EntropyLfsrW - 2 -: 4] : // refresh
                   {1'b0, lfsr_en_rand_q[3:1]};                // shift out

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      lfsr_en_rand_q <= '0;
    end else begin
      lfsr_en_rand_q <= lfsr_en_rand_d;
    end
  end

  // LFSR enable randomness ---------------------------------------------------

  // Randomness outputs =======================================================
  assign rand_data_o = lfsr_data_permuted;
  assign rand_aux_o = aux_rand_q;

  // entropy valid
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rand_valid_o <= 1'b 0;
    end else if (rand_valid_set) begin
      rand_valid_o <= 1'b 1;
    end else if (rand_valid_clear) begin
      rand_valid_o <= 1'b 0;
    end
  end

  // Let consumers know that the randomness will be valid in the next clock cycle.
  assign rand_early_o = rand_valid_set;

  `ASSUME(ConsumeNotAseertWhenNotReady_M, rand_consumed_i |-> rand_valid_o)

  // Randomness outputs -------------------------------------------------------

  // Remaining outputs
  assign count_error_o = hash_count_error | seed_idx_count_error;

  ///////////////////
  // State Machine //
  ///////////////////

  rand_st_e st, st_d;

  // State FF
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, st_d, st, rand_st_e, StRandReset)

  // State: Next State and Output Logic
  // SEC_CM: FSM.SPARSE
  always_comb begin
    st_d = st;
    sparse_fsm_error_o = 1'b 0;

    // Default Timer values
    timer_enable = 1'b 0;
    timer_update = 1'b 0;

    threshold_hit_clr = 1'b 0;

    // EDN request
    entropy_req_o = 1'b 0;

    // rand is valid when this logic expands the entropy.
    // FSM sets the valid signal, the signal is cleared by `consume` signal
    // or FSM clear signal.
    // Why split the signal to set and clear?
    // FSM only set the signal to make entropy valid while processing other
    // tasks such as EDN request.
    rand_valid_set   = 1'b 0;
    rand_valid_clear = 1'b 0;

    // mode_latch to store mode_i into mode_q
    mode_latch = 1'b 0;

    // lfsr_en: Let LFSR run
    // To save power, this logic enables LFSR when it needs entropy expansion.
    lfsr_en = 1'b 0;

    // lfsr_seed_en_red: Signal to update LFSR seed
    // LFSR seed can be updated by EDN or SW.
    lfsr_seed_en_red = '0;

    // Signal to track whether FSM should stay in StRandReady state or move on.
    ready_phase_d = ready_phase_q;

    // Auxiliary randomness control signals
    aux_update = 1'b 0;

    // Error
    err_o = '{valid: 1'b 0, code: ErrNone, info: '0};

    unique case (st)
      StRandReset: begin
        if (entropy_ready_i) begin

          // As SW ready, discard current dummy entropy and refresh.
          rand_valid_clear = 1'b 1;

          mode_latch = 1'b 1;
          // SW has configured KMAC
          unique case (mode_i)
            EntropyModeSw: begin
              st_d = StSwSeedWait;
            end

            EntropyModeEdn: begin
              st_d = StRandEdn;

              // Timer reset
              timer_update = 1'b 1;
            end

            default: begin
              // EntropyModeNone or other values
              // Error. No valid mode given, report to SW
              st_d = StRandErrIncorrectMode;
            end
          endcase
        end else begin
          st_d = StRandReset;

          // Setting the dummy rand gate until SW prepares.
          // This lets the Application Interface move forward out of reset
          // without SW intervention.
          rand_valid_set = 1'b 1;
        end
      end

      StRandReady: begin
        timer_enable = 1'b 1; // If limit is zero, timer won't work

        lfsr_en = lfsr_en_rand_q[0];

        if (rand_consumed_i &&
            ((fast_process_i && in_keyblock_i) || !fast_process_i)) begin
          // If fast_process is set, don't clear the rand valid, even
          // consumed. So, the logic does not expand the entropy again.
          // If fast_process is not set, then every rand_consume signal
          // triggers rand expansion.

          // Allow for two reads from the Keccak core. This is what is needed
          // per round.
          lfsr_en = 1'b 1;
          ready_phase_d = ~ready_phase_q;

          if (ready_phase_q) begin
            st_d = StRandGenerate;

            rand_valid_clear = 1'b 1;
          end else begin
            st_d = StRandReady;
          end
        end else if ((mode_q == EntropyModeEdn) &&
            (entropy_refresh_req_i || threshold_hit_q)) begin
          st_d = StRandEdn;

          // Timer reset
          timer_update = 1'b 1;

          // Clear the threshold as it refreshes the hash
          threshold_hit_clr = 1'b 1;
        end else begin
          st_d = StRandReady;
        end
      end

      StRandEdn: begin
        // Send request
        entropy_req_o = 1'b 1;

        // Wait timer
        timer_enable = 1'b 1;

        if (timer_expired && non_zero_wait_timer_limit) begin
          // If timer count is non-zero and expired;
          st_d = StRandErrWaitExpired;

        end else if (entropy_ack_i) begin
          lfsr_seed_en_red[seed_idx] = 1'b 1;

          if (lfsr_seed_done) begin
            st_d = StRandGenerate;

            if ((fast_process_i && in_keyblock_i) || !fast_process_i) begin
              lfsr_en = 1'b 1;
              rand_valid_clear = 1'b 1;
            end
          end else begin
            st_d = StRandEdn;
          end
        end else if (rand_consumed_i &&
            ((fast_process_i && in_keyblock_i) || !fast_process_i)) begin
          // Somehow, while waiting the EDN entropy, the KMAC or SHA3 logic
          // consumed the remained entropy. This can happen when the previous
          // SHA3/ KMAC op completed and this Entropy FSM has moved to this
          // state to refresh the entropy and the SW initiates another hash
          // operation while waiting for the EDN response.
          st_d = StRandEdn;

          rand_valid_clear = 1'b 1;
        end else begin
          st_d = StRandEdn;
        end
      end

      StSwSeedWait: begin
        lfsr_seed_en_red = seed_update_i;

        if (lfsr_seed_done) begin
          st_d = StRandGenerate;

          lfsr_en = 1'b 1;

          rand_valid_clear = 1'b 1;
        end else begin
          st_d = StSwSeedWait;
        end
      end

      StRandGenerate: begin
        // The current LFSR output is used as auxiliary randomness.
        aux_update = 1'b 1;

        // Advance the LFSR and set the valid bit. The next LFSR output will be
        // used for re-masking.
        lfsr_en = 1'b 1;
        rand_valid_set = 1'b 1;

        st_d = StRandReady;
      end

      StRandErrWaitExpired: begin
        st_d = StRandErr;

        err_o = '{ valid: 1'b 1,
                   code: ErrWaitTimerExpired,
                   info: 24'(timer_value)
                 };
      end

      StRandErrIncorrectMode: begin
        st_d = StRandErr;

        err_o = '{ valid: 1'b 1,
                   code: ErrIncorrectEntropyMode,
                   info: 24'(mode_q)
                 };
      end

      StRandErr: begin
        // Keep entropy signal valid to complete current hashing even with error
        rand_valid_set = 1'b 1;

        if (err_processed_i) begin
          st_d = StRandReset;

        end else begin
          st_d = StRandErr;
        end

      end

      StTerminalError: begin
        // this state is terminal
        st_d = st;
        sparse_fsm_error_o = 1'b 1;
      end

      default: begin
        st_d = StTerminalError;
        sparse_fsm_error_o = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      st_d = StTerminalError;
    end
  end
  `ASSERT_KNOWN(RandStKnown_A, st)

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      ready_phase_q <= '0;
    end else begin
      ready_phase_q <= ready_phase_d;
    end
  end

  // mubi4 sender

  assign entropy_configured = (st != StRandReset)
                            ? prim_mubi_pkg::MuBi4True
                            : prim_mubi_pkg::MuBi4False ;
  prim_mubi4_sender #(
    .AsyncOn(1'b0)
  ) u_entropy_configured (
    .clk_i,
    .rst_ni,

    .mubi_i (entropy_configured  ),
    .mubi_o (entropy_configured_o)
  );

  ////////////////
  // Assertions //
  ////////////////

  `ASSERT_INIT(EntropyLfsrWDivisble, NumChunksEntropyLfsr ==
      EntropyLfsrW / ChunkSizeEntropyLfsr)

  // We reseed one chunk of the entropy generator at a time. Therefore the
  // chunk size must match the data width of the software and EDN inputs.
  `ASSERT_INIT(ChunkSizeEntropyLfsrMatchesSw, ChunkSizeEntropyLfsr == 32)
  `ASSERT_INIT(ChunkSizeEntropyLfsrMatchesEdn, ChunkSizeEntropyLfsr ==
      edn_pkg::ENDPOINT_BUS_WIDTH)

// the code below is not meant to be synthesized,
// but it is intended to be used in simulation and FPV
`ifndef SYNTHESIS
  // Check that the supplied permutations are valid.
  logic [EntropyLfsrW-1:0] perm_test;
  initial begin : p_perm_check
    perm_test = '0;
    for (int k = 0; k < EntropyLfsrW; k++) begin
      perm_test[RndCnstLfsrPerm[k]] = 1'b1;
    end
    // All bit positions must be marked with 1.
    `ASSERT_I(PermutationCheck_A, &perm_test)
  end

  logic [ChunkSizeEntropyLfsr-1:0] perm_fwd_test;
  initial begin : p_perm_fwd_check
    perm_fwd_test = '0;
    for (int k = 0; k < ChunkSizeEntropyLfsr; k++) begin
      perm_fwd_test[RndCnstLfsrFwdPerm[k]] = 1'b1;
    end
    // All bit positions must be marked with 1.
    `ASSERT_I(PermutationCheck_A, &perm_fwd_test)
  end
`endif

endmodule : kmac_entropy


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// KMAC Error Checking logic
//
// `kmac_err` module checks the SW introduced errors.
//  1. SW command sequencing error.
//  2. SW configuration error.
//
// ## SW Command Sequencing Error
//
// KMAC assumes the application interface and the SW register interface to
// follow the specific sequence. It expects the requester to send the `Start`
// command then push the message body. The `Process` command follows the message
// body. The SW may issue `Run` command if it needs the digest result more than
// a block rate. Then SW completes the hash operation with `Done` command.
//
// This `kmac_err` module checks if the SW issues the correct command. If not,
// it reports the error via ERR_CODE register.
//
// However, the logic does not prevent the error-ed command to be propagated.
// The unexpected commands are filtered by each individual submodule.
//
// st := { Idle, MsgFeed, Processing, Absorbed, Squeeze}
//
// allowed := {
//   Idle :      { Start     },
//   MsgFeed:    { Process   },
//   Processing: { None      },
//   Absorbed:   { Run, Done },
//   Squeeze:    { None      }
// }
//
// ## SW Configuration Error
//
// `kmac_errchk` module checks if SW configured correct combinations of the
// configuration registers when the hashing operation begins.
//
// 1. Mode & Strength combinations
// 2. Kmac Prefix
// * sideload & key_valid -> Checker in kmac_core

`include "prim_assert.sv"

module kmac_errchk
  import kmac_pkg::*;
  import sha3_pkg::sha3_mode_e;
  import sha3_pkg::keccak_strength_e;
#(
  parameter bit EnMasking = 1'b 1
) (
  input clk_i,
  input rst_ni,

  // Configurations
  input sha3_mode_e       cfg_mode_i,
  input keccak_strength_e cfg_strength_i,

  input        kmac_en_i,
  input [47:0] cfg_prefix_6B_i, // first 6B of PREFIX

  // If the signal below is set, errchk propagates the command to the rest of
  // the blocks even with err_modestrength.
  input        cfg_en_unsupported_modestrength_i,

  // Entropy Ready Status to check if SW initiated the hahs without entropy cfg
  input        entropy_ready_pulse_i,

  // SW commands: Only valid command is sent out to the rest of the modules
  input  kmac_cmd_e sw_cmd_i,
  output kmac_cmd_e sw_cmd_o,

  // Status from KMAC_APP
  input app_active_i,

  // Status from SHA3 core
  input prim_mubi_pkg::mubi4_t sha3_absorbed_i,
  input keccak_done_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  // Error processed indicator
  input err_processed_i,

  output err_t error_o,
  output logic sparse_fsm_error_o
);

  // sha3_pkg::sha3_mode_e
  import sha3_pkg::L128;
  import sha3_pkg::L224;
  import sha3_pkg::L256;
  import sha3_pkg::L384;
  import sha3_pkg::L512;

  // sha3_pkg::keccak_strength_e
  import sha3_pkg::Sha3;
  import sha3_pkg::Shake;
  import sha3_pkg::CShake;

  /////////////////
  // Definitions //
  /////////////////
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 5 -n 6 \
  //      -s 2239170217 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (50.00%)
  //  4: |||||||||||||||| (40.00%)
  //  5: |||| (10.00%)
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 5
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 4
  //
  localparam int StateWidth = 6;
  typedef enum logic [StateWidth-1:0] {
    StIdle = 6'b001101,
    StMsgFeed = 6'b110001,
    StProcessing = 6'b010110,
    StAbsorbed = 6'b100010,
    StSqueezing = 6'b111100,
    StTerminalError = 6'b011011
  } st_e;
  st_e st, st_d;

  localparam int StateWidthL = 3;
  typedef enum logic [StateWidthL-1:0] {
    StIdleL,
    StMsgFeedL,
    StProcessingL,
    StAbsorbedL,
    StSqueezingL,
    StErrorL
  } st_logical_e;
  st_logical_e stL;


  /////////////
  // Signals //
  /////////////

  // `err_swsequence` occurs when SW issues wrong command
  logic err_swsequence;

  // `err_modestrength` occcurs when Mode & Strength combinations are not
  // allowed. This error does not block the hashing operation.
  // UnexpectedModeStrength may stop the processing based on CFG
  // The error raises when SW issues CmdStart.
  logic err_modestrength;

  // `err_prefix` occurs when the first 6B of !!PREFIX is not
  // `encode_string("KMAC")` and kmac is enabled. This error does not block the
  // KMAC operation.
  logic err_prefix;

  // `err_entropy_ready` occurs when SW initiated the hashing op. without
  // configuring the entropy. This error may happen only when EnMasking is
  // set.
  logic err_entropy_ready;

  // entropy_ready is a pulse signal. Logic needs to store the state.
  logic cfg_entropy_ready;

  // Signal to block the SW command propagation
  logic block_swcmd;

  ///////////////////
  // Error Checker //
  ///////////////////

  // SW sequence Error
  // info field: Current state, Received command
  // SEC_CM: FSM.SPARSE
  always_comb begin
    err_swsequence = 1'b 0;
    sparse_fsm_error_o = 1'b 0;

    unique case (st)
      StIdle: begin
        // Allow Start command only
        if (!(sw_cmd_i inside {CmdNone, CmdStart})) begin
          err_swsequence = 1'b 1;
        end
      end

      StMsgFeed: begin
        // Allow Process only
        if (!(sw_cmd_i inside {CmdNone, CmdProcess})) begin
          err_swsequence = 1'b 1;
        end
      end

      StProcessing: begin
        if (sw_cmd_i != CmdNone) begin
          err_swsequence = 1'b 1;
        end
      end

      StAbsorbed: begin
        // Allow ManualRun and Done
        if (!(sw_cmd_i inside {CmdNone, CmdManualRun, CmdDone})) begin
          err_swsequence = 1'b 1;
        end
      end

      StSqueezing: begin
        if (sw_cmd_i != CmdNone) begin
          err_swsequence = 1'b 1;
        end
      end

      StTerminalError: begin
        err_swsequence = 1'b 0;
        sparse_fsm_error_o = 1'b 1;
      end

      default: begin
        err_swsequence = 1'b 0;
        sparse_fsm_error_o = 1'b 1;
      end
    endcase
  end

  assign block_swcmd =  (err_swsequence)
                     || (err_modestrength
                         && !cfg_en_unsupported_modestrength_i)
                     || err_entropy_ready;

  // sw_cmd_o latch
  // To reduce the command path delay, sw_cmd is latched here
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni)           sw_cmd_o <= CmdNone;
    else if (!block_swcmd) sw_cmd_o <= sw_cmd_i;
  end

  // Mode & Strength
  always_comb begin : check_modestrength
    err_modestrength = 1'b 0;

    if (st == StIdle && st_d == StMsgFeed) begin
      // When moving to the next stage, checks the config
      if (!((cfg_mode_i == Sha3 &&
             cfg_strength_i inside {L224, L256, L384, L512}) ||
            ((cfg_mode_i == Shake || cfg_mode_i == CShake) &&
             (cfg_strength_i inside {L128, L256})))) begin
        err_modestrength = 1'b 1;
      end
    end
  end : check_modestrength


  // Check prefix 6B is `encode_string("KMAC")`
  always_comb begin : check_prefix
    err_prefix = 1'b 0;

    if (st == StIdle && st_d == StMsgFeed && kmac_en_i) begin
      if (cfg_prefix_6B_i != EncodedStringKMAC) begin
        err_prefix = 1'b 1;
      end
    end
  end : check_prefix

  if (EnMasking) begin : g_entropy_chk

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni)              cfg_entropy_ready <= 1'b 0;
      else if (err_processed_i) cfg_entropy_ready <= 1'b 0;
      else if (entropy_ready_pulse_i && st == StIdle) begin
        cfg_entropy_ready <= 1'b 1;
      end
    end

    always_comb begin : check_entropy_ready
      err_entropy_ready = 1'b 0;

      if (st == StIdle && st_d == StMsgFeed && kmac_en_i) begin
        if (!cfg_entropy_ready) begin
          err_entropy_ready = 1'b 1;
        end
      end
    end : check_entropy_ready

  end else begin : g_pseudo_entropy_chk

    // If EnMasking is 0, entropy module is not generated.
    // tying the error signal to 0.
    assign err_entropy_ready = 1'b 0;

    assign cfg_entropy_ready = 1'b 1;

    logic unused_cfg_entropy_ready;
    assign unused_cfg_entropy_ready = cfg_entropy_ready;

  end

  always_comb begin : recode_st
    unique case (st)
      StIdle       : stL = StIdleL;
      StMsgFeed    : stL = StMsgFeedL;
      StProcessing : stL = StProcessingL;
      StAbsorbed   : stL = StAbsorbedL;
      StSqueezing  : stL = StSqueezingL;
      default      : stL = StErrorL;
    endcase
  end : recode_st

  // Return error code
  err_t err;
  always_comb begin : err_return
    err = '{valid: 1'b0, code: ErrNone, info: '0};

    priority case (1'b 1)
      err_swsequence: begin
        err = '{ valid: 1'b 1,
                 code: ErrSwCmdSequence,
                 info: {5'h0,
                        {err_swsequence, err_modestrength, err_prefix},
                        {5'h 0, stL},
                        {2'b0, sw_cmd_i}
                       }
               };
      end

      err_modestrength: begin
        err = '{ valid: 1'b 1,
                 code:  ErrUnexpectedModeStrength,
                 info:  { 5'h 0,
                          {err_swsequence, err_modestrength, err_prefix},
                          8'h 0,
                          {2'b 00, cfg_mode_i},
                          {1'b 0,  cfg_strength_i}
                        }
               };
      end

      err_prefix: begin
        err = '{ valid: 1'b 1,
                 code:  ErrIncorrectFunctionName,
                 info:  { 5'h 0,
                          {err_swsequence, err_modestrength, err_prefix},
                          16'h 0000
                        }
               };
      end

      err_entropy_ready: begin
        err = '{ valid: 1'b 1,
                 code:  ErrSwHashingWithoutEntropyReady,
                 info:  { 8'({ err_entropy_ready,
                               err_swsequence,
                               err_modestrength,
                               err_prefix}),
                          16'({kmac_en_i, cfg_entropy_ready})
                        }
               };
      end

      default: begin
        err = '{valid: 1'b0, code: ErrNone, info: '0};
      end
    endcase
  end : err_return

  assign error_o = err;

  // If below failed, revise err_swsequence error response info field.
  `ASSERT_INIT(ExpectedStSwCmdBits_A, $bits(st) == StateWidth && $bits(sw_cmd_i) == 6)

  // If failed, revise err_modestrength error info field.
  `ASSERT_INIT(ExpectedModeStrengthBits_A,
               $bits(cfg_mode_i) == 2 && $bits(cfg_strength_i) == 3)


  ///////////////////
  // State Machine //
  ///////////////////
  st_e st_gated_d;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, st_gated_d, st, st_e, StIdle)

  // ICEBOX(#14631): Move block_swcmd to PRIM_FLOP_SPARSE_FSM()
  //
  // It would be better to place this condition (block_swcmd) in `always_ff`
  // block to clearly indicate the clock gating condition. However, the
  // statemachine uses the sparse encoding scheme and macro. It prevents any
  // latch enable signals.
  assign st_gated_d = (block_swcmd) ? st : st_d ;

  always_comb begin : next_state
    st_d = st;

    unique case (st)
      StIdle: begin
        if (!app_active_i && sw_cmd_i == CmdStart) begin
          // Proceed to the next state only when the SW issues the Start command
          // in a valid period.
          st_d = StMsgFeed;
        end
      end

      StMsgFeed: begin
        if (sw_cmd_i == CmdProcess) begin
          st_d = StProcessing;
        end
      end

      StProcessing: begin
        if (prim_mubi_pkg::mubi4_test_true_strict(sha3_absorbed_i)) begin
          st_d = StAbsorbed;
        end
      end

      StAbsorbed: begin
        if (sw_cmd_i == CmdManualRun) begin
          st_d = StSqueezing;
        end else if (sw_cmd_i == CmdDone) begin
          st_d = StIdle;
        end
      end

      StSqueezing: begin
        if (keccak_done_i) begin
          st_d = StAbsorbed;
        end
      end

      StTerminalError: begin
        // this state is terminal
        st_d = st;
      end

      default: begin
        // this state is terminal
        st_d = StTerminalError;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en_i != lc_ctrl_pkg::Off) begin
      st_d = StTerminalError;
    end
  end : next_state
  `ASSERT_KNOWN(StKnown_A, st)

endmodule : kmac_errchk


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// KMAC/SHA3

`include "prim_assert.sv"

module kmac
  import kmac_pkg::*;
  import kmac_reg_pkg::*;
#(
  // EnMasking: Enable masking security hardening inside keccak_round
  // If it is enabled, the result digest will be two set of 1600bit.
  parameter bit EnMasking = 1,

  // In case EnMasking == 0, this defines whether SW can provide a masked key or whether Share 1 of
  // the SW key is simply ignored. In case EnMasking == 1, this parameter has no meaning, always
  // both shares of the key provided by SW are used.
  // This is useful to allow both for area-optimized unmasked designs as well as unmasked designs
  // having a SW interface fully compatible with the masked design.
  parameter bit SwKeyMasked = 0,

  // Command delay, useful for SCA measurements only. A value of e.g. 40 allows the processor to go
  // into sleep before KMAC starts operation. If a value > 0 is chosen, the processor can provide
  // two commands subsquently and then go to sleep. The second command is buffered internally and
  // will be presented to the hardware SecCmdDelay number of cycles after the first one.
  parameter int SecCmdDelay = 0,

  // Accept SW message when idle and before receiving a START command. Useful for SCA only.
  parameter bit SecIdleAcceptSwMsg = 1'b0,

  parameter lfsr_perm_t RndCnstLfsrPerm = RndCnstLfsrPermDefault,
  parameter lfsr_seed_t RndCnstLfsrSeed = RndCnstLfsrSeedDefault,
  parameter lfsr_fwd_perm_t RndCnstLfsrFwdPerm = RndCnstLfsrFwdPermDefault,
  parameter msg_perm_t  RndCnstMsgPerm  = RndCnstMsgPermDefault,

  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}}
) (
  input clk_i,
  input rst_ni,

  input rst_shadowed_ni,

  input clk_edn_i,
  input rst_edn_ni,

  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // KeyMgr sideload (secret key) interface
  input keymgr_pkg::hw_key_req_t keymgr_key_i,

  // KeyMgr KDF data path
  input  app_req_t [NumAppIntf-1:0] app_i,
  output app_rsp_t [NumAppIntf-1:0] app_o,

  // EDN interface
  output edn_pkg::edn_req_t entropy_o,
  input  edn_pkg::edn_rsp_t entropy_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t lc_escalate_en_i,

  // interrupts
  output logic intr_kmac_done_o,
  output logic intr_fifo_empty_o,
  output logic intr_kmac_err_o,

  // parameter consistency check with keymgr
  output logic en_masking_o,

  // Idle signal
  output prim_mubi_pkg::mubi4_t idle_o
);

  ////////////////
  // Parameters //
  ////////////////
  localparam int Share = (EnMasking) ? 2 : 1 ;
  localparam int SwKeyShare = (EnMasking || SwKeyMasked) ? 2 : 1;

  /////////////////
  // Definitions //
  /////////////////
  // This state machine is to track the current process based on SW input and
  // KMAC operation.
  // Encoding generated with:
  // $ ./util/design/sparse-fsm-encode.py -d 3 -m 6 -n 6 \
  //      -s 1966361510 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (53.33%)
  //  4: ||||||||||||||| (40.00%)
  //  5: || (6.67%)
  //  6: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 5
  // Minimum Hamming weight: 2
  // Maximum Hamming weight: 5
  //
  localparam int StateWidth = 6;
  typedef enum logic [StateWidth-1:0] {
    // Idle state
    KmacIdle = 6'b001011,

    // When software writes CmdStart @ KmacIdle and kmac_en, FSM moves to this
    KmacPrefix = 6'b000110,

    // When SHA3 engine processes Key block, FSM moves to here.
    KmacKeyBlock = 6'b111110,

    // Message Feed
    KmacMsgFeed = 6'b010101,

    // Complete and squeeze
    KmacDigest = 6'b101101,

    // Error
    KmacTerminalError = 6'b110000

  } kmac_st_e;

  kmac_st_e kmac_st, kmac_st_d;

  /////////////
  // Signals //
  /////////////
  kmac_reg2hw_t reg2hw;
  kmac_hw2reg_t hw2reg;

  // devmode ties to 1 as KMAC should be operated at the beginning for ROM_CTRL.
  logic devmode;
  assign devmode = 1'b 1;

  // Window
  typedef enum int {
    WinState   = 0,
    WinMsgFifo = 1
  } tl_window_e;

  tlul_pkg::tl_h2d_t tl_win_h2d[2];
  tlul_pkg::tl_d2h_t tl_win_d2h[2];

  // SHA3 core control signals and its response.
  // Sequence: start --> process(multiple) --> get absorbed event --> {run -->} done
  logic sha3_start, sha3_run, unused_sha3_squeeze;
  prim_mubi_pkg::mubi4_t sha3_done;
  prim_mubi_pkg::mubi4_t sha3_done_d;
  prim_mubi_pkg::mubi4_t sha3_absorbed;

  // Indicate one block processed
  logic sha3_block_processed;

  // EStatus for entropy
  logic entropy_in_keyblock;

  // Application interface logic generates absorbed from sha3_absorbed.
  // It is active only if SW initiates the hashing engine.
  prim_mubi_pkg::mubi4_t app_absorbed;
  logic event_absorbed;

  sha3_pkg::sha3_st_e sha3_fsm;

  // Prefix: kmac_pkg defines Prefix based on N size and S size.
  // Then computes left_encode(len(N)) size and left_encode(len(S))
  // For given default value 32, 256 bits, the max
  // encode_string(N) || encode_string(S) is 328. So 11 Prefix registers are
  // created.
  logic [sha3_pkg::NSRegisterSize*8-1:0] reg_ns_prefix;
  logic [sha3_pkg::NSRegisterSize*8-1:0] ns_prefix;

  // NumWordsPrefix from kmac_reg_pkg
  `ASSERT_INIT(PrefixRegSameToPrefixPkg_A,
               kmac_reg_pkg::NumWordsPrefix*4 == sha3_pkg::NSRegisterSize)

  // NumEntriesMsgFifo from kmac_reg_pkg must match calculated MsgFifoDepth
  // from kmac_pkg.
  `ASSERT_INIT(NumEntriesRegSameToNumEntriesPkg_A,
               kmac_reg_pkg::NumEntriesMsgFifo == kmac_pkg::MsgFifoDepth)

  // NumBytesMsgFifoEntry from kmac_reg_pkg must match the MsgWidth calculated
  // in kmac_pkg (although MsgWidth is in bits, so we multiply by 8).
  `ASSERT_INIT(EntrySizeRegSameToEntrySizePkg_A,
               kmac_reg_pkg::NumBytesMsgFifoEntry * 8 == kmac_pkg::MsgWidth)

  // Output state: this is used to redirect the digest to KeyMgr or Software
  // depends on the configuration.
  logic state_valid;
  logic [sha3_pkg::StateW-1:0] state [Share];

  // state is de-muxed in keymgr interface logic.
  // the output from keymgr logic goes into staterd module to be visible to SW
  logic reg_state_valid;
  logic [sha3_pkg::StateW-1:0] reg_state [Share];

  // SHA3 Entropy interface
  logic sha3_rand_valid, sha3_rand_early, sha3_rand_consumed;
  logic [sha3_pkg::StateW/2-1:0] sha3_rand_data;
  logic sha3_rand_aux;

  // FIFO related signals
  logic msgfifo_empty, msgfifo_full;
  logic [kmac_pkg::MsgFifoDepthW-1:0] msgfifo_depth;

  logic                          msgfifo_valid       ;
  logic [kmac_pkg::MsgWidth-1:0] msgfifo_data [Share];
  logic [kmac_pkg::MsgStrbW-1:0] msgfifo_strb        ;
  logic                          msgfifo_ready       ;

  if (EnMasking) begin : gen_msgfifo_data_masked
    // In Masked mode, the input message data is split into two shares.
    // Only concern, however, here is the secret key. So message can be
    // put into only one share and other is 0.
    assign msgfifo_data[1] = '0;
  end

  // TL-UL Adapter(MSG_FIFO) signals
  logic        tlram_req;
  logic        tlram_gnt;
  logic        tlram_we;
  logic [8:0]  tlram_addr;   // NOT_READ
  logic [31:0] tlram_wdata;
  logic [31:0] tlram_wmask;
  logic [31:0] tlram_rdata;
  logic        tlram_rvalid;
  logic [1:0]  tlram_rerror;
  logic [31:0] tlram_wdata_endian;
  logic [31:0] tlram_wmask_endian;

  logic                          sw_msg_valid;
  logic [kmac_pkg::MsgWidth-1:0] sw_msg_data ;
  logic [kmac_pkg::MsgWidth-1:0] sw_msg_mask ;
  logic                          sw_msg_ready;

  // KeyMgr interface to MSG_FIFO
  logic                          mux2fifo_valid;
  logic [kmac_pkg::MsgWidth-1:0] mux2fifo_data ;
  logic [kmac_pkg::MsgWidth-1:0] mux2fifo_mask ;
  logic                          mux2fifo_ready;

  // KMAC to SHA3 core
  logic                          msg_valid       ;
  logic [kmac_pkg::MsgWidth-1:0] msg_data [Share];
  logic [kmac_pkg::MsgWidth-1:0] msg_data_masked [Share];
  logic [kmac_pkg::MsgStrbW-1:0] msg_strb        ;
  logic                          msg_ready       ;

  // Process control signals
  // Process pulse propagates from register to SHA3 engine one by one.
  // Each module (MSG_FIFO, KMAC core, SHA3 core) generates the process pulse
  // after flushing internal data to the next module.
  logic reg2msgfifo_process, msgfifo2kmac_process, kmac2sha3_process;


  // Secret Key signals
  logic [MaxKeyLen-1:0] sw_key_data_reg [SwKeyShare];
  logic [MaxKeyLen-1:0] sw_key_data [Share];
  key_len_e             sw_key_len;
  logic [MaxKeyLen-1:0] key_data [Share];
  key_len_e             key_len;

  // SHA3 Mode, Strength, KMAC enable for app interface
  logic                       reg_kmac_en,         app_kmac_en;
  sha3_pkg::sha3_mode_e       reg_sha3_mode,       app_sha3_mode;
  sha3_pkg::keccak_strength_e reg_keccak_strength, app_keccak_strength;

  // RegIF of enabling unsupported mode & strength
  logic cfg_en_unsupported_modestrength;

  // Indicating AppIntf is active. This signal is used to check SW error
  logic app_active;

  // Command
  // sw_cmd is the command written by SW
  // checked_sw_cmd is checked in the kmac_errchk module.
  //   Invalid command is filtered out in the module.
  // kmac_cmd is generated in KeyMgr interface.
  // If SW initiates the KMAC/SHA3, kmac_cmd represents SW command,
  // if KeyMgr drives the data, kmac_cmd is controled in the state machine
  // in KeyMgr interface logic.
  kmac_cmd_e sw_cmd, checked_sw_cmd, kmac_cmd, cmd_q;
  logic      cmd_update;

  // Entropy configurations
  logic [9:0]  wait_timer_prescaler;
  logic [15:0] wait_timer_limit;
  logic        entropy_refresh_req;
  logic [NumSeedsEntropyLfsr-1:0]       entropy_seed_update;
  logic [NumSeedsEntropyLfsr-1:0][31:0] entropy_seed_data;

  logic [HashCntW-1:0] entropy_hash_threshold;
  logic [HashCntW-1:0] entropy_hash_cnt;
  logic                entropy_hash_clr;

  logic entropy_ready;
  entropy_mode_e entropy_mode;
  logic entropy_fast_process;

  prim_mubi_pkg::mubi4_t entropy_configured;

  // Message Masking
  logic msg_mask_en, cfg_msg_mask;
  logic [MsgWidth-1:0] msg_mask;

  // SHA3 Error response
  sha3_pkg::err_t sha3_err;

  // KeyMgr Error response
  kmac_pkg::err_t app_err;

  // Entropy Generator Error
  kmac_pkg::err_t entropy_err;

  // Error checker
  kmac_pkg::err_t errchecker_err;

  // MsgFIFO Error
  kmac_pkg::err_t msgfifo_err;

  logic err_processed;

  logic alert_fatal, alert_recov_operation;
  logic alert_intg_err;

  // Life cycle
  localparam int unsigned NumLcSyncCopies = 6;
  lc_ctrl_pkg::lc_tx_t [NumLcSyncCopies-1:0] lc_escalate_en_sync;
  lc_ctrl_pkg::lc_tx_t [NumLcSyncCopies-1:0] lc_escalate_en;

  //////////////////////////////////////
  // Connecting Register IF to logics //
  //////////////////////////////////////

  // Function-name N and Customization input string S
  always_comb begin
    for (int i = 0 ; i < NumWordsPrefix; i++) begin
      reg_ns_prefix[32*i+:32] = reg2hw.prefix[i].q;
    end
  end

  // Create a lint error to reduce the risk of accidentally enabling this feature.
  `ASSERT_STATIC_LINT_ERROR(KmacSecCmdDelayNonDefault, SecCmdDelay == 0)

  if (SecCmdDelay > 0) begin : gen_cmd_delay_buf
    // Delay and buffer commands for SCA measurements.
    localparam int unsigned WidthCounter = $clog2(SecCmdDelay+1);
    logic [WidthCounter-1:0] count_d, count_q;
    logic                    counting_d, counting_q;
    logic                    cmd_buf_empty;
    kmac_cmd_e               cmd_buf_q;

    assign cmd_buf_empty = (cmd_buf_q == CmdNone);

    // When seeing a write to the cmd register, we start counting. We stop counting once the
    // counter has expired and the command buffer is empty.
    assign counting_d = reg2hw.cmd.cmd.qe          ? 1'b1 :
                        cmd_update & cmd_buf_empty ? 1'b0 : counting_q;

    // Clear counter upon writes to the cmd register or if the specified delay is reached.
    assign count_d = reg2hw.cmd.cmd.qe ? '0             :
                     cmd_update        ? '0             :
                     counting_q        ? count_q + 1'b1 : count_q;

    // The manual run command cannot be delayed. Software expects this to be triggered immediately
    // and will poll the status register to wait for the SHA3 engine to return back to the squeeze
    // state.
    assign cmd_update = (cmd_q == CmdManualRun)                    ? 1'b1 :
                        (count_q == SecCmdDelay[WidthCounter-1:0]) ? 1'b1 : 1'b0;

    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        count_q    <= '0;
        counting_q <= 1'b0;
      end else begin
        count_q    <= count_d;
        counting_q <= counting_d;
      end
    end

    // cmd.q is valid while cmd.qe is high, meaning it needs to be registered. We buffer one
    // additional command such that software can write START followed by PROCESS and then go to
    // sleep.
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        cmd_q     <= CmdNone;
        cmd_buf_q <= CmdNone;
      end else begin
        if (reg2hw.cmd.cmd.qe && cmd_update) begin
          // New write & counter expired.
          cmd_q     <= cmd_buf_q;
          cmd_buf_q <= kmac_cmd_e'(reg2hw.cmd.cmd.q);

        end else if (reg2hw.cmd.cmd.qe) begin
          // New write.
          if (counting_q == 1'b0) begin
            cmd_q     <= kmac_cmd_e'(reg2hw.cmd.cmd.q);
          end else begin
            cmd_buf_q <= kmac_cmd_e'(reg2hw.cmd.cmd.q);
          end

        end else if (cmd_update) begin
          // Counter expired.
          cmd_q     <= cmd_buf_q;
          cmd_buf_q <= CmdNone;
        end
      end
    end

  end else begin : gen_no_cmd_delay_buf
    // Directly forward signals from register IF.
    assign cmd_update = reg2hw.cmd.cmd.qe;
    assign cmd_q      = kmac_cmd_e'(reg2hw.cmd.cmd.q);
  end

  // Command signals
  assign sw_cmd = (cmd_update) ? cmd_q : CmdNone;
  `ASSERT_KNOWN(KmacCmd_A, sw_cmd)
  always_comb begin
    sha3_start = 1'b 0;
    sha3_run = 1'b 0;
    sha3_done_d = prim_mubi_pkg::MuBi4False;
    reg2msgfifo_process = 1'b 0;

    unique case (kmac_cmd)
      CmdStart: begin
        sha3_start = 1'b 1;
      end

      CmdProcess: begin
        reg2msgfifo_process = 1'b 1;
      end

      CmdManualRun: begin
        sha3_run = 1'b 1;
      end

      CmdDone: begin
        sha3_done_d = prim_mubi_pkg::MuBi4True;
      end

      CmdNone: begin
        // inactive state
      end

      default: begin
      end
    endcase
  end

  // Status register ==========================================================
  // status.squeeze is valid only when SHA3 engine completes the Absorb and not
  // running the manual keccak rounds. This status is for SW to determine when
  // to read the STATE values.
  assign hw2reg.status.sha3_idle.d     = sha3_fsm == sha3_pkg::StIdle;
  assign hw2reg.status.sha3_absorb.d   = sha3_fsm == sha3_pkg::StAbsorb;
  assign hw2reg.status.sha3_squeeze.d  = sha3_fsm == sha3_pkg::StSqueeze;

  // FIFO related status
  assign hw2reg.status.fifo_depth.d[MsgFifoDepthW-1:0] = msgfifo_depth;
  if ($bits(hw2reg.status.fifo_depth.d) != MsgFifoDepthW) begin : gen_fifo_depth_tie
    assign hw2reg.status.fifo_depth.d[$bits(hw2reg.status.fifo_depth.d)-1:MsgFifoDepthW] = '0;
  end
  assign hw2reg.status.fifo_empty.d  = msgfifo_empty;
  assign hw2reg.status.fifo_full.d   = msgfifo_full;

  // Configuration Register
  logic engine_stable;
  assign engine_stable = sha3_fsm == sha3_pkg::StIdle;

  // SEC_CM: CFG_SHADOWED.CONFIG.REGWEN
  assign hw2reg.cfg_regwen.d = engine_stable;

  // Secret Key
  // Secret key is defined as external register. So the logic latches when SW
  // writes to KEY_SHARE0 , KEY_SHARE1 registers.
  // SEC_CM: SW_KEY.KEY.MASKING
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      sw_key_data_reg[0] <= '0;
    end else if (engine_stable) begin
      for (int j = 0 ; j < MaxKeyLen/32 ; j++) begin
        if (reg2hw.key_share0[j].qe) begin
          sw_key_data_reg[0][32*j+:32] <= reg2hw.key_share0[j].q;
        end
      end // for j
    end // else if engine_stable
  end // always_ff

  if (EnMasking || SwKeyMasked) begin : gen_key_share1_reg
    always_ff @(posedge clk_i or negedge rst_ni) begin
      if (!rst_ni) begin
        sw_key_data_reg[1] <= '0;
      end else if (engine_stable) begin
        for (int j = 0 ; j < MaxKeyLen/32 ; j++) begin
          if (reg2hw.key_share1[j].qe) begin
            sw_key_data_reg[1][32*j+:32] <= reg2hw.key_share1[j].q;
          end
        end // for j
      end // else if engine_stable
    end // always_ff
  end else begin : gen_no_key_share1_reg
    logic unused_key_share1;
    assign unused_key_share1 = ^reg2hw.key_share1;
  end

  if (EnMasking || !SwKeyMasked) begin : gen_key_forward
    // Forward all available key shares as is.
    assign sw_key_data = sw_key_data_reg;
  end else begin : gen_key_unmask
    // Masking is disabled but the SW still provides the key in two shares.
    // Unmask the key for processing.
    assign sw_key_data[0] = sw_key_data_reg[0] ^ sw_key_data_reg[1];
  end

  assign sw_key_len = key_len_e'(reg2hw.key_len.q);

  // Entropy configurations
  assign wait_timer_prescaler = reg2hw.entropy_period.prescaler.q;
  assign wait_timer_limit     = reg2hw.entropy_period.wait_timer.q;
  assign entropy_refresh_req = reg2hw.cmd.entropy_req.q
                            && reg2hw.cmd.entropy_req.qe;
  for (genvar i = 0; i < NumSeedsEntropyLfsr; i++) begin : gen_entropy_seed
    assign entropy_seed_update[i] = reg2hw.entropy_seed[i].qe;
    assign entropy_seed_data[i] = reg2hw.entropy_seed[i].q;
  end

  assign entropy_hash_threshold = reg2hw.entropy_refresh_threshold_shadowed.q;
  assign hw2reg.entropy_refresh_hash_cnt.de = 1'b 1;
  assign hw2reg.entropy_refresh_hash_cnt.d  = entropy_hash_cnt;

  assign entropy_hash_clr = reg2hw.cmd.hash_cnt_clr.qe
                         && reg2hw.cmd.hash_cnt_clr.q;

  // Entropy config
  assign entropy_ready = reg2hw.cfg_shadowed.entropy_ready.q
                       & reg2hw.cfg_shadowed.entropy_ready.qe;
  assign entropy_mode  = entropy_mode_e'(reg2hw.cfg_shadowed.entropy_mode.q);
  assign entropy_fast_process = reg2hw.cfg_shadowed.entropy_fast_process.q;

  // msg_mask_en turns on the message LFSR when KMAC is enabled.
  assign cfg_msg_mask = reg2hw.cfg_shadowed.msg_mask.q;
  assign msg_mask_en = cfg_msg_mask & msg_valid & msg_ready;

  // Enable unsupported mode & strength combination
  assign cfg_en_unsupported_modestrength =
    reg2hw.cfg_shadowed.en_unsupported_modestrength.q;

  `ASSERT(EntropyReadyLatched_A, $rose(entropy_ready) |=> !entropy_ready)

  // Idle control (registered output)
  // The logic checks idle of SHA3 engine, MSG_FIFO, KMAC_CORE, KEYMGR interface
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      idle_o <= prim_mubi_pkg::MuBi4True;
    end else if ((sha3_fsm == sha3_pkg::StIdle) && (msgfifo_empty || SecIdleAcceptSwMsg)) begin
      idle_o <= prim_mubi_pkg::MuBi4True;
    end else begin
      idle_o <= prim_mubi_pkg::MuBi4False;
    end
  end

  // Clear the error processed
  assign err_processed = reg2hw.cfg_shadowed.err_processed.q
                       & reg2hw.cfg_shadowed.err_processed.qe;

  // Make sure the field has latch in reg_top
  `ASSERT(ErrProcessedLatched_A, $rose(err_processed) |=> !err_processed)

  // App mode, strength, kmac_en
  assign reg_kmac_en         = reg2hw.cfg_shadowed.kmac_en.q;
  assign reg_sha3_mode       = sha3_pkg::sha3_mode_e'(reg2hw.cfg_shadowed.mode.q);
  assign reg_keccak_strength = sha3_pkg::keccak_strength_e'(reg2hw.cfg_shadowed.kstrength.q);

  ///////////////
  // Interrupt //
  ///////////////

  logic event_msgfifo_empty, msgfifo_empty_q;

  // Hash process absorbed interrupt
  // Convert mubi4_t to logic to generate interrupts
  assign event_absorbed = prim_mubi_pkg::mubi4_test_true_strict(app_absorbed);

  prim_intr_hw #(.Width(1)) intr_kmac_done (
    .clk_i,
    .rst_ni,
    .event_intr_i           (event_absorbed),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.kmac_done.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.kmac_done.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.kmac_done.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.kmac_done.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.kmac_done.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.kmac_done.d),
    .intr_o                 (intr_kmac_done_o)
  );

  `ASSERT(Sha3AbsorbedPulse_A,
    $rose(prim_mubi_pkg::mubi4_test_true_strict(sha3_absorbed)) |=>
      prim_mubi_pkg::mubi4_test_false_strict(sha3_absorbed))

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) msgfifo_empty_q <= 1'b1;
    else         msgfifo_empty_q <= msgfifo_empty;
  end

  assign event_msgfifo_empty = ~msgfifo_empty_q & msgfifo_empty;

  prim_intr_hw #(.Width(1)) intr_fifo_empty (
    .clk_i,
    .rst_ni,
    .event_intr_i           (event_msgfifo_empty),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.fifo_empty.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.fifo_empty.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.fifo_empty.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.fifo_empty.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.fifo_empty.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.fifo_empty.d),
    .intr_o                 (intr_fifo_empty_o)
  );

  // Error
  // As of now, only SHA3 error exists. More error codes will be added.

  logic event_error;
  assign event_error = sha3_err.valid    | app_err.valid
                     | entropy_err.valid | errchecker_err.valid
                     ;

  // Assing error code to the register
  assign hw2reg.err_code.de = event_error;

  always_comb begin
    hw2reg.err_code.d = '0;

    priority case (1'b 1)
      // app_err has the highest priority. If SW issues an incorrect command
      // while app is in active state, the error from AppIntf is passed
      // through.
      app_err.valid: begin
        hw2reg.err_code.d = {app_err.code, app_err.info};
      end

      errchecker_err.valid: begin
        hw2reg.err_code.d = {errchecker_err.code , errchecker_err.info};
      end

      sha3_err.valid: begin
        hw2reg.err_code.d = {sha3_err.code , sha3_err.info};
      end

      entropy_err.valid: begin
        hw2reg.err_code.d = {entropy_err.code, entropy_err.info};
      end

      msgfifo_err.valid: begin
        hw2reg.err_code.d = {msgfifo_err.code, msgfifo_err.info};
      end

      default: begin
        hw2reg.err_code.d = '0;
      end
    endcase
  end

  // Counter errors
  logic counter_error, sha3_count_error, key_index_error;
  logic msgfifo_counter_error;
  logic kmac_entropy_hash_counter_error;
  assign counter_error = sha3_count_error
                       | kmac_entropy_hash_counter_error
                       | key_index_error
                       | msgfifo_counter_error;

  assign msgfifo_counter_error = msgfifo_err.valid;

  // State Errors
  logic sparse_fsm_error;
  logic sha3_state_error, kmac_errchk_state_error;
  logic kmac_core_state_error, kmac_app_state_error;
  logic kmac_entropy_state_error, kmac_state_error;
  assign sparse_fsm_error = sha3_state_error
                          | kmac_errchk_state_error
                          | kmac_core_state_error
                          | kmac_app_state_error
                          | kmac_entropy_state_error
                          | kmac_state_error;

  // Control Signal Integrity Errors
  logic control_integrity_error;
  logic sha3_storage_rst_error;
  assign control_integrity_error = sha3_storage_rst_error;

  prim_intr_hw #(.Width(1)) intr_kmac_err (
    .clk_i,
    .rst_ni,
    .event_intr_i           (event_error),
    .reg2hw_intr_enable_q_i (reg2hw.intr_enable.kmac_err.q),
    .reg2hw_intr_test_q_i   (reg2hw.intr_test.kmac_err.q),
    .reg2hw_intr_test_qe_i  (reg2hw.intr_test.kmac_err.qe),
    .reg2hw_intr_state_q_i  (reg2hw.intr_state.kmac_err.q),
    .hw2reg_intr_state_de_o (hw2reg.intr_state.kmac_err.de),
    .hw2reg_intr_state_d_o  (hw2reg.intr_state.kmac_err.d),
    .intr_o                 (intr_kmac_err_o)
  );

  ///////////////////
  // State Machine //
  ///////////////////

  // State FF
  `PRIM_FLOP_SPARSE_FSM(u_state_regs, kmac_st_d, kmac_st, kmac_st_e, KmacIdle)

  always_comb begin
    // Default value
    kmac_st_d = kmac_st;

    entropy_in_keyblock = 1'b 0;
    kmac_state_error = 1'b 0;

    unique case (kmac_st)
      KmacIdle: begin
        if (kmac_cmd == CmdStart) begin
          // If cSHAKE turned on
          if (sha3_pkg::CShake == app_sha3_mode) begin
            kmac_st_d = KmacPrefix;
          end else begin
            // Jump to Msg feed directly
            kmac_st_d = KmacMsgFeed;
          end
        end else begin
          kmac_st_d = KmacIdle;
        end
      end

      KmacPrefix: begin
        // Wait until SHA3 processes one block
        if (sha3_block_processed) begin
          kmac_st_d = (app_kmac_en) ? KmacKeyBlock : KmacMsgFeed ;
        end else begin
          kmac_st_d = KmacPrefix;
        end
      end

      KmacKeyBlock: begin
        entropy_in_keyblock = 1'b 1;
        if (sha3_block_processed) begin
          kmac_st_d = KmacMsgFeed;
        end else begin
          kmac_st_d = KmacKeyBlock;
        end
      end

      KmacMsgFeed: begin
        // If absorbed, move to Digest
        if (prim_mubi_pkg::mubi4_test_true_strict(sha3_absorbed) &&
          prim_mubi_pkg::mubi4_test_true_strict(sha3_done)) begin
          // absorbed and done can be asserted at a cycle if Applications have
          // requested the hash operation. kmac_app FSM issues CmdDone command
          // if it receives absorbed signal.
          kmac_st_d = KmacIdle;
        end else if (prim_mubi_pkg::mubi4_test_true_strict(sha3_absorbed) &&
          prim_mubi_pkg::mubi4_test_false_loose(sha3_done)) begin
          kmac_st_d = KmacDigest;
        end else begin
          kmac_st_d = KmacMsgFeed;
        end
      end

      KmacDigest: begin
        // SW can manually run it, wait till done
        if (prim_mubi_pkg::mubi4_test_true_strict(sha3_done)) begin
          kmac_st_d = KmacIdle;
        end else begin
          kmac_st_d = KmacDigest;
        end
      end

      KmacTerminalError: begin
        //this state is terminal
        kmac_st_d = KmacTerminalError;
        kmac_state_error = 1'b 1;
      end

      default: begin
        kmac_st_d = KmacTerminalError;
        kmac_state_error = 1'b 1;
      end
    endcase

    // SEC_CM: FSM.GLOBAL_ESC, FSM.LOCAL_ESC
    // Unconditionally jump into the terminal error state
    // if the life cycle controller triggers an escalation.
    if (lc_escalate_en[0] != lc_ctrl_pkg::Off) begin
      kmac_st_d = KmacTerminalError;
    end
  end
  `ASSERT_KNOWN(KmacStKnown_A, kmac_st)

  ///////////////
  // Instances //
  ///////////////

  // KMAC core
  kmac_core #(
    .EnMasking (EnMasking)
  ) u_kmac_core (
    .clk_i,
    .rst_ni,

    // from Msg FIFO
    .fifo_valid_i (msgfifo_valid),
    .fifo_data_i  (msgfifo_data ),
    .fifo_strb_i  (msgfifo_strb ),
    .fifo_ready_o (msgfifo_ready),

    // to SHA3 core
    .msg_valid_o  (msg_valid),
    .msg_data_o   (msg_data ),
    .msg_strb_o   (msg_strb ),
    .msg_ready_i  (msg_ready),

    // Configurations
    .kmac_en_i  (app_kmac_en),
    .mode_i     (app_sha3_mode),
    .strength_i (app_keccak_strength),

    // Secret key interface
    .key_data_i (key_data),
    .key_len_i  (key_len ),

    // Controls
    .start_i   (sha3_start          ),
    .process_i (msgfifo2kmac_process),
    .done_i    (sha3_done           ),
    .process_o (kmac2sha3_process   ),

    // LC escalation
    .lc_escalate_en_i (lc_escalate_en[1]),

    // Error detection
    .sparse_fsm_error_o (kmac_core_state_error),
    .key_index_error_o  (key_index_error)
  );

  // SHA3 hashing engine

  // msg_data masking
  if (EnMasking == 1) begin: g_msg_mask
    logic [MsgWidth-1:0] msg_mask_permuted;

    // Permute the LFSR output to avoid same lfsr applied to multiple times
    always_comb begin
      msg_mask_permuted = '0;
      for (int unsigned i = 0 ; i < MsgWidth ; i++) begin
        // Loop through the MsgPerm constant and swap between the bits
        msg_mask_permuted[i] = msg_mask[RndCnstMsgPerm[i]];
      end
    end

    for (genvar i = 0 ; i < Share ; i++) begin: g_msg_data_mask
      assign msg_data_masked[i] = msg_data[i]
                                ^ ({MsgWidth{cfg_msg_mask}} & msg_mask_permuted);
    end : g_msg_data_mask
  end else begin : g_no_msg_mask
    assign msg_data_masked[0] = msg_data[0];

    logic unused_msgmask;
    assign unused_msgmask = ^{msg_mask, cfg_msg_mask, msg_mask_en};
  end
  sha3 #(
    .EnMasking (EnMasking)
  ) u_sha3 (
    .clk_i,
    .rst_ni,

    // MSG_FIFO interface (or from KMAC)
    .msg_valid_i (msg_valid),
    .msg_data_i  (msg_data_masked ),
    .msg_strb_i  (msg_strb ),
    .msg_ready_o (msg_ready),

    // Entropy interface
    .rand_valid_i    (sha3_rand_valid),
    .rand_early_i    (sha3_rand_early),
    .rand_data_i     (sha3_rand_data),
    .rand_aux_i      (sha3_rand_aux),
    .rand_consumed_o (sha3_rand_consumed),

    // N, S: Used in cSHAKE mode
    .ns_data_i       (ns_prefix),

    // Configurations
    .mode_i     (app_sha3_mode),
    .strength_i (app_keccak_strength),

    // Controls (CMD register)
    .start_i    (sha3_start       ),
    .process_i  (kmac2sha3_process),
    .run_i      (sha3_run         ),
    .done_i     (sha3_done        ),

    // LC escalation
    .lc_escalate_en_i (lc_escalate_en[2]),

    .absorbed_o  (sha3_absorbed),
    .squeezing_o (unused_sha3_squeeze),

    .block_processed_o (sha3_block_processed),

    .sha3_fsm_o (sha3_fsm),

    .state_valid_o (state_valid),
    .state_o       (state), // [Share]

    .error_o                    (sha3_err),
    .sparse_fsm_error_o         (sha3_state_error),
    .count_error_o              (sha3_count_error),
    .keccak_storage_rst_error_o (sha3_storage_rst_error)
  );

  // MSG_FIFO window interface to FIFO interface ===============================
  // Tie the read path
  assign tlram_rvalid = 1'b 0;
  assign tlram_rdata = '0;
  assign tlram_rerror = '0;

  // Convert endian here
  //    prim_packer always packs to the right(bit0). If the input DWORD is
  //    big-endian, it needs to be swapped to little-endian to maintain the
  //    order. Internal SHA3(Keccak) runs in little-endian in contrast to HMAC
  //    So, no endian-swap after prim_packer.
  assign tlram_wdata_endian = conv_endian32(tlram_wdata,
                                reg2hw.cfg_shadowed.msg_endianness.q);
  assign tlram_wmask_endian = conv_endian32(tlram_wmask,
                                reg2hw.cfg_shadowed.msg_endianness.q);

  // TL Adapter
  tlul_adapter_sram #(
    .SramAw ($clog2(MsgWindowDepth)),
    .SramDw (MsgWindowWidth),
    .Outstanding (1),
    .ByteAccess  (1),
    .ErrOnRead   (1)
  ) u_tlul_adapter_msgfifo (
    .clk_i,
    .rst_ni,
    .en_ifetch_i (prim_mubi_pkg::MuBi4False),
    .tl_i        (tl_win_h2d[WinMsgFifo]),
    .tl_o        (tl_win_d2h[WinMsgFifo]),

    .req_o       (tlram_req),
    .req_type_o  (),
    .gnt_i       (tlram_gnt),
    .we_o        (tlram_we ),
    .addr_o      (tlram_addr),
    .wdata_o     (tlram_wdata),
    .wmask_o     (tlram_wmask),
    .intg_error_o(           ),
    .rdata_i     (tlram_rdata),
    .rvalid_i    (tlram_rvalid),
    .rerror_i    (tlram_rerror)
  );

  assign sw_msg_valid = tlram_req & tlram_we ;
  if (MsgWidth == MsgWindowWidth) begin : gen_sw_msg_samewidth
    assign sw_msg_data  = tlram_wdata_endian ;
    assign sw_msg_mask  = tlram_wmask_endian ;
  end else begin : gen_sw_msg_diff
    assign sw_msg_data = {{MsgWidth-MsgWindowWidth{1'b0}}, tlram_wdata_endian};
    assign sw_msg_mask = {{MsgWidth-MsgWindowWidth{1'b0}}, tlram_wmask_endian};
  end
  assign tlram_gnt    = sw_msg_ready ;

  logic unused_tlram_addr;
  assign unused_tlram_addr = &{1'b0, tlram_addr};

  // Application interface Mux/Demux
  kmac_app #(
    .EnMasking(EnMasking),
    .SecIdleAcceptSwMsg(SecIdleAcceptSwMsg)
  ) u_app_intf (
    .clk_i,
    .rst_ni,

    .reg_key_data_i (sw_key_data),
    .reg_key_len_i  (sw_key_len),

    .reg_prefix_i (reg_ns_prefix),

    .reg_kmac_en_i         (reg_kmac_en),
    .reg_sha3_mode_i       (reg_sha3_mode),
    .reg_keccak_strength_i (reg_keccak_strength),

    // data from tl_adapter
    .sw_valid_i (sw_msg_valid),
    .sw_data_i  (sw_msg_data),
    .sw_mask_i  (sw_msg_mask),
    .sw_ready_o (sw_msg_ready),

    // KeyMgr sideloaded key interface
    .keymgr_key_i,

    // Application data in / digest out interface
    .app_i,
    .app_o,

    // Secret Key output to KMAC Core
    .key_data_o (key_data),
    .key_len_o  (key_len),

    // to MSG_FIFO
    .kmac_valid_o (mux2fifo_valid),
    .kmac_data_o  (mux2fifo_data),
    .kmac_mask_o  (mux2fifo_mask),
    .kmac_ready_i (mux2fifo_ready),

    // to KMAC Core
    .kmac_en_o (app_kmac_en),

    // to SHA3 Core
    .sha3_prefix_o     (ns_prefix),
    .sha3_mode_o       (app_sha3_mode),
    .keccak_strength_o (app_keccak_strength),

    // Keccak state from SHA3 core
    .keccak_state_valid_i (state_valid),
    .keccak_state_i       (state),

    // to STATE TL Window
    .reg_state_valid_o    (reg_state_valid),
    .reg_state_o          (reg_state),

    // Configuration: Sideloaded Key
    .keymgr_key_en_i      (reg2hw.cfg_shadowed.sideload.q),

    .absorbed_i (sha3_absorbed), // from SHA3
    .absorbed_o (app_absorbed),  // to SW

    .app_active_o(app_active),

    .error_i         (sha3_err.valid),
    .err_processed_i (err_processed),

    // Command interface
    .sw_cmd_i (checked_sw_cmd),
    .cmd_o    (kmac_cmd),

    // Status
    .entropy_ready_i (entropy_configured),

    // LC escalation
    .lc_escalate_en_i (lc_escalate_en[3]),

    // Error report
    .error_o            (app_err),
    .sparse_fsm_error_o (kmac_app_state_error)

  );

  // Message FIFO
  kmac_msgfifo #(
    .OutWidth  (kmac_pkg::MsgWidth),
    .MsgDepth  (kmac_pkg::MsgFifoDepth),
    .EnMasking (EnMasking)
  ) u_msgfifo (
    .clk_i,
    .rst_ni,

    .fifo_valid_i (mux2fifo_valid),
    .fifo_data_i  (mux2fifo_data),
    .fifo_mask_i  (mux2fifo_mask),
    .fifo_ready_o (mux2fifo_ready),

    .msg_valid_o (msgfifo_valid),
    .msg_data_o  (msgfifo_data[0]),
    .msg_strb_o  (msgfifo_strb),
    .msg_ready_i (msgfifo_ready),

    .fifo_empty_o (msgfifo_empty), // intr and status
    .fifo_full_o  (msgfifo_full),  // connected to status only
    .fifo_depth_o (msgfifo_depth),

    .clear_i (sha3_done),

    .process_i (reg2msgfifo_process ),
    .process_o (msgfifo2kmac_process),

    .err_o (msgfifo_err)
  );

  logic [sha3_pkg::StateW-1:0] reg_state_tl [Share];
  always_comb begin
    for (int i = 0 ; i < Share; i++) begin
      reg_state_tl[i] = reg_state_valid ? reg_state[i] : 'b0;
    end
  end

  // State (Digest) reader
  kmac_staterd #(
    .AddrW     (9), // 512B
    .EnMasking (EnMasking)
  ) u_staterd (
    .clk_i,
    .rst_ni,

    .tl_i (tl_win_h2d[WinState]),
    .tl_o (tl_win_d2h[WinState]),

    .state_i (reg_state_tl),

    .endian_swap_i (reg2hw.cfg_shadowed.state_endianness.q)
  );

  // Error checker
  kmac_errchk #(
    .EnMasking (EnMasking)
  ) u_errchk (
    .clk_i,
    .rst_ni,

    // Configurations
    .cfg_mode_i    (reg_sha3_mode      ),
    .cfg_strength_i(reg_keccak_strength),

    .kmac_en_i      (reg_kmac_en        ),
    .cfg_prefix_6B_i(reg_ns_prefix[47:0]), // first 6B of PREFIX

    .cfg_en_unsupported_modestrength_i (cfg_en_unsupported_modestrength),

    .entropy_ready_pulse_i (entropy_ready),

    // SW commands
    .sw_cmd_i(sw_cmd),
    .sw_cmd_o(checked_sw_cmd),

    // Status from KMAC_APP
    .app_active_i(app_active),

    // Status from SHA3 core
    .sha3_absorbed_i(sha3_absorbed       ),
    .keccak_done_i  (sha3_block_processed),

    // LC escalation
    .lc_escalate_en_i (lc_escalate_en[4]),

    .err_processed_i (err_processed),

    .error_o            (errchecker_err),
    .sparse_fsm_error_o (kmac_errchk_state_error)
  );

  // Entropy Generator
  if (EnMasking == 1) begin : gen_entropy

    logic entropy_req, entropy_ack;
    logic [edn_pkg::ENDPOINT_BUS_WIDTH-1:0] entropy_data;
    logic unused_entropy_fips;

    // Synchronize EDN interface
    prim_sync_reqack_data #(
      .Width(edn_pkg::ENDPOINT_BUS_WIDTH),
      .DataSrc2Dst(1'b0),
      .DataReg(1'b0)
    ) u_prim_sync_reqack_data (
      .clk_src_i (clk_i),
      .rst_src_ni(rst_ni),
      .clk_dst_i (clk_edn_i),
      .rst_dst_ni(rst_edn_ni),
      .req_chk_i ((kmac_entropy_state_error == 1'b0) && (entropy_err.valid == 1'b0)),
      .src_req_i (entropy_req),
      .src_ack_o (entropy_ack),
      .dst_req_o (entropy_o.edn_req),
      .dst_ack_i (entropy_i.edn_ack),
      .data_i    (entropy_i.edn_bus),
      .data_o    (entropy_data)
    );

    // We don't track whether the entropy is pre-FIPS or not inside KMAC.
    assign unused_entropy_fips = entropy_i.edn_fips;

    kmac_entropy #(
     .RndCnstLfsrPerm(RndCnstLfsrPerm),
     .RndCnstLfsrSeed(RndCnstLfsrSeed),
     .RndCnstLfsrFwdPerm(RndCnstLfsrFwdPerm)
    ) u_entropy (
      .clk_i,
      .rst_ni,

      // EDN interface
      .entropy_req_o (entropy_req),
      .entropy_ack_i (entropy_ack),
      .entropy_data_i(entropy_data),

      // Entropy to internal logic (DOM AND)
      .rand_valid_o    (sha3_rand_valid),
      .rand_early_o    (sha3_rand_early),
      .rand_data_o     (sha3_rand_data),
      .rand_aux_o      (sha3_rand_aux),
      .rand_consumed_i (sha3_rand_consumed),

      // Status from internal logic
      //// KMAC secret block handling indicator
      .in_keyblock_i (entropy_in_keyblock),

      // Configuration
      .mode_i          (entropy_mode),
      .entropy_ready_i (entropy_ready),
      .fast_process_i  (entropy_fast_process),

      //// Entropy refresh period in clk cycles
      .wait_timer_prescaler_i (wait_timer_prescaler),
      .wait_timer_limit_i     (wait_timer_limit),

      //// Message Masking
      .msg_mask_en_i (msg_mask_en),
      .msg_mask_o    (msg_mask),

      //// SW update of seed
      .seed_update_i         (entropy_seed_update),
      .seed_data_i           (entropy_seed_data),
      .entropy_refresh_req_i (entropy_refresh_req),

      // Status
      .hash_cnt_o       (entropy_hash_cnt),
      .hash_cnt_clr_i   (entropy_hash_clr),
      .hash_threshold_i (entropy_hash_threshold),

      .entropy_configured_o (entropy_configured),

      // LC escalation
      .lc_escalate_en_i (lc_escalate_en[5]),

      // Error
      .err_o              (entropy_err),
      .sparse_fsm_error_o (kmac_entropy_state_error),
      .count_error_o      (kmac_entropy_hash_counter_error),
      .err_processed_i    (err_processed)
    );
  end else begin : gen_empty_entropy
    // If Masking is not used, no need of entropy. Ignore inputs and config; tie output to 0.
    edn_pkg::edn_rsp_t unused_entropy_input;
    entropy_mode_e     unused_entropy_mode;
    logic              unused_entropy_fast_process;

    assign unused_entropy_input        = entropy_i;
    assign unused_entropy_mode         = entropy_mode;
    assign unused_entropy_fast_process = entropy_fast_process;

    assign entropy_o = '{default: '0};

    logic unused_sha3_rand_consumed;
    assign sha3_rand_valid = 1'b 1;
    assign sha3_rand_early = 1'b 1;
    assign sha3_rand_data = '0;
    assign sha3_rand_aux = '0;
    assign unused_sha3_rand_consumed = sha3_rand_consumed;

    logic [NumSeedsEntropyLfsr-1:0]       unused_seed_update;
    logic [NumSeedsEntropyLfsr-1:0][31:0] unused_seed_data;
    logic [31:0] unused_refresh_period;
    logic unused_entropy_refresh_req;
    assign unused_seed_data = entropy_seed_data;
    assign unused_seed_update = entropy_seed_update;
    assign unused_refresh_period = ^{wait_timer_limit, wait_timer_prescaler};
    assign unused_entropy_refresh_req = entropy_refresh_req;

    logic unused_entropy_hash;
    assign unused_entropy_hash = ^{entropy_hash_clr, entropy_hash_threshold};
    assign entropy_hash_cnt = '0;

    assign entropy_err = '{valid: 1'b 0, code: ErrNone, info: '0};

    assign kmac_entropy_state_error = 1'b 0;
    assign kmac_entropy_hash_counter_error  = 1'b 0;

    logic [1:0] unused_entropy_status;
    assign unused_entropy_status = entropy_in_keyblock;

    // If Masking is off, always entropy configured
    assign entropy_configured = prim_mubi_pkg::MuBi4True;
  end

  // MUBI4 buf
  prim_mubi4_sender #(
    .AsyncOn (0)
  ) u_sha3_done_sender (
    .clk_i,
    .rst_ni,
    .mubi_i (sha3_done_d),
    .mubi_o (sha3_done)
  );

  // Register top
  logic [NumAlerts-1:0] alert_test, alerts, alerts_q;

  logic shadowed_storage_err, shadowed_update_err;
  kmac_reg_top u_reg (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni,

    .tl_i,
    .tl_o,

    .tl_win_o (tl_win_h2d),
    .tl_win_i (tl_win_d2h),

    .reg2hw,
    .hw2reg,

    // SEC_CM: CFG_SHADOWED.CONFIG.SHADOW
    .shadowed_storage_err_o (shadowed_storage_err),
    .shadowed_update_err_o  (shadowed_update_err),
    // SEC_CM: BUS.INTEGRITY
    .intg_err_o             (alert_intg_err),

    .devmode_i (devmode)
  );

  logic unused_cfg_shadowed_qe;
  assign unused_cfg_shadowed_qe = ^{
    reg2hw.cfg_shadowed.kmac_en.qe                     ,
    reg2hw.cfg_shadowed.kstrength.qe                   ,
    reg2hw.cfg_shadowed.mode.qe                        ,
    reg2hw.cfg_shadowed.msg_endianness.qe              ,
    reg2hw.cfg_shadowed.state_endianness.qe            ,
    reg2hw.cfg_shadowed.sideload.qe                    ,
    reg2hw.cfg_shadowed.entropy_mode.qe                ,
    reg2hw.cfg_shadowed.entropy_fast_process.qe        ,
    reg2hw.cfg_shadowed.msg_mask.qe                    ,
    reg2hw.cfg_shadowed.en_unsupported_modestrength.qe
    };

  // Alerts
  assign alert_test = {
    reg2hw.alert_test.fatal_fault_err.q
      & reg2hw.alert_test.fatal_fault_err.qe,    // [1]
    reg2hw.alert_test.recov_operation_err.q
      & reg2hw.alert_test.recov_operation_err.qe // [0]
  };

  assign alerts = {
    alert_fatal,           // Alerts[1]
    alert_recov_operation  // Alerts[0]
    };

  assign alert_recov_operation = shadowed_update_err;

  // The recoverable alert is observable via status register until the KMAC operation is restarted
  // by re-writing the Control Register.
  logic status_alert_recov_ctrl_update_err;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      status_alert_recov_ctrl_update_err <= 1'b 0;
    end else if (alert_recov_operation) begin
      status_alert_recov_ctrl_update_err <= 1'b 1;
    end else if (err_processed) begin
      status_alert_recov_ctrl_update_err <= 1'b 0;
    end
  end

  assign hw2reg.status.alert_recov_ctrl_update_err.d  = status_alert_recov_ctrl_update_err;

  assign alert_fatal = shadowed_storage_err
                     | alert_intg_err
                     | sparse_fsm_error
                     | counter_error
                     | control_integrity_error
                     ;

  // Make the fatal alert observable via status register.
  // Cannot be reset except the hardware reset
  logic status_alert_fatal_fault;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      status_alert_fatal_fault <= 1'b 0;
    end else if (alert_fatal) begin
      status_alert_fatal_fault <= 1'b 1;
    end
  end
  assign hw2reg.status.alert_fatal_fault.d  = status_alert_fatal_fault;

  for (genvar i = 0; i < NumAlerts; i++) begin : gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i)
    ) u_prim_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i] ),
      .alert_req_i   ( alerts[i]     ),
      .alert_ack_o   (               ),
      .alert_state_o (               ),
      .alert_rx_i    ( alert_rx_i[i] ),
      .alert_tx_o    ( alert_tx_o[i] )
    );
  end

  // Below assumes NumAlerts == 2
  `ASSERT_INIT(NumAlerts2_A, NumAlerts == 2)

  always_ff @(posedge clk_i or negedge rst_ni) begin
  // break up the combinatorial path for local escalation
    if (!rst_ni) begin
      alerts_q[1] <= 1'b0;
    end else if (alerts[1]) begin
      // fatal alerts cannot be cleared
      alerts_q[1] <= 1'b1;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
  // break up the combinatorial path for local escalation
    if (!rst_ni) begin
      alerts_q[0] <= 1'b0;
    end else begin
      // recoverable alerts can be cleared so just latch the value
      alerts_q[0] <= alerts[0];
    end
  end

  // Latched recoverable alert[0] is not used. Rather removing above,
  // keep alert_q[1:0] and make alert_q[0] unused (lint waive).
  logic unused_alerts_q0;
  assign unused_alerts_q0 = alerts_q[0];

  // SEC_CM: LC_ESCALATE_EN.INTERSIG.MUBI, FSM.GLOBAL_ESC, FSM.LOCAL_ESC
  lc_ctrl_pkg::lc_tx_t alert_to_lc_tx;
  assign alert_to_lc_tx = lc_ctrl_pkg::lc_tx_bool_to_lc_tx(alerts_q[1]);
  for (genvar i = 0; i < NumLcSyncCopies; i++) begin : gen_or_alert_lc_sync
      assign lc_escalate_en[i] = lc_ctrl_pkg::lc_tx_or_hi(alert_to_lc_tx, lc_escalate_en_sync[i]);
  end

  // Synchronize life cycle input
  prim_lc_sync #(
    .NumCopies (NumLcSyncCopies)
  ) u_prim_lc_sync (
    .clk_i,
    .rst_ni,
    .lc_en_i ( lc_escalate_en_i    ),
    .lc_en_o ( lc_escalate_en_sync )
  );

  assign en_masking_o = EnMasking;

  ////////////////
  // Assertions //
  ////////////////

  // Assert known for output values
  `ASSERT_KNOWN(KmacDone_A, intr_kmac_done_o)
  `ASSERT_KNOWN(FifoEmpty_A, intr_fifo_empty_o)
  `ASSERT_KNOWN(KmacErr_A, intr_kmac_err_o)
  `ASSERT_KNOWN(TlODValidKnown_A, tl_o.d_valid)
  `ASSERT_KNOWN(TlOAReadyKnown_A, tl_o.a_ready)
  `ASSERT_KNOWN(AlertKnownO_A, alert_tx_o)
  `ASSERT_KNOWN(EnMaskingKnown_A, en_masking_o)

  // Parameter as desired
  `ASSERT_INIT(SecretKeyDivideBy32_A, (kmac_pkg::MaxKeyLen % 32) == 0)

  // Command input should be sparse
  `ASSUME(CmdSparse_M, reg2hw.cmd.cmd.qe |-> reg2hw.cmd.cmd.q inside {CmdStart, CmdProcess,
                                                                CmdManualRun,CmdDone, CmdNone})

  // redundant counter error
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(SentMsgCountCheck_A, u_sha3.u_pad.u_sentmsg_count,
                                         alert_tx_o[1])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(RoundCountCheck_A, u_sha3.u_keccak.u_round_count,
                                         alert_tx_o[1])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(KeyIndexCountCheck_A, u_kmac_core.u_key_index_count,
                                         alert_tx_o[1])

  // Sparse FSM state error
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(KmacCoreFsmCheck_A, u_kmac_core.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(KmacAppFsmCheck_A, u_app_intf.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(SHA3FsmCheck_A, u_sha3.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(SHA3padFsmCheck_A, u_sha3.u_pad.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(KeccackFsmCheck_A, u_sha3.u_keccak.u_state_regs,
                                       alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(ErrorCheckFsmCheck_A, u_errchk.u_state_regs, alert_tx_o[1])
  `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(KmacFsmCheck_A, u_state_regs, alert_tx_o[1])

  // prim is only instantiated if masking is enabled
  if (EnMasking == 1) begin : g_testassertion
    `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(EntropyFsmCheck_A, gen_entropy.u_entropy.u_state_regs,
                                         alert_tx_o[1])

    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(HashCountCheck_A, gen_entropy.u_entropy.u_hash_count,
                                         alert_tx_o[1])
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(SeedIdxCountCheck_A,
                                           gen_entropy.u_entropy.u_seed_idx_count,
                                           alert_tx_o[1])

    // MsgFifo.Packer
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(
      PackerCountCheck_A,
      u_msgfifo.u_packer.g_pos_dupcnt.u_pos,
      alert_tx_o[1]
    )

    // MsgFifo.Fifo
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(
      MsgFifoWptrCheck_A,
      u_msgfifo.u_msgfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_wptr,
      alert_tx_o[1]
    )
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(
      MsgFifoRptrCheck_A,
      u_msgfifo.u_msgfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_rptr,
      alert_tx_o[1]
    )
  end

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A, u_reg, alert_tx_o[1])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module rom_ctrl_regs_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output rom_ctrl_reg_pkg::rom_ctrl_regs_reg2hw_t reg2hw, // Write
  input  rom_ctrl_reg_pkg::rom_ctrl_regs_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import rom_ctrl_reg_pkg::* ;

  localparam int AW = 7;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [17:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(18)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic alert_test_we;
  logic alert_test_wd;
  logic fatal_alert_cause_checker_error_qs;
  logic fatal_alert_cause_integrity_error_qs;
  logic [31:0] digest_0_qs;
  logic [31:0] digest_1_qs;
  logic [31:0] digest_2_qs;
  logic [31:0] digest_3_qs;
  logic [31:0] digest_4_qs;
  logic [31:0] digest_5_qs;
  logic [31:0] digest_6_qs;
  logic [31:0] digest_7_qs;
  logic [31:0] exp_digest_0_qs;
  logic [31:0] exp_digest_1_qs;
  logic [31:0] exp_digest_2_qs;
  logic [31:0] exp_digest_3_qs;
  logic [31:0] exp_digest_4_qs;
  logic [31:0] exp_digest_5_qs;
  logic [31:0] exp_digest_6_qs;
  logic [31:0] exp_digest_7_qs;

  // Register instances
  // R[alert_test]: V(True)
  logic alert_test_qe;
  logic [0:0] alert_test_flds_we;
  assign alert_test_qe = &alert_test_flds_we;
  prim_subreg_ext #(
    .DW    (1)
  ) u_alert_test (
    .re     (1'b0),
    .we     (alert_test_we),
    .wd     (alert_test_wd),
    .d      ('0),
    .qre    (),
    .qe     (alert_test_flds_we[0]),
    .q      (reg2hw.alert_test.q),
    .ds     (),
    .qs     ()
  );
  assign reg2hw.alert_test.qe = alert_test_qe;


  // R[fatal_alert_cause]: V(False)
  //   F[checker_error]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_checker_error (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.checker_error.de),
    .d      (hw2reg.fatal_alert_cause.checker_error.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_checker_error_qs)
  );

  //   F[integrity_error]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_fatal_alert_cause_integrity_error (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.fatal_alert_cause.integrity_error.de),
    .d      (hw2reg.fatal_alert_cause.integrity_error.d),

    // to internal hardware
    .qe     (),
    .q      (),
    .ds     (),

    // to register interface (read)
    .qs     (fatal_alert_cause_integrity_error_qs)
  );


  // Subregister 0 of Multireg digest
  // R[digest_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[0].de),
    .d      (hw2reg.digest[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_0_qs)
  );


  // Subregister 1 of Multireg digest
  // R[digest_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[1].de),
    .d      (hw2reg.digest[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_1_qs)
  );


  // Subregister 2 of Multireg digest
  // R[digest_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[2].de),
    .d      (hw2reg.digest[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_2_qs)
  );


  // Subregister 3 of Multireg digest
  // R[digest_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[3].de),
    .d      (hw2reg.digest[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_3_qs)
  );


  // Subregister 4 of Multireg digest
  // R[digest_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[4].de),
    .d      (hw2reg.digest[4].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_4_qs)
  );


  // Subregister 5 of Multireg digest
  // R[digest_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[5].de),
    .d      (hw2reg.digest[5].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_5_qs)
  );


  // Subregister 6 of Multireg digest
  // R[digest_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[6].de),
    .d      (hw2reg.digest[6].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_6_qs)
  );


  // Subregister 7 of Multireg digest
  // R[digest_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_digest_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.digest[7].de),
    .d      (hw2reg.digest[7].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.digest[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (digest_7_qs)
  );


  // Subregister 0 of Multireg exp_digest
  // R[exp_digest_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[0].de),
    .d      (hw2reg.exp_digest[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_0_qs)
  );


  // Subregister 1 of Multireg exp_digest
  // R[exp_digest_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[1].de),
    .d      (hw2reg.exp_digest[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_1_qs)
  );


  // Subregister 2 of Multireg exp_digest
  // R[exp_digest_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[2].de),
    .d      (hw2reg.exp_digest[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_2_qs)
  );


  // Subregister 3 of Multireg exp_digest
  // R[exp_digest_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[3].de),
    .d      (hw2reg.exp_digest[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_3_qs)
  );


  // Subregister 4 of Multireg exp_digest
  // R[exp_digest_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[4].de),
    .d      (hw2reg.exp_digest[4].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_4_qs)
  );


  // Subregister 5 of Multireg exp_digest
  // R[exp_digest_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[5].de),
    .d      (hw2reg.exp_digest[5].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_5_qs)
  );


  // Subregister 6 of Multireg exp_digest
  // R[exp_digest_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[6].de),
    .d      (hw2reg.exp_digest[6].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_6_qs)
  );


  // Subregister 7 of Multireg exp_digest
  // R[exp_digest_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_exp_digest_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.exp_digest[7].de),
    .d      (hw2reg.exp_digest[7].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.exp_digest[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (exp_digest_7_qs)
  );



  logic [17:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == ROM_CTRL_ALERT_TEST_OFFSET);
    addr_hit[ 1] = (reg_addr == ROM_CTRL_FATAL_ALERT_CAUSE_OFFSET);
    addr_hit[ 2] = (reg_addr == ROM_CTRL_DIGEST_0_OFFSET);
    addr_hit[ 3] = (reg_addr == ROM_CTRL_DIGEST_1_OFFSET);
    addr_hit[ 4] = (reg_addr == ROM_CTRL_DIGEST_2_OFFSET);
    addr_hit[ 5] = (reg_addr == ROM_CTRL_DIGEST_3_OFFSET);
    addr_hit[ 6] = (reg_addr == ROM_CTRL_DIGEST_4_OFFSET);
    addr_hit[ 7] = (reg_addr == ROM_CTRL_DIGEST_5_OFFSET);
    addr_hit[ 8] = (reg_addr == ROM_CTRL_DIGEST_6_OFFSET);
    addr_hit[ 9] = (reg_addr == ROM_CTRL_DIGEST_7_OFFSET);
    addr_hit[10] = (reg_addr == ROM_CTRL_EXP_DIGEST_0_OFFSET);
    addr_hit[11] = (reg_addr == ROM_CTRL_EXP_DIGEST_1_OFFSET);
    addr_hit[12] = (reg_addr == ROM_CTRL_EXP_DIGEST_2_OFFSET);
    addr_hit[13] = (reg_addr == ROM_CTRL_EXP_DIGEST_3_OFFSET);
    addr_hit[14] = (reg_addr == ROM_CTRL_EXP_DIGEST_4_OFFSET);
    addr_hit[15] = (reg_addr == ROM_CTRL_EXP_DIGEST_5_OFFSET);
    addr_hit[16] = (reg_addr == ROM_CTRL_EXP_DIGEST_6_OFFSET);
    addr_hit[17] = (reg_addr == ROM_CTRL_EXP_DIGEST_7_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(ROM_CTRL_REGS_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(ROM_CTRL_REGS_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(ROM_CTRL_REGS_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(ROM_CTRL_REGS_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(ROM_CTRL_REGS_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(ROM_CTRL_REGS_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(ROM_CTRL_REGS_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(ROM_CTRL_REGS_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(ROM_CTRL_REGS_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(ROM_CTRL_REGS_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(ROM_CTRL_REGS_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(ROM_CTRL_REGS_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(ROM_CTRL_REGS_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(ROM_CTRL_REGS_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(ROM_CTRL_REGS_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(ROM_CTRL_REGS_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(ROM_CTRL_REGS_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(ROM_CTRL_REGS_PERMIT[17] & ~reg_be)))));
  end

  // Generate write-enables
  assign alert_test_we = addr_hit[0] & reg_we & !reg_error;

  assign alert_test_wd = reg_wdata[0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = alert_test_we;
    reg_we_check[1] = 1'b0;
    reg_we_check[2] = 1'b0;
    reg_we_check[3] = 1'b0;
    reg_we_check[4] = 1'b0;
    reg_we_check[5] = 1'b0;
    reg_we_check[6] = 1'b0;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = 1'b0;
    reg_we_check[9] = 1'b0;
    reg_we_check[10] = 1'b0;
    reg_we_check[11] = 1'b0;
    reg_we_check[12] = 1'b0;
    reg_we_check[13] = 1'b0;
    reg_we_check[14] = 1'b0;
    reg_we_check[15] = 1'b0;
    reg_we_check[16] = 1'b0;
    reg_we_check[17] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = '0;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = fatal_alert_cause_checker_error_qs;
        reg_rdata_next[1] = fatal_alert_cause_integrity_error_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = digest_0_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = digest_1_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = digest_2_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = digest_3_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = digest_4_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = digest_5_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = digest_6_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = digest_7_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = exp_digest_0_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = exp_digest_1_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = exp_digest_2_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = exp_digest_3_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = exp_digest_4_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = exp_digest_5_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = exp_digest_6_qs;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = exp_digest_7_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module rom_ctrl_rom_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t64 tl_i,
  output tlul_pkg::tl_d2h_t64 tl_o,

  // Output port for window
  output tlul_pkg::tl_h2d_t64 tl_win_o,
  input  tlul_pkg::tl_d2h_t64 tl_win_i,

  // To HW

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import rom_ctrl_reg_pkg::* ;


  // Add an unloaded flop to make use of clock / reset
  // This is done to specifically address lint complaints of unused clocks/resets
  // Since the flop is unloaded it will be removed during synthesis
  logic unused_reg;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      unused_reg <= '0;
    end else begin
      unused_reg <= tl_i.a_valid;
    end
  end



  // Since there are no registers in this block, commands are routed through to windows which
  // can report their own integrity errors.
  assign intg_err_o = 1'b0;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t64 tl_o_pre;

  //zdr: del tlul_rsp_intg_gen
  // tlul_rsp_intg_gen #(
  //   .EnableRspIntgGen(0),
  //   .EnableDataIntgGen(0)
  // ) u_rsp_intg_gen (
  //   .tl_i(tl_o_pre),
  //   .tl_o(tl_o)
  // );
  assign tl_o = tl_o_pre;

  assign tl_win_o = tl_i;
  assign tl_o_pre = tl_win_i;

  // Unused signal tieoff
  // devmode_i is not used if there are no registers
  logic unused_devmode;
  assign unused_devmode = ^devmode_i;
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

module rom_ctrl
  import rom_ctrl_reg_pkg::NumAlerts;
  import prim_rom_pkg::rom_cfg_t;
#(
  parameter                       BootRomInitFile = "",
  parameter logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b1}},
  parameter bit [63:0]            RndCnstScrNonce = '0,
  parameter bit [127:0]           RndCnstScrKey = '0,

  // Disable all (de)scrambling operation. This disables both the scrambling block and the boot-time
  // checker. Don't use this in a real chip, but it's handy for small FPGA targets where we don't
  // want to spend area on unused scrambling.
  parameter bit                   SecDisableScrambling = 1'b0
) (
  input  clk_i,
  input  rst_ni,

  // ROM configuration parameters
  input  rom_cfg_t rom_cfg_i,

  input  tlul_pkg::tl_h2d_t64 rom_tl_i,
  output tlul_pkg::tl_d2h_t64 rom_tl_o,

  input  tlul_pkg::tl_h2d_t regs_tl_i,
  output tlul_pkg::tl_d2h_t regs_tl_o,

  // Alerts
  input  prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i,
  output prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o,

  // Connections to other blocks
  output rom_ctrl_pkg::pwrmgr_data_t pwrmgr_data_o,
  output rom_ctrl_pkg::keymgr_data_t keymgr_data_o,
  input  kmac_pkg::app_rsp_t         kmac_data_i,
  output kmac_pkg::app_req_t         kmac_data_o
);

  import rom_ctrl_pkg::*;
  import rom_ctrl_reg_pkg::*;
  import prim_mubi_pkg::mubi4_t, prim_mubi_pkg::MuBi4True;
  import prim_util_pkg::vbits;

  `define CLK_WAIT_BOUNDS ##[MIN_CLK_WAIT_CYCLES:MAX_CLK_WAIT_CYCLES]
  // ROM_CTRL_ROM_SIZE is auto-generated by regtool and comes from the bus window size, measured in
  // bytes of content (i.e. 4 times the number of 32 bit words).
  localparam int unsigned RomSizeByte = ROM_CTRL_ROM_SIZE;
  localparam int unsigned RomSizeWords = RomSizeByte >> 2;
  localparam int unsigned RomIndexWidth = vbits(RomSizeWords);

  // DataWidth is normally 39, representing 32 bits of actual data plus 7 ECC check bits. If
  // scrambling is disabled ("insecure mode"), we store a raw 32-bit image and generate ECC check
  // bits on the fly.
  localparam int unsigned DataWidth = SecDisableScrambling ? 32 : 64;

  mubi4_t                   rom_select_bus;

  logic [RomIndexWidth-1:0] rom_rom_index, rom_prince_index;
  logic                     rom_req;
  logic [DataWidth-1:0]     rom_scr_rdata;
  logic [DataWidth-1:0]     rom_clr_rdata;
  logic                     rom_rvalid;

  logic [RomIndexWidth-1:0] bus_rom_rom_index, bus_rom_prince_index;
  logic                     bus_rom_req;
  logic                     bus_rom_gnt;
  logic [DataWidth-1:0]     bus_rom_rdata;
  logic                     bus_rom_rvalid, bus_rom_rvalid_raw;

  logic [RomIndexWidth-1:0] checker_rom_index;
  logic                     checker_rom_req;
  logic [DataWidth-1:0]     checker_rom_rdata;

  logic                     internal_alert;

  // Pack / unpack kmac connection data ========================================

  logic [63:0]              kmac_rom_data;
  logic                     kmac_rom_rdy;
  logic                     kmac_rom_vld;
  logic                     kmac_rom_last;
  logic                     kmac_done;
  logic [255:0]             kmac_digest;
  logic                     kmac_err;

  if (!SecDisableScrambling) begin : gen_kmac_scramble_enabled
    // The usual situation, with scrambling enabled. Collect up output signals for kmac and split up
    // the input struct into separate signals.

    // Neglecting any first / last block effects, and assuming that ROM_CTRL can always fill the
    // KMAC message FIFO while a KMAC round is running, the total processing time for a 32kB ROM is
    // calculated as follows:
    //
    // (Padding Overhead) x (ROM Size) / (Block Size) x (Block Processing Time + KMAC Absorb Time)
    //
    // ROM_CTRL can only read out one 32 or 39 bit (with ECC) word per cycle, so if we were to zero
    // pad this to align with the 64bit KMAC interface, the padding overhead would amount to 2x
    // in this equation:
    //
    // 2 x 32 kByte / (1600 bit - 2x 256bit) x (96 cycles + (1600 bit - 2x 256bit) / 64bit)) =
    // 2 x 32 x 1024 x 8bit / 1088bit x (96 cycles + 17 cycles) =
    // 2 x 262144 bit / 1088 bit x 113 cycles =
    // 2 x 27226.35 cycles
    //
    // Luckily, the KMAC interface allows to transmit data with a byte enable mask, and only the
    // enabled bytes will be packed into the message FIFO. Assuming that the processing is the
    // bottleneck, we can thus reduce the overhead of 2x in that equation to 1x or 5/8x if we only
    // set 4 or 5 byte enables (4 for 32bit, 5 for 39bit)!
    localparam int NumBytes = (DataWidth + 7) / 8;

    // SEC_CM: MEM.DIGEST
    assign kmac_data_o = '{valid: kmac_rom_vld,
                           data: kmac_rom_data,
                           strb: kmac_pkg::MsgStrbW'({NumBytes{1'b1}}),
                           last: kmac_rom_last};

    assign kmac_rom_rdy = kmac_data_i.ready;
    assign kmac_done = kmac_data_i.done;
    assign kmac_digest = kmac_data_i.digest_share0[255:0] ^ kmac_data_i.digest_share1[255:0];
    assign kmac_err = kmac_data_i.error;

    logic unused_kmac_digest;
    assign unused_kmac_digest = ^{
      kmac_data_i.digest_share0[kmac_pkg::AppDigestW-1:256],
      kmac_data_i.digest_share1[kmac_pkg::AppDigestW-1:256]
    };

  end : gen_kmac_scramble_enabled
  else begin : gen_kmac_scramble_disabled
    // Scrambling is disabled. Stub out all KMAC connections and waive the ignored signals.

    assign kmac_data_o = '0;
    assign kmac_rom_rdy = 1'b0;
    assign kmac_done = 1'b0;
    assign kmac_digest = '0;
    assign kmac_err = 1'b0;

    logic unused_kmac_inputs;
    assign unused_kmac_inputs = ^{kmac_data_i};

    logic unused_kmac_outputs;
    assign unused_kmac_outputs = ^{kmac_rom_vld, kmac_rom_data, kmac_rom_last};

  end : gen_kmac_scramble_disabled

  // TL interface ==============================================================

  tlul_pkg::tl_h2d_t64 tl_rom_h2d_upstream, tl_rom_h2d_downstream;
  tlul_pkg::tl_d2h_t64 tl_rom_d2h;

  logic  rom_reg_integrity_error;

  rom_ctrl_rom_reg_top u_rom_top (
    .clk_i,
    .rst_ni,
    .tl_i       (rom_tl_i),
    .tl_o       (rom_tl_o),
    .tl_win_o   (tl_rom_h2d_upstream),
    .tl_win_i   (tl_rom_d2h),

    .intg_err_o (rom_reg_integrity_error),    // SEC_CM: BUS.INTEGRITY

    .devmode_i  (1'b1)
  );

  // This buffer ensures that when we calculate bus_rom_prince_index by snooping on
  // tl_rom_h2d_upstream, we get a value that's buffered from the thing that goes into both the ECC
  // check and the addr_o output of u_tl_adapter_rom. That way, an injected 1- or 2-bit fault that
  // affects bus_rom_prince_index must either affect the ECC check (causing it to fail) OR it cannot
  // affect bus_rom_rom_index (so the address-tweakable scrambling will mean the read probably gets
  // garbage).
  //
  // SEC_CM: CTRL.REDUN
  prim_buf #(
    .Width($bits(tlul_pkg::tl_h2d_t64))
  ) u_tl_rom_h2d_buf (
    .in_i (tl_rom_h2d_upstream),
    .out_o (tl_rom_h2d_downstream)
  );

  // Bus -> ROM adapter ========================================================

  logic rom_integrity_error;

  tlul_adapter_sram64 #(
    .SramAw(RomIndexWidth),
    .SramDw(64),
    .Outstanding(2),
    .ByteAccess(0),
    .ErrOnWrite(1),
    .CmdIntgCheck(0),
    .EnableRspIntgGen(0),
    .EnableDataIntgGen(SecDisableScrambling),
    .EnableDataIntgPt(SecDisableScrambling), // SEC_CM: BUS.INTEGRITY
    .SecFifoPtr      (1)                      // SEC_CM: TLUL_FIFO.CTR.REDUN
  ) u_tl_adapter_rom (
    .clk_i,
    .rst_ni,

    .tl_i         (tl_rom_h2d_downstream),
    .tl_o         (tl_rom_d2h),
    .en_ifetch_i  (prim_mubi_pkg::MuBi4True),
    .req_o        (bus_rom_req),
    .req_type_o   (),
    .gnt_i        (bus_rom_gnt),
    .we_o         (),
    .addr_o       (bus_rom_rom_index),
    .wdata_o      (),
    .wmask_o      (),
    .intg_error_o (rom_integrity_error),
    .rdata_i      (bus_rom_rdata),
    .rvalid_i     (bus_rom_rvalid),
    .rerror_i     (2'b00)
  );

  // Snoop on the "upstream" TL transaction to infer the address to pass to the PRINCE cipher.
  // zdr: addr 2-> 3 for 64bit
  assign bus_rom_prince_index = (tl_rom_h2d_upstream.a_valid ?
                                 tl_rom_h2d_upstream.a_address[3 +: RomIndexWidth] :
                                 '0);

  // Unless there has been an injected fault, bus_rom_prince_index and bus_rom_rom_index should have
  // the same value.
  `ASSERT(BusRomIndicesMatch_A, bus_rom_prince_index == bus_rom_rom_index)

  // The mux ===================================================================

  logic mux_alert;

  rom_ctrl_mux #(
    .AW (RomIndexWidth),
    .DW (DataWidth)
  ) u_mux (
    .clk_i,
    .rst_ni,
    .sel_bus_i         (rom_select_bus),
    .bus_rom_addr_i    (bus_rom_rom_index),
    .bus_prince_addr_i (bus_rom_prince_index),
    .bus_req_i         (bus_rom_req),
    .bus_gnt_o         (bus_rom_gnt),
    .bus_rdata_o       (bus_rom_rdata),
    .bus_rvalid_o      (bus_rom_rvalid_raw),
    .chk_addr_i        (checker_rom_index),
    .chk_req_i         (checker_rom_req),
    .chk_rdata_o       (checker_rom_rdata),
    .rom_rom_addr_o    (rom_rom_index),
    .rom_prince_addr_o (rom_prince_index),
    .rom_req_o         (rom_req),
    .rom_scr_rdata_i   (rom_scr_rdata),
    .rom_clr_rdata_i   (rom_clr_rdata),
    .rom_rvalid_i      (rom_rvalid),
    .alert_o           (mux_alert)
  );

  // Squash all responses from the ROM to the bus if there's an internal integrity error from the
  // checker FSM or the mux. This avoids having to handle awkward corner cases in the mux: if
  // something looks bad, we'll complain and hang the bus transaction.
  //
  // Note that the two signals that go into internal_alert are both sticky. The mux explicitly
  // latches its alert_o output and the checker FSM jumps to an invalid scrap state when it sees an
  // error which, in turn, sets checker_alert.
  //
  // SEC_CM: BUS.LOCAL_ESC
  assign bus_rom_rvalid = bus_rom_rvalid_raw & !internal_alert;

  // The ROM itself ============================================================

  if (!SecDisableScrambling) begin : gen_rom_scramble_enabled

    // SEC_CM: MEM.SCRAMBLE
    rom_ctrl_scrambled_rom #(
      .MemInitFile (BootRomInitFile),
      .Width       (DataWidth),
      .Depth       (RomSizeWords),
      .ScrNonce    (RndCnstScrNonce),
      .ScrKey      (RndCnstScrKey)
    ) u_rom (
      .clk_i,
      .rst_ni,
      .req_i         (rom_req),
      .rom_addr_i    (rom_rom_index),
      .prince_addr_i (rom_prince_index),
      .rvalid_o      (rom_rvalid),
      .scr_rdata_o   (rom_scr_rdata),
      .clr_rdata_o   (rom_clr_rdata),
      .cfg_i         (rom_cfg_i)
    );

  end : gen_rom_scramble_enabled
  else begin : gen_rom_scramble_disabled

    // If scrambling is disabled then instantiate a normal ROM primitive (no PRINCE cipher etc.).
    // Note that this "raw memory" doesn't have ECC bits either.

    prim_rom_adv #(
      .Width       (DataWidth),
      .Depth       (RomSizeWords),
      .MemInitFile (BootRomInitFile)
    ) u_rom (
      .clk_i,
      .rst_ni,
      .req_i    (rom_req),
      .addr_i   (rom_rom_index),
      .rvalid_o (rom_rvalid),
      .rdata_o  (rom_scr_rdata),
      .cfg_i    (rom_cfg_i)
    );

    // There's no scrambling, so "scrambled" and "clear" rdata are equal.
    assign rom_clr_rdata = rom_scr_rdata;

    // Since we're not generating a keystream, we don't use the rom_prince_index at all
    logic unused_prince_index;
    assign unused_prince_index = ^rom_prince_index;

  end : gen_rom_scramble_disabled

  // Zero expand checker rdata to pass to KMAC
  assign kmac_rom_data = {{64-DataWidth{1'b0}}, checker_rom_rdata};

  // Register block ============================================================

  rom_ctrl_regs_reg2hw_t reg2hw;
  rom_ctrl_regs_hw2reg_t hw2reg;
  logic                  reg_integrity_error;

  rom_ctrl_regs_reg_top u_reg_regs (
    .clk_i,
    .rst_ni,
    .tl_i       (regs_tl_i),
    .tl_o       (regs_tl_o),
    .reg2hw     (reg2hw),
    .hw2reg     (hw2reg),
    .intg_err_o (reg_integrity_error),    // SEC_CM: BUS.INTEGRITY
    .devmode_i  (1'b1)
   );

  // The checker FSM ===========================================================

  logic [255:0] digest_q, exp_digest_q;
  logic [255:0] digest_d;
  logic         digest_de;
  logic [63:0]  exp_digest_word_d;
  logic         exp_digest_de;
  logic [1:0]   exp_digest_idx;

  logic         checker_alert;

  if (!SecDisableScrambling) begin : gen_fsm_scramble_enabled

    rom_ctrl_fsm #(
      .RomDepth (RomSizeWords),
      .TopCount (4)
    ) u_checker_fsm (
      .clk_i,
      .rst_ni,
      .digest_i             (digest_q),
      .exp_digest_i         (exp_digest_q),
      .digest_o             (digest_d),
      .digest_vld_o         (digest_de),
      .exp_digest_o         (exp_digest_word_d),
      .exp_digest_vld_o     (exp_digest_de),
      .exp_digest_idx_o     (exp_digest_idx),
      .pwrmgr_data_o        (pwrmgr_data_o),
      .keymgr_data_o        (keymgr_data_o),
      .kmac_rom_rdy_i       (kmac_rom_rdy),
      .kmac_rom_vld_o       (kmac_rom_vld),
      .kmac_rom_last_o      (kmac_rom_last),
      .kmac_done_i          (kmac_done),
      .kmac_digest_i        (kmac_digest),
      .kmac_err_i           (kmac_err),
      .rom_select_bus_o     (rom_select_bus),
      .rom_addr_o           (checker_rom_index),
      .rom_req_o            (checker_rom_req),
      .rom_data_i           (checker_rom_rdata[63:0]),
      .alert_o              (checker_alert)
    );

  end : gen_fsm_scramble_enabled
  else begin : gen_fsm_scramble_disabled

    // If scrambling is disabled, there's no checker FSM.

    assign digest_d = '0;
    assign digest_de = 1'b0;
    assign exp_digest_word_d = '0;
    assign exp_digest_de = 1'b0;
    assign exp_digest_idx = '0;

    assign pwrmgr_data_o = PWRMGR_DATA_DEFAULT;
    // Send something other than '1 or '0 because the key manager has an "all ones" and an "all
    // zeros" check.
    assign keymgr_data_o = '{data: {128{2'b10}}, valid: 1'b1};

    assign kmac_rom_vld = 1'b0;
    assign kmac_rom_last = 1'b0;

    // Always grant access to the bus. Setting this to a constant should mean the mux gets
    // synthesized away completely.
    assign rom_select_bus = MuBi4True;

    assign checker_rom_index = '0;
    assign checker_rom_req = 1'b0;
    assign checker_alert = 1'b0;

    logic unused_fsm_inputs;
    assign unused_fsm_inputs = ^{kmac_rom_rdy, kmac_done, kmac_digest, digest_q, exp_digest_q};

  end : gen_fsm_scramble_disabled

  // // Register data =============================================================

  // // DIGEST and EXP_DIGEST registers

  // // Repack signals to convert between the view expected by rom_ctrl_reg_pkg for CSRs and the view
  // // expected by rom_ctrl_fsm. Register 0 of a multi-reg appears as the low bits of the packed data.
  // for (genvar i = 0; i < 8; i++) begin: gen_csr_digest
  //   localparam int unsigned TopBitInt = 32 * i + 31;
  //   localparam bit [7:0] TopBit = TopBitInt[7:0];

  //   assign hw2reg.digest[i].d = digest_d[TopBit -: 32];
  //   assign hw2reg.digest[i].de = digest_de;

  //   assign hw2reg.exp_digest[i].d = exp_digest_word_d;
  //   assign hw2reg.exp_digest[i].de = exp_digest_de && (i[2:0] == exp_digest_idx);

  //   assign digest_q[TopBit -: 32] = reg2hw.digest[i].q;
  //   assign exp_digest_q[TopBit -: 32] = reg2hw.exp_digest[i].q;
  // end

  // Register data =============================================================

  // DIGEST and EXP_DIGEST registers

  // Repack signals to convert between the view expected by rom_ctrl_reg_pkg for CSRs and the view
  // expected by rom_ctrl_fsm. Register 0 of a multi-reg appears as the low bits of the packed data.
  for (genvar i = 0; i < 4; i++) begin: gen_csr_digest
    localparam int unsigned TopBitInt = 64 * i + 63;  // Change from 32 to 64
    localparam bit [7:0] TopBit = TopBitInt[7:0];

    assign hw2reg.digest[2*i].d = digest_d[TopBit -: 32];  // Low 32 bits
    assign hw2reg.digest[2*i].de = digest_de;

    assign hw2reg.digest[2*i+1].d = digest_d[TopBit - 32 -: 32];  // High 32 bits
    assign hw2reg.digest[2*i+1].de = digest_de;

    assign hw2reg.exp_digest[2*i].d = exp_digest_word_d[63:32];
    assign hw2reg.exp_digest[2*i].de = exp_digest_de && (i[1:0] == exp_digest_idx);

    assign hw2reg.exp_digest[2*i+1].d = exp_digest_word_d[31:0];
    assign hw2reg.exp_digest[2*i+1].de = exp_digest_de && (i[1:0] == exp_digest_idx);

    assign digest_q[TopBit -: 32] = reg2hw.digest[2*i].q;
    assign digest_q[TopBit - 32 -: 32] = reg2hw.digest[2*i+1].q;

    assign exp_digest_q[TopBit -: 32] = reg2hw.exp_digest[2*i].q;
    assign exp_digest_q[TopBit - 32 -: 32] = reg2hw.exp_digest[2*i+1].q;
  end

  logic bus_integrity_error;
  assign bus_integrity_error = rom_reg_integrity_error | rom_integrity_error | reg_integrity_error;

  assign internal_alert = checker_alert | mux_alert;

  // FATAL_ALERT_CAUSE register
  assign hw2reg.fatal_alert_cause.checker_error.d  = internal_alert;
  assign hw2reg.fatal_alert_cause.checker_error.de = internal_alert;
  assign hw2reg.fatal_alert_cause.integrity_error.d  = bus_integrity_error;
  assign hw2reg.fatal_alert_cause.integrity_error.de = bus_integrity_error;

  // Alert generation ==========================================================

  logic [NumAlerts-1:0] alert_test;
  assign alert_test[AlertFatal] = reg2hw.alert_test.q &
                                  reg2hw.alert_test.qe;

  logic [NumAlerts-1:0] alerts;
  assign alerts[AlertFatal] = bus_integrity_error | checker_alert | mux_alert;

  for (genvar i = 0; i < NumAlerts; i++) begin: gen_alert_tx
    prim_alert_sender #(
      .AsyncOn(AlertAsyncOn[i]),
      .IsFatal(i == AlertFatal)
    ) u_alert_sender (
      .clk_i,
      .rst_ni,
      .alert_test_i  ( alert_test[i] ),
      .alert_req_i   ( alerts[i]     ),
      .alert_ack_o   (               ),
      .alert_state_o (               ),
      .alert_rx_i    ( alert_rx_i[i] ),
      .alert_tx_o    ( alert_tx_o[i] )
    );
  end

  // Asserts ===================================================================
  //
  // "ROM" TL interface: The d_valid and a_ready signals should be unconditionally defined. The
  // other signals in rom_tl_o (which are the other D channel signals) should be defined if d_valid.
  `ASSERT_KNOWN(RomTlODValidKnown_A, rom_tl_o.d_valid)
  `ASSERT_KNOWN(RomTlOAReadyKnown_A, rom_tl_o.a_ready)
  `ASSERT_KNOWN_IF(RomTlODDataKnown_A, rom_tl_o, rom_tl_o.d_valid)

  // "regs" TL interface: The d_valid and a_ready signals should be unconditionally defined. The
  // other signals in rom_tl_o (which are the other D channel signals) should be defined if d_valid.
  `ASSERT_KNOWN(RegsTlODValidKnown_A, regs_tl_o.d_valid)
  `ASSERT_KNOWN(RegsTlOAReadyKnown_A, regs_tl_o.a_ready)
  `ASSERT_KNOWN_IF(RegsTlODDataKnown_A, regs_tl_o, regs_tl_o.d_valid)

  // The assert_tx_o output should have a known value when out of reset
  `ASSERT_KNOWN(AlertTxOKnown_A, alert_tx_o)

  // Assertions to check that we've wired up our alert bits correctly
  if (!SecDisableScrambling) begin : gen_asserts_with_scrambling
    `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CompareFsmAlert_A,
                                         gen_fsm_scramble_enabled.
                                         u_checker_fsm.u_compare.u_state_regs,
                                         alert_tx_o[AlertFatal])
    `ASSERT_PRIM_FSM_ERROR_TRIGGER_ALERT(CheckerFsmAlert_A,
                                         gen_fsm_scramble_enabled.
                                         u_checker_fsm.u_state_regs,
                                         alert_tx_o[AlertFatal])
    `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(CompareAddrCtrCheck_A,
                                           gen_fsm_scramble_enabled.
                                           u_checker_fsm.u_compare.u_prim_count_addr,
                                           alert_tx_o[AlertFatal])
  end

  // The pwrmgr_data_o output (the "done" and "good" signals) should have a known value when out of
  // reset. (In theory, the "good" signal could be unknown when !done, but the stronger and simpler
  // assertion is also true, so we use that)
  `ASSERT_KNOWN(PwrmgrDataOKnown_A, pwrmgr_data_o)

  // The valid signal for keymgr_data_o should always be known when out of reset. The rest of the
  // struct (a data signal) should be known whenever the valid signal is true.
  `ASSERT_KNOWN(KeymgrDataOValidKnown_A, keymgr_data_o.valid)
  `ASSERT_KNOWN_IF(KeymgrDataODataKnown_A, keymgr_data_o, keymgr_data_o.valid)

  // The valid signal for kmac_data_o should always be known when out of reset. The rest of the
  // struct (data, strb and last) should be known whenever the valid signal is true.
  `ASSERT_KNOWN(KmacDataOValidKnown_A, kmac_data_o.valid)
  `ASSERT_KNOWN_IF(KmacDataODataKnown_A, kmac_data_o, kmac_data_o.valid)

  // Check that pwrmgr_data_o.good is stable when kmac_data_o.valid is asserted
  `ASSERT(StabilityChkKmac_A, kmac_data_o.valid && $past(kmac_data_o.valid)
          |-> $stable(pwrmgr_data_o.good))

  // Check that pwrmgr_data_o.good is stable when keymgr_data_o.valid is asserted
  `ASSERT(StabilityChkkeymgr_A, keymgr_data_o.valid && $past(keymgr_data_o.valid)
          |-> $stable(pwrmgr_data_o.good))

  // Check that pwrmgr_data_o.done is never de-asserted once asserted
  `ASSERT(PwrmgrDataChk_A, $rose(pwrmgr_data_o.done == prim_mubi_pkg::MuBi4True) |->
          always !$fell(pwrmgr_data_o.done == prim_mubi_pkg::MuBi4True),
          clk_i, !rst_ni || internal_alert)

  // Check that keymgr_data_o.valid is never de-asserted once asserted
  `ASSERT(KeymgrValidChk_A, $rose(keymgr_data_o.valid) |-> always !$fell(keymgr_data_o.valid),
          clk_i, !rst_ni || internal_alert)

  // Check that rom_tl_o.d_valid is not asserted unless pwrmgr_data_o.done is asseterd.
  // This check ensures that all tl accesses are blocked until rom check is completed. You might
  // think we could check for a_ready, but that doesn't work because the TL to SRAM adapter has a
  // 1-entry cache that accepts the transaction (but doesn't reply)
  `ASSERT(TlAccessChk_A,
          (pwrmgr_data_o.done == prim_mubi_pkg::MuBi4False) |->
          (!rom_tl_o.d_valid || (rom_tl_o.d_valid && rom_tl_o.d_error)))

  // Check that whenever there is an alert triggered and FSM state is Invalid, there is no response
  // to read requests.
  if (!SecDisableScrambling) begin : gen_fsm_scramble_enabled_asserts

    `ASSERT(BusLocalEscChk_A,
            (gen_fsm_scramble_enabled.u_checker_fsm.state_d == rom_ctrl_pkg::Invalid)
            |-> always(!bus_rom_rvalid))
  end

  // Alert assertions for reg_we onehot check
  `ASSERT_PRIM_REG_WE_ONEHOT_ERROR_TRIGGER_ALERT(RegWeOnehotCheck_A,
                                                 u_reg_regs, alert_tx_o[AlertFatal])

  // Alert assertions for redundant counters.
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(FifoWptrCheck_A,
      u_tl_adapter_rom.u_rspfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_wptr,
      alert_tx_o[AlertFatal])
  `ASSERT_PRIM_COUNT_ERROR_TRIGGER_ALERT(FifoRptrCheck_A,
      u_tl_adapter_rom.u_rspfifo.gen_normal_fifo.u_fifo_cnt.gen_secure_ptrs.u_rptr,
      alert_tx_o[AlertFatal])
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

//
// The comparator inside the ROM checker
//
// This module is in charge of comparing the digest that was computed over the ROM data with the
// expected digest stored in the top few words.
//

`include "prim_assert.sv"

module rom_ctrl_compare
  import prim_mubi_pkg::mubi4_t;
#(
  parameter int NumWords = 2
) (
  input logic                        clk_i,
  input logic                        rst_ni,

  input logic                        start_i,
  output logic                       done_o,
  output mubi4_t                     good_o,

  // CSR inputs for DIGEST and EXP_DIGEST. Ordered with word 0 as LSB.
  input logic [NumWords*64-1:0]      digest_i,
  input logic [NumWords*64-1:0]      exp_digest_i,

  // To alert system
  output logic                       alert_o
);

  import prim_util_pkg::vbits;
  import prim_mubi_pkg::mubi4_bool_to_mubi;

  `ASSERT_INIT(NumWordsPositive_A, 0 < NumWords)

  localparam int AW = vbits(NumWords);

  localparam int unsigned LastAddrInt = NumWords - 1;
  localparam bit [AW-1:0] LastAddr    = LastAddrInt[AW-1:0];

  logic          addr_incr;
  logic [AW-1:0] addr_q;

  // This module must wait until triggered by a write to start_i. At that point, it cycles through
  // the words of DIGEST and EXP_DIGEST, comparing them to one another and passing each digest word
  // to the key manager. Finally, it gets to the Done state.
  //
  // States:
  //
  //    Waiting
  //    Checking
  //    Done
  //
  // Encoding generated with:
  // $ util/design/sparse-fsm-encode.py -d 3 -m 3 -n 5 -s 1 --language=sv
  //
  // Hamming distance histogram:
  //
  //  0: --
  //  1: --
  //  2: --
  //  3: |||||||||||||||||||| (66.67%)
  //  4: |||||||||| (33.33%)
  //  5: --
  //
  // Minimum Hamming distance: 3
  // Maximum Hamming distance: 4
  // Minimum Hamming weight: 1
  // Maximum Hamming weight: 3
  //
  // SEC_CM: FSM.SPARSE
  typedef enum logic [4:0] {
    Waiting  = 5'b00100,
    Checking = 5'b10010,
    Done     = 5'b11001
  } state_e;

  state_e state_q, state_d;
  logic   matches_q, matches_d;
  logic   fsm_alert;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, state_e, Waiting)

  always_comb begin
    state_d = state_q;
    fsm_alert = 1'b0;
    unique case (state_q)
      Waiting: begin
        if (start_i) state_d = Checking;
      end
      Checking: begin
        if (addr_q == LastAddr) state_d = Done;
      end
      Done: begin
        // Final state
      end
      default: fsm_alert = 1'b1;
    endcase
  end

  // start_i should only be signalled when we're in the Waiting state
  //
  // SEC_CM: COMPARE.CTRL_FLOW.CONSISTENCY
  logic start_alert;
  assign start_alert = start_i && (state_q != Waiting);

  // addr_q should be zero when we're in the Waiting state
  //
  // SEC_CM: COMPARE.CTR.CONSISTENCY
  logic wait_addr_alert;
  assign wait_addr_alert = (state_q == Waiting) && (addr_q != '0);

  // addr_q should be LastAddr when we're in the Done state
  //
  // SEC_CM: COMPARE.CTR.CONSISTENCY
  logic done_addr_alert;
  assign done_addr_alert = (state_q == Done) && (addr_q != LastAddr);

  // Increment addr_q on each cycle except the last when in Checking. The prim_count primitive
  // doesn't overflow but in case NumWords is not a power of 2, we need to take care of this
  // ourselves.
  assign addr_incr = (state_q == Checking) && (addr_q != LastAddr);

  // SEC_CM: COMPARE.CTR.REDUN
  logic addr_ctr_alert;
  prim_count #(
    .Width(AW)
  ) u_prim_count_addr (
    .clk_i,
    .rst_ni,
    .clr_i(1'b0),
    .set_i(1'b0),
    .set_cnt_i('0),
    .incr_en_i(addr_incr),
    .decr_en_i(1'b0),
    .step_i(AW'(1)),
    .cnt_o(addr_q),
    .cnt_next_o(),
    .err_o(addr_ctr_alert)
  );

  logic [AW+5-1:0] digest_idx;
  logic [31:0]     digest_word, exp_digest_word;
  assign digest_idx = {addr_q, 5'd31};
  assign digest_word = digest_i[digest_idx -: 32];
  assign exp_digest_word = exp_digest_i[digest_idx -: 32];

  assign matches_d = matches_q && (digest_word == exp_digest_word);
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      matches_q <= 1'b1;
    end else begin
      if (state_q == Checking) begin
        matches_q <= matches_d;
      end
    end
  end

  assign done_o = (state_q == Done);

  // Instantiate an explicit prim_mubi4_sender for the good signal. The logic is that we don't want
  // to make the actual check multi-bit (doing so properly would mean replicating the 32-bit
  // comparator) but we *do* want to make sure a synthesis tool doesn't optimize away the 4-bit
  // signal. The barrier from the primitive ensures that won't happen.
  prim_mubi4_sender
  u_done_sender (
    .clk_i,
    .rst_ni,
    .mubi_i (mubi4_bool_to_mubi(matches_q)),
    .mubi_o (good_o)
  );

  assign alert_o = fsm_alert | start_alert | wait_addr_alert | done_addr_alert | addr_ctr_alert;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

//
// A counter module that drives the ROM accesses from the checker.
//
// This module doesn't need state hardening: an attacker that glitches its behaviour can stall the
// chip or read ROM data in the wrong order. Assuming we've picked a key for the ROM that ensures
// all words have different values, exploiting a glitch in this module to hide a ROM modification
// would still need a pre-image attack on SHA-3.
//
// RomDepth is the number of words in the ROM. RomTopCount is the number of those words (at the top
// of the address space) that are considered part of the expected hash.
//
// When it comes out of reset, the module starts reading from address zero. Once the reading is
// done, it will signal done_o. The surrounding (hardened) design should check that done_o never has
// a high -> low transition.
//
// The read_addr_o signal should be connected to the stateful mux that controls access to ROM. This
// mux gives access to the rom_ctrl_counter until done_o is asserted. The data_addr_o signal gives
// the address of the ROM word that was just read.
//
// The data_* signals are used to handshake with KMAC, although the surrounding FSM will step in
// once we've got to the top of memory. The counter uses the output buffer on the ROM instance to
// hold data and drives rom_addr_o and data_vld_o to make a rdy/vld interface with the ROM output.
// This interface should signal things correctly until done_o goes high. data_last_nontop_o is set
// on the last word before the top RomTopCount words.
//

`include "prim_assert.sv"

module rom_ctrl_counter
  import prim_util_pkg::vbits;
#(
  parameter int RomDepth = 16,
  parameter int RomTopCount = 2
) (
  input                        clk_i,
  input                        rst_ni,

  output                       done_o,

  output [vbits(RomDepth)-1:0] read_addr_o,
  output                       read_req_o,

  output [vbits(RomDepth)-1:0] data_addr_o,

  input                        data_rdy_i,
  output                       data_last_nontop_o
);

  // The number of ROM entries that should be hashed. We assume there are at least 2, so that we can
  // register the data_last_nontop_o signal.
  localparam int RomNonTopCount = RomDepth - RomTopCount;

  `ASSERT_INIT(TopCountValid_A, 1 <= RomTopCount && RomTopCount < RomDepth)
  `ASSERT_INIT(NonTopCountValid_A, 2 <= RomNonTopCount)

  localparam int AW = vbits(RomDepth);

  localparam int unsigned TopAddrInt = RomDepth - 1;
  localparam int unsigned TNTAddrInt = RomNonTopCount - 2;

  localparam bit [AW-1:0] TopAddr = TopAddrInt[AW-1:0];
  localparam bit [AW-1:0] TNTAddr = TNTAddrInt[AW-1:0];

  logic          go;
  logic          req_q, vld_q;
  logic [AW-1:0] addr_q, addr_d;
  logic          done_q, done_d;
  logic          last_nontop_q, last_nontop_d;

  assign done_d = addr_q == TopAddr;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      done_q <= 1'b0;
    end else begin
      done_q <= done_d;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      addr_q        <= '0;
      last_nontop_q <= 1'b0;
    end else if (go) begin
      addr_q        <= addr_d;
      last_nontop_q <= last_nontop_d;
    end
  end

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      req_q <= 1'b0;
      vld_q <= 1'b0;
    end else begin
      // The first ROM request goes out immediately after reset (once we reach the top of ROM, we
      // signal done_o, after which the request signal is unused). We could clear it again when we
      // are done, but there's no need: the mux will switch away from us anyway.
      req_q <= 1'b1;

      // ROM data is valid from one cycle after the request goes out.
      vld_q <= req_q;
    end
  end

  assign go = data_rdy_i & vld_q & ~done_d;

  assign addr_d        = addr_q + {{AW-1{1'b0}}, 1'b1};
  assign last_nontop_d = addr_q == TNTAddr;

  assign done_o             = done_q;
  assign read_addr_o        = go ? addr_d : addr_q;
  assign read_req_o         = req_q;
  assign data_addr_o        = addr_q;
  assign data_last_nontop_o = last_nontop_q;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

//
// The ROM checker FSM module
//

`include "prim_assert.sv"

module rom_ctrl_fsm
  import prim_mubi_pkg::mubi4_t;
  import prim_util_pkg::vbits;
  import rom_ctrl_pkg::*;
#(
  parameter int RomDepth = 16,
  parameter int TopCount = 8
) (
  input logic                        clk_i,
  input logic                        rst_ni,

  // CSR inputs for DIGEST and EXP_DIGEST. To make the indexing look nicer, these are ordered so
  // that DIGEST_0 is the bottom 32 bits (they get reversed while we're shuffling around the wires
  // in rom_ctrl).
  input logic [TopCount*64-1:0]      digest_i,
  input logic [TopCount*64-1:0]      exp_digest_i,

  // CSR outputs for DIGEST and EXP_DIGEST. Ordered with word 0 as LSB.
  output logic [TopCount*64-1:0]     digest_o,
  output logic                       digest_vld_o,
  output logic [63:0]                exp_digest_o,
  output logic                       exp_digest_vld_o,
  output logic [vbits(TopCount)-1:0] exp_digest_idx_o,

  // To power manager and key manager
  output pwrmgr_data_t pwrmgr_data_o,
  output keymgr_data_t keymgr_data_o,

  // To KMAC (ROM data)
  input logic                        kmac_rom_rdy_i,
  output logic                       kmac_rom_vld_o,
  output logic                       kmac_rom_last_o,

  // To KMAC (digest data)
  input logic                        kmac_done_i,
  input logic [TopCount*64-1:0]      kmac_digest_i,
  input logic                        kmac_err_i,

  // To ROM mux
  output mubi4_t                     rom_select_bus_o,
  output logic [vbits(RomDepth)-1:0] rom_addr_o,
  output logic                       rom_req_o,

  // Raw bits from ROM
  input logic [63:0]                 rom_data_i,

  // To alert system
  output logic                       alert_o
);

  import prim_mubi_pkg::mubi4_test_true_loose;
  import prim_mubi_pkg::MuBi4False, prim_mubi_pkg::MuBi4True;

  localparam int AW = vbits(RomDepth);
  localparam int TAW = vbits(TopCount);

  localparam int unsigned TopStartAddrInt = RomDepth - TopCount;
  localparam bit [AW-1:0] TopStartAddr    = TopStartAddrInt[AW-1:0];

  // The counter / address generator
  logic          counter_done;
  logic [AW-1:0] counter_read_addr;
  logic          counter_read_req;
  logic [AW-1:0] counter_data_addr;
  logic          counter_data_rdy;
  logic          counter_lnt;
  rom_ctrl_counter #(
    .RomDepth (RomDepth),
    .RomTopCount (TopCount)
  ) u_counter (
    .clk_i              (clk_i),
    .rst_ni             (rst_ni),
    .done_o             (counter_done),
    .read_addr_o        (counter_read_addr),
    .read_req_o         (counter_read_req),
    .data_addr_o        (counter_data_addr),
    .data_rdy_i         (counter_data_rdy),
    .data_last_nontop_o (counter_lnt)
  );

  // The compare block (responsible for comparing CSR data and forwarding it to the key manager)
  logic   start_checker_q;
  logic   checker_done, checker_alert;
  mubi4_t checker_good;
  rom_ctrl_compare #(
    .NumWords  (TopCount)
  ) u_compare (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .start_i      (start_checker_q),
    .done_o       (checker_done),
    .good_o       (checker_good),
    .digest_i     (digest_i),
    .exp_digest_i (exp_digest_i),
    .alert_o      (checker_alert)
  );

  // Main FSM
  //
  // There are the following logical states
  //
  //    ReadingLow:   We're reading the low part of ROM and passing it to KMAC
  //    ReadingHigh:  We're reading the high part of ROM and waiting for KMAC
  //    RomAhead:     We've finished reading the high part of ROM, but are still waiting for KMAC
  //    KmacAhead:    KMAC is done, but we're still reading the high part of ROM
  //    Checking:     We are comparing DIGEST and EXP_DIGEST and sending data to keymgr
  //    Done:         Terminal state
  //    Invalid:      Terminal and invalid state (only reachable by a glitch)
  //
  // The FSM is linear, except for the branch where reading the high part of ROM races with getting
  // the result back from KMAC.
  //
  //     digraph fsm {
  //       ReadingLow -> ReadingHigh;
  //       ReadingHigh -> RomAhead;
  //       ReadingHigh -> KmacAhead;
  //       RomAhead -> Checking;
  //       KmacAhead -> Checking;
  //       Checking -> Done;
  //       Done [peripheries=2];
  //     }
  // SEC_CM: FSM.SPARSE
  // SEC_CM: INTERSIG.MUBI

  fsm_state_e state_d, state_q;
  logic       fsm_alert;

  `PRIM_FLOP_SPARSE_FSM(u_state_regs, state_d, state_q, fsm_state_e, ReadingLow)

  always_comb begin
    state_d = state_q;
    fsm_alert = 1'b0;

    unique case (state_q)
      ReadingLow: begin
        // Switch to ReadingHigh when counter_lnt is true and kmac_rom_rdy_i & kmac_rom_vld_o
        // (implying that the transaction went through)
        if (counter_lnt && kmac_rom_rdy_i && kmac_rom_vld_o) begin
          state_d = ReadingHigh;
        end
      end

      ReadingHigh: begin
        unique case ({kmac_done_i, counter_done})
          2'b01: state_d = RomAhead;
          2'b10: state_d = kmac_err_i ? Invalid : KmacAhead;
          2'b11: state_d = kmac_err_i ? Invalid : Checking;
          default: ; // No change
        endcase
      end

      RomAhead: begin
        if (kmac_done_i) state_d = kmac_err_i ? Invalid : Checking;
      end

      KmacAhead: begin
        if (counter_done) state_d = Checking;
      end

      Checking: begin
        if (checker_done) state_d = Done;
      end

      Done: begin
        // Final state
      end

      default: begin
        // An invalid state (includes the explicit Invalid state)
        fsm_alert = 1'b1;
        state_d = Invalid;
      end
    endcase

    // Consistency checks for done signals.
    //
    // If checker_done is high in a state other than Checking or Done then something has gone wrong
    // and we ran the check early. Similarly, counter_done should only be high after we've left
    // ReadingLow. Finally, kmac_done_i should only be high in ReadingHigh or RomAhead. If any of
    // these consistency requirements don't hold, jump to the Invalid state. This will also raise an
    // alert on the following cycle.
    //
    // SEC_CM: CHECKER.CTRL_FLOW.CONSISTENCY
    if ((checker_done && !(state_q inside {Checking, Done})) ||
        (counter_done && state_q == ReadingLow) ||
        (kmac_done_i && !(state_q inside {ReadingHigh, RomAhead}))) begin
      state_d = Invalid;
    end

    // Jump to an invalid state if sending out an alert for any other reason
    //
    // SEC_CM: CHECKER.FSM.LOCAL_ESC
    if (alert_o) begin
      state_d = Invalid;
    end
  end

  // The in_state_done signal is supposed to be true iff we're in FSM state Done. Grabbing just the
  // bottom 4 bits of state_q is equivalent to "mubi4_bool_to_mubi(state_q == Done)" except that it
  // doesn't have a 1-bit signal on the way.
  logic [9:0] state_q_bits;
  logic       unused_state_q_top_bits;
  assign state_q_bits = {state_q};
  assign unused_state_q_top_bits = ^state_q_bits[9:4];

  mubi4_t in_state_done;
  assign in_state_done = mubi4_t'(state_q_bits[3:0]);

  // Route digest signals coming back from KMAC straight to the CSRs
  assign digest_o     = kmac_digest_i;
  assign digest_vld_o = kmac_done_i;

  // Snoop on ROM reads to populate EXP_DIGEST, one word at a time
  logic reading_top;
  logic [AW-1:0] rel_addr_wide;
  logic [TAW-1:0] rel_addr;

  assign reading_top = (state_q == ReadingHigh || state_q == KmacAhead) & ~counter_done;
  assign rel_addr_wide = counter_data_addr - TopStartAddr;
  assign rel_addr = rel_addr_wide[TAW-1:0];

  // The top bits of rel_addr_wide should always be zero if we're reading the top bits (because TAW
  // bits should be enough to encode the difference between counter_data_addr and TopStartAddr)
  `ASSERT(RelAddrWide_A, exp_digest_vld_o |-> ~|rel_addr_wide[AW-1:TAW])
  logic unused_top_rel_addr_wide;
  assign unused_top_rel_addr_wide = |rel_addr_wide[AW-1:TAW];

  assign exp_digest_o = rom_data_i;
  assign exp_digest_vld_o = reading_top;
  assign exp_digest_idx_o = rel_addr;

  // The 'done' signal for pwrmgr is asserted once we get into the Done state. The 'good' signal
  // compes directly from the checker.
  assign pwrmgr_data_o = '{done: in_state_done, good: checker_good};

  // Pass the digest all-at-once to the keymgr. The loose check means that glitches will add
  // spurious edges to the valid signal that can be caught at the other end.
  assign keymgr_data_o = '{data: digest_i, valid: mubi4_test_true_loose(in_state_done)};

  // KMAC rom data interface
  logic kmac_rom_vld_d, kmac_rom_vld_q;
  always_comb begin
    // There will be valid data to pass to KMAC on each cycle after a counter request has gone out
    // when we were in state ReadingLow. That data goes out (causing us to drop the valid signal) if
    // KMAC was ready. Note that this formulation allows kmac_rom_vld_q to be high even if we're not
    // in the ReadingLow state: if something goes wrong and we get faulted into Invalid then we'll
    // still correctly send the end of the KMAC transaction.
    kmac_rom_vld_d = kmac_rom_vld_q;
    if (kmac_rom_rdy_i) begin
      kmac_rom_vld_d = 0;
    end
    if (counter_read_req && state_q == ReadingLow && !counter_lnt) begin
      kmac_rom_vld_d = 1;
    end
  end
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      kmac_rom_vld_q <= 0;
    end else begin
      kmac_rom_vld_q <= kmac_rom_vld_d;
    end
  end

  assign counter_data_rdy = kmac_rom_rdy_i | (state_q inside {ReadingHigh, KmacAhead});
  assign kmac_rom_vld_o = kmac_rom_vld_q;
  assign kmac_rom_last_o = counter_lnt;

  // The "last" flag is signalled when we're reading the last word in the first part of the ROM. As
  // a quick consistency check, this should only happen when the "valid" flag is also high.
  `ASSERT(LastImpliesValid_A, kmac_rom_last_o |-> kmac_rom_vld_o,
          clk_i, !rst_ni || (state_q == Invalid))

  // Start the checker when transitioning into the "Checking" state
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      start_checker_q <= 1'b0;
    end else begin
      start_checker_q <= (state_q != Checking) && (state_d == Checking);
    end
  end

  // The counter is supposed to run from zero up to the top of memory and then tell us that it's
  // done with the counter_done signal. We would like to be sure that no-one can fiddle with the
  // counter address once the hash has been computed (if they could subvert the mux as well, this
  // would allow them to generate a useful wrong address for a fetch). Fortunately, doing so would
  // cause the counter_done signal to drop again and we *know* that it should stay high when our FSM
  // is in the Done state.
  //
  // SEC_CM: CHECKER.CTR.CONSISTENCY
  logic unexpected_counter_change;
  assign unexpected_counter_change = mubi4_test_true_loose(in_state_done) & !counter_done;

  // We keep control of the ROM mux from reset until we're done.
  assign rom_select_bus_o = in_state_done;

  assign rom_addr_o = counter_read_addr;
  assign rom_req_o = counter_read_req;

  assign alert_o = fsm_alert | checker_alert | unexpected_counter_change;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

//
// The mux to select between ROM inputs
//

module rom_ctrl_mux
  import prim_mubi_pkg::mubi4_t;
#(
  parameter int AW = 8,
  parameter int DW = 39
) (
  input logic           clk_i,
  input logic           rst_ni,

  // Select signal saying whether access is granted to the bus. This module raises an alert (by
  // setting alert_o) if the signal isn't an allowed value or if the selection switches back from
  // the bus to the checker.
  input mubi4_t         sel_bus_i,

  // Interface for bus
  input logic [AW-1:0]  bus_rom_addr_i,
  input logic [AW-1:0]  bus_prince_addr_i,
  input logic           bus_req_i,
  output logic          bus_gnt_o,
  output logic [DW-1:0] bus_rdata_o,
  output logic          bus_rvalid_o,

  // Interface for ROM checker
  input logic [AW-1:0]  chk_addr_i,
  input logic           chk_req_i,
  output logic [DW-1:0] chk_rdata_o,

  // Interface for ROM
  output logic [AW-1:0] rom_rom_addr_o,
  output logic [AW-1:0] rom_prince_addr_o,
  output logic          rom_req_o,
  input logic [DW-1:0]  rom_scr_rdata_i,
  input logic [DW-1:0]  rom_clr_rdata_i,
  input logic           rom_rvalid_i,

  // Alert output
  //
  // This isn't latched in this module because it feeds into a fatal alert at top-level, whose
  // sender will latch it anyway.
  output logic          alert_o
);

  import prim_mubi_pkg::*;

  // Track the state of the mux up to the current cycle. This is a "1-way" mux, which means that
  // we never switch from the bus back to the checker.
  //
  // We also have a version that's delayed by a single cycle to allow a check that sel_bus_q is
  // never reset from True to False.
  logic [3:0] sel_bus_q_raw, sel_bus_qq_raw;
  mubi4_t     sel_bus_q, sel_bus_qq;

  prim_flop #(.Width (4), .ResetValue ({MuBi4False}))
  u_sel_bus_q_flop (
    .clk_i,
    .rst_ni,
    .d_i (mubi4_or_hi(sel_bus_q, sel_bus_i)),
    .q_o (sel_bus_q_raw)
  );
  assign sel_bus_q = mubi4_t'(sel_bus_q_raw);

  prim_flop #(.Width (4), .ResetValue ({MuBi4False}))
  u_sel_bus_qq_flop (
    .clk_i,
    .rst_ni,
    .d_i (sel_bus_q),
    .q_o (sel_bus_qq_raw)
  );
  assign sel_bus_qq = mubi4_t'(sel_bus_qq_raw);

  // Spot if the sel_bus_i signal or its register version has a corrupt value.
  //
  // SEC_CM: MUX.MUBI
  logic sel_invalid;
  assign sel_invalid = mubi4_test_invalid(sel_bus_i) || mubi4_test_invalid(sel_bus_q);

  // Spot if the select signal switches back to the checker once we've switched to the bus. Doing so
  // will have no lasting effect because of how we calculate sel_bus_q) but isn't supposed to
  // happen, so we want to trigger an alert.
  //
  // SEC_CM: MUX.CONSISTENCY
  logic sel_reverted;
  assign sel_reverted = mubi4_test_true_loose(sel_bus_q) & mubi4_test_false_loose(sel_bus_i);

  // Spot if the sel_bus_q signal has reverted somehow.
  //
  // SEC_CM: MUX.CONSISTENCY
  logic sel_q_reverted;
  assign sel_q_reverted = mubi4_test_true_loose(sel_bus_qq) & mubi4_test_false_loose(sel_bus_q);

  logic alert_q, alert_d;

  assign alert_d = sel_invalid | sel_reverted | sel_q_reverted;

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      alert_q <= 0;
    end else begin
      alert_q <= alert_q | alert_d;
    end
  end

  assign alert_o = alert_q;

  // The bus can have access every cycle, from when the select signal switches to the bus.
  assign bus_gnt_o    = mubi4_test_true_strict(sel_bus_i);
  assign bus_rdata_o  = rom_clr_rdata_i;
  // A high rom_rvalid_i is a response to a bus request if the select signal pointed at the bus on
  // the previous cycle.
  assign bus_rvalid_o = mubi4_test_true_strict(sel_bus_q) & rom_rvalid_i;

  assign chk_rdata_o = rom_scr_rdata_i;

  assign rom_req_o         = mubi4_test_true_strict(sel_bus_i) ? bus_req_i         : chk_req_i;
  assign rom_rom_addr_o    = mubi4_test_true_strict(sel_bus_i) ? bus_rom_addr_i    : chk_addr_i;
  assign rom_prince_addr_o = mubi4_test_true_strict(sel_bus_i) ? bus_prince_addr_i : chk_addr_i;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`include "prim_assert.sv"

//
// A scrambled ROM. This is scrambled with a fixed key, passed in as a parameter (this parameter
// will be a compile-time random constant).
//
// This code follows the structure of prim_ram_1p_scr.sv (although it's much simplified because the
// key is fixed and we don't support writes). For more information about what is going on, see that
// file. Using the parameter names in prim_ram_1p_scr, we have NumPrinceRoundsHalf = 2 (so
// approximately 5 effective rounds), NumDiffRounds = 2 and NumAddrScrRounds = 2 (enabling address
// scrambling with 2 rounds).
//
// There are two input address ports (rom_addr_i and prince_addr_i). These are expected to be
// connected to signals that are logically the same. The first is used as an input to the physical
// ROM index. The second is used when calculating the address-tweakable keystream. The trick is that
// you can mitigate fault-injection attacks that corrupt the address by splitting it somewhere
// "upstream". If a fault-injection only corrupts one of the two addresses, the result will be
// garbage.

module rom_ctrl_scrambled_rom
  import prim_rom_pkg::rom_cfg_t;
#(
  // The initial contents of the ROM. This is used for synthesis. For simulation, this is not used;
  // instead, the simulator loads the contents of ROM over DPI.
  //
  // In either case, the input file should be scrambled. That is, it should contain the bits that
  // will appear in the physical ROM.
  parameter MemInitFile = "",

  // The width of ROM words in bits
  parameter int Width = 40,

  // The number of words in the ROM
  parameter int Depth = 16,

  // The nonce for data and address scrambling
  parameter bit [63:0] ScrNonce = '0,

  // The (fixed) key for the PRINCE cipher
  parameter bit [127:0] ScrKey = '0,

  localparam int Aw = $clog2(Depth)
) (
  input logic              clk_i,
  input logic              rst_ni,

  input  logic             req_i,
  input  logic [Aw-1:0]    rom_addr_i,
  input  logic [Aw-1:0]    prince_addr_i,
  output logic             rvalid_o,
  output logic [Width-1:0] scr_rdata_o,
  output logic [Width-1:0] clr_rdata_o,

  input rom_cfg_t          cfg_i
);

  /////////////////////////////////////
  // Anchor incoming seeds and constants
  /////////////////////////////////////
  localparam int TotalAnchorWidth = $bits(ScrNonce) +
                                    $bits(ScrKey);

  logic [63:0] scr_nonce;
  logic [127:0] scr_key;

  prim_sec_anchor_buf #(
    .Width(TotalAnchorWidth)
  ) u_seed_anchor (
    .in_i({ScrNonce,
           ScrKey}),
    .out_o({scr_nonce,
            scr_key})
  );

  logic [63-Aw:0] data_scr_nonce;
  logic [Aw-1:0] addr_scr_nonce;
  assign data_scr_nonce = scr_nonce[63-Aw:0];
  assign addr_scr_nonce = scr_nonce[63-:Aw];

  // Parameter Checks ==========================================================

  // The depth needs to be a power of 2 to use address scrambling
  `ASSERT_INIT(DepthPow2Check_A, (Depth & (Depth - 1)) == 0)
  // We only support a width up to 64
  `ASSERT_INIT(MaxWidthCheck_A, Width <= 64)

  // Address scrambling ========================================================

  logic [Aw-1:0] addr_scr;
  prim_subst_perm #(
    .DataWidth (Aw),
    .NumRounds (2),
    .Decrypt   (0)
  ) u_sp_addr (
    .data_i (rom_addr_i),
    .key_i  (addr_scr_nonce),
    .data_o (addr_scr)
  );

  // Keystream generation ======================================================

  logic [63:0] keystream;

  prim_prince #(
    .DataWidth      (64),
    .KeyWidth       (128),
    .NumRoundsHalf  (2),
    .HalfwayDataReg (1'b1),
    .HalfwayKeyReg  (1'b1)
  ) u_prince (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),
    .valid_i (req_i),
    .data_i  ({data_scr_nonce, prince_addr_i}),
    .key_i   (scr_key),
    .dec_i   (1'b0),
    .data_o  (keystream),
    .valid_o ()
  );

  if (Width < 64) begin : gen_unread_keystream
    // Ignore top bits of keystream: we just use the bottom Width bits.
    logic unused_top_keystream;
    assign unused_top_keystream = ^keystream[63:Width];
  end

  // The physical ROM ==========================================================

  logic [Width-1:0] rdata_scr;

  prim_rom_adv #(
    .Width       (Width),
    .Depth       (Depth),
    .MemInitFile (MemInitFile)
  ) u_rom (
    .clk_i    (clk_i),
    .rst_ni   (rst_ni),
    .req_i    (req_i),
    .addr_i   (addr_scr),
    .rvalid_o (rvalid_o),
    .rdata_o  (rdata_scr),
    .cfg_i    (cfg_i)
  );

  assign scr_rdata_o = rdata_scr;

  // Data scrambling ===========================================================

  logic [Width-1:0] rdata_xor;

  prim_subst_perm #(
    .DataWidth (Width),
    .NumRounds (2),
    .Decrypt   (1)
  ) u_sp_data (
    .data_i (rdata_scr),
    .key_i  ('0),
    .data_o (rdata_xor)
  );

  // XOR rdata with keystream ==================================================

  assign clr_rdata_o = rdata_xor ^ keystream[Width-1:0];

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// ------------------- W A R N I N G: A U T O - G E N E R A T E D   C O D E !! -------------------//
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED WITH THE FOLLOWING COMMAND:
//
// util/topgen.py -t hw/top_earlgrey/data/top_earlgrey.hjson \
//                -o hw/top_earlgrey/ \
//                --rnd_cnst_seed 4881560218908238235


package top_earlgrey_rnd_cnst_rot_pkg;

  ////////////////////////////////////////////
  // otp_ctrl
  ////////////////////////////////////////////
  // Compile-time random bits for initial LFSR seed
  parameter otp_ctrl_pkg::lfsr_seed_t RndCnstOtpCtrlLfsrSeed = {
    40'hCB_0157A3AC
  };

  // Compile-time random permutation for LFSR output
  parameter otp_ctrl_pkg::lfsr_perm_t RndCnstOtpCtrlLfsrPerm = {
    240'h3946_DF803226_3D64E474_A1A11054_1E61A557_70D0A331_10222592_C19479D2
  };

  // Compile-time random permutation for scrambling key/nonce register reset value
  parameter otp_ctrl_pkg::scrmbl_key_init_t RndCnstOtpCtrlScrmblKeyInit = {
    256'h605FEFE9_977B00B6_FDC21D57_7A172D04_7DCF0EEB_BDD268AF_D4E2506D_F1D0603F
  };

  ////////////////////////////////////////////
  // lc_ctrl
  ////////////////////////////////////////////
  // Compile-time random bits for lc state group diversification value
  parameter lc_ctrl_pkg::lc_keymgr_div_t RndCnstLcCtrlLcKeymgrDivInvalid = {
    128'h9CD62F17_8ADC74D5_3D8AD0B6_00E7A1DD
  };

  // Compile-time random bits for lc state group diversification value
  parameter lc_ctrl_pkg::lc_keymgr_div_t RndCnstLcCtrlLcKeymgrDivTestDevRma = {
    128'h2F1A43C0_3DD4FF9B_887AB752_1CA6CBD8
  };

  // Compile-time random bits for lc state group diversification value
  parameter lc_ctrl_pkg::lc_keymgr_div_t RndCnstLcCtrlLcKeymgrDivProduction = {
    128'hD7107BAB_98B07574_3F7AEBA8_1E1C4EC8
  };

  // Compile-time random bits used for invalid tokens in the token mux
  parameter lc_ctrl_pkg::lc_token_mux_t RndCnstLcCtrlInvalidTokens = {
    256'hEBDEEE29_11062E03_9F8C7E1A_FA78A1D4_2886CC89_AE759CF8_65B22A5F_28DE2ECA,
    256'h36AFC2E8_A402302C_BDCF2B48_19AFAA0A_11CB6837_1EEF174D_98315696_C49A8EF5,
    256'h3C96F11E_4F43FFD4_21E456B4_D6A9D1D2_AB4A836F_1545EBF5_0FF87BC3_FE8473A3,
    256'hB8A698EB_44C3B582_1FC5BAE3_E1BD5972_3B69B2D7_B5330424_C30845EB_1F7A5EEF
  };

  ////////////////////////////////////////////
  // alert_handler
  ////////////////////////////////////////////
  // These LFSR parameters have been generated with
  // $ util/design/gen-lfsr-seed.py --width 32 --seed 2700182644
  localparam int LfsrWidth = 32;
  typedef logic [LfsrWidth-1:0]                        lfsr_seed_t;
  typedef logic [LfsrWidth-1:0][$clog2(LfsrWidth)-1:0] lfsr_perm_t;
  localparam lfsr_seed_t RndCnstLfsrSeedDefault = 32'he96064e5;
  localparam lfsr_perm_t RndCnstLfsrPermDefault =
      160'hebd1e5d4a1cee5afdb866a9c7a0278b899020d31;
  // Compile-time random bits for initial LFSR seed
  parameter lfsr_seed_t RndCnstAlertHandlerLfsrSeed = {
    32'h762A1F91
  };

  // Compile-time random permutation for LFSR output
  parameter lfsr_perm_t RndCnstAlertHandlerLfsrPerm = {
    160'h375ED89D_2A1D3286_2F7A7785_F940950C_C1CBDB05
  };

  ////////////////////////////////////////////
  // sram_ctrl_ret_aon
  ////////////////////////////////////////////
  // Compile-time random reset value for SRAM scrambling key.
  parameter otp_ctrl_pkg::sram_key_t RndCnstSramCtrlRetAonSramKey = {
    128'h3925A2B2_B291A984_70716274_C976B810
  };

  // Compile-time random reset value for SRAM scrambling nonce.
  parameter otp_ctrl_pkg::sram_nonce_t RndCnstSramCtrlRetAonSramNonce = {
    128'h6DD974CC_66D7F9C8_518EEFB7_5AC6B952
  };

  // Compile-time random bits for initial LFSR seed
  // parameter sram_ctrl_pkg::lfsr_seed_t RndCnstSramCtrlRetAonLfsrSeed = {
  //   32'h8242CE57
  // };

  // Compile-time random permutation for LFSR output
  // parameter sram_ctrl_pkg::lfsr_perm_t RndCnstSramCtrlRetAonLfsrPerm = {
  //   160'h9EB0A8F5_24A38F50_A1658338_21DF3607_BEF3365B
  // };

  ////////////////////////////////////////////
  // flash_ctrl
  ////////////////////////////////////////////
  // Compile-time random bits for default address key
  // parameter flash_ctrl_pkg::flash_key_t RndCnstFlashCtrlAddrKey = {
  //   128'h4B9E2FC1_918D324C_4CFB1A95_698EA1EB
  // };

  // // Compile-time random bits for default data key
  // parameter flash_ctrl_pkg::flash_key_t RndCnstFlashCtrlDataKey = {
  //   128'h7868F849_707838F5_47A2C2A6_4A91A9D7
  // };

  // Compile-time random bits for default seeds
  // parameter flash_ctrl_pkg::all_seeds_t RndCnstFlashCtrlAllSeeds = {
  //   256'h03429D8D_73DEDB65_D2B0751B_90255CCD_E50A2C9A_B31CAFB7_5C007285_A0AE495E,
  //   256'h2F5F51FD_2ACF2129_01174C95_76A112CE_A79B5228_2399833D_A888C025_46E72EB6
  // };

  // // Compile-time random bits for initial LFSR seed
  // parameter flash_ctrl_pkg::lfsr_seed_t RndCnstFlashCtrlLfsrSeed = {
  //   32'hF09A26A1
  // };

  // // Compile-time random permutation for LFSR output
  // parameter flash_ctrl_pkg::lfsr_perm_t RndCnstFlashCtrlLfsrPerm = {
  //   160'h8D51F377_9EA63579_4CE550B2_476E096B_C165846C
  // };

  ////////////////////////////////////////////
  // aes
  ////////////////////////////////////////////
  // Default seed of the PRNG used for register clearing.
  // parameter aes_pkg::clearing_lfsr_seed_t RndCnstAesClearingLfsrSeed = {
  //   64'h690709F0_9E8597D2
  // };

  // // Permutation applied to the LFSR of the PRNG used for clearing.
  // parameter aes_pkg::clearing_lfsr_perm_t RndCnstAesClearingLfsrPerm = {
  //   128'h18C91866_7BFD0701_C2E7C825_AD6C5429,
  //   256'h18C8E8BB_AA737B5F_CFB7A8A6_CD054048_BF9B54A1_4CFF8E69_DC8DE000_F65C955B
  // };

  // // Permutation applied to the clearing PRNG output for clearing the second share of registers.
  // parameter aes_pkg::clearing_lfsr_perm_t RndCnstAesClearingSharePerm = {
  //   128'hF8633CFD_E5AFA6B5_07549420_EAED688C,
  //   256'h110A9306_B63992EA_71787DC9_F634CC30_916F7B48_4A6E3195_D37BB278_8F153E40
  // };

  // // Default seed of the PRNG used for masking.
  // parameter aes_pkg::masking_lfsr_seed_t RndCnstAesMaskingLfsrSeed = {
  //   160'hEBDB78AA_E822F2F4_44DF087B_34854B57_FA1B481B
  // };

  // // Permutation applied to the concatenated LFSRs of the PRNG used for masking.
  // parameter aes_pkg::masking_lfsr_perm_t RndCnstAesMaskingLfsrPerm = {
  //   256'h35211013_03181580_8909584F_6726255D_0417556D_9E2A2273_41642E82_6136760C,
  //   256'h4E9B0616_931F514C_8D0B793D_66428130_37878800_20024950_2B68999D_0A6F864D,
  //   256'h4A94193F_54293A1A_63774685_2833577D_1C323974_9C0F2C05_31834027_1E705E1B,
  //   256'h758E453E_7B52906A_8C8A9848_5B11122F_622D083B_569A9153_781D9223_8F6E385F,
  //   256'h47957F96_4B847E24_7A726065_97597C3C_075A4371_6C0E5C69_340D8B44_6B14019F
  // };

  ////////////////////////////////////////////
  // kmac
  ////////////////////////////////////////////
  // Compile-time random data for LFSR default seed
  parameter kmac_pkg::lfsr_seed_t RndCnstKmacLfsrSeed = {
    32'h48F16180,
    256'h90982699_8ACE3628_C0CF0E58_B7088571_8609FA79_565DCBA5_40ADED8C_8D5560AF,
    256'h97340EA9_29AAE07C_399BB65D_74BD1FF1_6F281690_2BBE7ED5_4814F745_1C011AFB,
    256'hB712B66E_42C19103_58162E3F_B2368EBD_E95C97FA_3B0E8F66_29A16E94_D4E43991
  };

  // Compile-time random permutation for LFSR output
  parameter kmac_pkg::lfsr_perm_t RndCnstKmacLfsrPerm = {
    64'hC116F8EC_1BB4A423,
    256'h18778492_5ADD5D7F_1736506F_13C55AB6_AB1A7075_10497A2A_30AAF41D_15E7B06A,
    256'h0605324A_931E4CA2_06B335F1_26DC4205_9684F991_522E8483_09936099_5DB9A761,
    256'h86A6CB55_A44A6637_901577FC_4838501B_71F8534B_27EC9C6B_CF3C31AE_BCA3A810,
    256'h266D6010_89E99C92_C7CC3EBD_711A5036_8D938C71_D234E9E5_644C636E_E1AE0B88,
    256'hCE78281D_70E775FC_1EB389EB_C09F7C1D_1AD4052B_89680D14_11EE2B68_C35E576B,
    256'h91112650_C8FE9C0E_5371C1B1_6E89371E_5B48E601_7A5460A5_833A78AF_684C4E02,
    256'h9C1D62FA_5A2C4C98_468F60C2_09967AA8_276072C0_90C3B20F_1BAC1804_4271BC55,
    256'hA5CA5265_DDF621B0_6B5613D0_ACC0EE00_90A6904D_29992B4C_87F7D1D9_359DEB94,
    256'h8AB24825_91DAB12E_A3B060A1_4F1B144A_43DE23A1_7587C94B_B0118C6F_F38A6360,
    256'h5C998B17_1151D0CA_38BDC3C3_E1C0184C_F029215B_1A78E4A2_5014B29E_3042E567,
    256'h9EBB4D62_B791C625_E5F4787B_4B68A4D2_D0866A29_ADA8AC86_D280510C_D399D229,
    256'h7148CBAC_A4C39BD3_7C136EC3_56E1171B_8B7460FA_8800950E_886C8F79_D43A5B6F,
    256'hA9758987_9F779682_ABA5EC58_FD5C4D5A_FA47B36C_1AB24FB0_ED461EE3_13949320,
    256'hA8572862_24082384_6B223D9F_50263D66_411455E1_FE6FDEF8_74801A26_82100C5D,
    256'h1F92FCCC_3A8E56DA_4A2F6DD3_C22D052C_286D9214_8A11F66A_A345732D_530FD9C0,
    256'h0E3C3E69_6B9DCD43_44033698_A6E877F4_B3556330_06CC1726_49BDEDC7_4EBA68C1,
    256'h236D33C9_1531C9D0_E221820D_9219DDC0_A45781A0_A9E15A7C_AD53DC81_42FB8413,
    256'h00D1A693_269C3DCB_46A51AC4_070B2923_987A6122_45AA5CAF_DCC89AF3_4F53C666,
    256'h4B068DDB_5A2E054B_B26E8E0F_59F47D0E_B7C31762_A11C5937_E82FADAB_A4A98B41,
    256'h82D37190_AD21A858_2383E7C7_C6172E81_F9EE6E21_64675464_9547336E_35619128,
    256'hD0AA1DAA_4A418549_C5A3D9E1_7DAFE195_22459691_12227A93_679A0006_5DC9B103,
    256'hBF4EF30A_4E6FA1CB_854C7ADD_0A552FB9_8954E9DB_6CD96BBE_B9B1F081_E00D5954,
    256'hA1756301_05F5ED3B_7D71E085_09685F24_9300A00D_09B6D94B_946C695B_B5706C06,
    256'hA866273B_B55F134D_19FCB953_99B46EBC_1D53F240_8B09417A_E0665515_04203018,
    256'hDA29406C_02E5919E_0EB185BC_41D789D9_E3A57C8C_B1410E89_21D29C54_E0244E4C,
    256'h611C0DE8_16AE9798_6AFC6459_A2C5681D_B48357E7_38B02F1D_3104AF12_D58415A4,
    256'h712D138C_FE70570B_3E0C8F96_E2D41049_89A0BA28_AA5A55F4_7C0A47E2_21AC2AE2,
    256'h544D6281_48FB29E3_C2D6B59C_02819412_E1EE5DC7_2545193F_EA567542_369473B4,
    256'hD8638274_A22F162D_B6A8C0AA_8B48B249_9230A188_DEBA5607_3DBC94D0_0B61C266,
    256'h8B63F0A9_9E454000_2B750F58_4E8368E6_7B5C064C_C98A3131_3B8D4A46_A628EFC6,
    256'h3214C371_F7282854_AF8B797A_41CC5629_95038A5C_14128AA7_E03EF942_AF63ECC4
  };

  // Compile-time random permutation for forwarding LFSR state
  parameter kmac_pkg::lfsr_fwd_perm_t RndCnstKmacLfsrFwdPerm = {
    160'h6C52BADA_026047A3_4F972E09_20768872_9FBCF8FF
  };

  // Compile-time random permutation for LFSR Message output
  parameter kmac_pkg::msg_perm_t RndCnstKmacMsgPerm = {
    128'hE16CB1A4_455785BD_0DC24673_FD21EADF,
    256'hE99C19F0_E0090DAF_78E94915_8B4C20F8_EE8944FB_00A9FA45_D07D2F5A_3CB2B6B9
  };

  ////////////////////////////////////////////
  // otbn
  ////////////////////////////////////////////
  // Default seed of the PRNG used for URND.
  parameter otbn_pkg::urnd_prng_seed_t RndCnstOtbnUrndPrngSeed = {
    256'h173B0217_51142EB3_0B9482BD_8E7D31D3_E1A2619D_66EF6CB9_16FD6C86_4A510AED
  };

  // Compile-time random reset value for IMem/DMem scrambling key.
  parameter otp_ctrl_pkg::otbn_key_t RndCnstOtbnOtbnKey = {
    128'h83D2D2E2_4871C35E_3AEABAE7_7182CDEF
  };

  // Compile-time random reset value for IMem/DMem scrambling nonce.
  parameter otp_ctrl_pkg::otbn_nonce_t RndCnstOtbnOtbnNonce = {
    64'hF9F77516_F1177315
  };

  ////////////////////////////////////////////
  // keymgr
  ////////////////////////////////////////////
  // Compile-time random bits for initial LFSR seed
  parameter keymgr_pkg::lfsr_seed_t RndCnstKeymgrLfsrSeed = {
    64'h733AFFA7_32F4C491
  };

  // Compile-time random permutation for LFSR output
  parameter keymgr_pkg::lfsr_perm_t RndCnstKeymgrLfsrPerm = {
    128'h2C629940_F4ED827C_37884C63_AA6A4E74,
    256'h55EC93C2_1BB87712_ED5D4CA1_E274C8DD_B953F0FE_03A46F59_8AC1E1A0_9FCFD865
  };

  // Compile-time random permutation for entropy used in share overriding
  parameter keymgr_pkg::rand_perm_t RndCnstKeymgrRandPerm = {
    160'h5216C347_ED2DE7AA_0BD0C6EB_D905EEB7_3203A483
  };

  // Compile-time random bits for revision seed
  parameter keymgr_pkg::seed_t RndCnstKeymgrRevisionSeed = {
    256'h414C190A_D0A09D14_4FFC0C0F_EA081CEF_945B641F_096B9F3E_9A494BA3_5FCFEF0D
  };

  // Compile-time random bits for creator identity seed
  parameter keymgr_pkg::seed_t RndCnstKeymgrCreatorIdentitySeed = {
    256'hFB223E8A_B704F249_EE3FA822_276C45E5_88ED40CF_52C8FAE2_D054A711_49771822
  };

  // Compile-time random bits for owner intermediate identity seed
  parameter keymgr_pkg::seed_t RndCnstKeymgrOwnerIntIdentitySeed = {
    256'h2EC37360_E23D4DDA_559ADABC_F099937F_EBBF048F_AC328BA1_BDEE0CAC_A987BE4A
  };

  // Compile-time random bits for owner identity seed
  parameter keymgr_pkg::seed_t RndCnstKeymgrOwnerIdentitySeed = {
    256'h4ABF486B_16740B20_BC32B13F_F07A13FF_21CE605E_0AC01985_8F73D707_CD0EC1D3
  };

  // Compile-time random bits for software generation seed
  parameter keymgr_pkg::seed_t RndCnstKeymgrSoftOutputSeed = {
    256'h3DAAEF20_E285FA65_8FDD1B42_6C037151_B16C8D44_4C444F39_6F4479CB_795CF94B
  };

  // Compile-time random bits for hardware generation seed
  parameter keymgr_pkg::seed_t RndCnstKeymgrHardOutputSeed = {
    256'h9E409D18_381BD5D5_6821E298_5E479971_05C4900F_25557467_5985B210_E1A968E4
  };

  // Compile-time random bits for generation seed when aes destination selected
  parameter keymgr_pkg::seed_t RndCnstKeymgrAesSeed = {
    256'h5E5B35E4_60FDAF1F_F382AB01_95E33689_D99BCEBF_2B79B683_9264EDF4_DE2B39F3
  };

  // Compile-time random bits for generation seed when kmac destination selected
  parameter keymgr_pkg::seed_t RndCnstKeymgrKmacSeed = {
    256'h94059891_A38BD1D1_6C763BBD_90347E58_152D7FCA_99380365_25AAA3F8_9E3DE8F1
  };

  // Compile-time random bits for generation seed when otbn destination selected
  parameter keymgr_pkg::seed_t RndCnstKeymgrOtbnSeed = {
    256'h278645E1_1D7CAC76_310205E1_9CD3F2ED_294A279F_3C6D0649_A905CC9B_10A67A16
  };

  // Compile-time random bits for generation seed when no CDI is selected
  parameter keymgr_pkg::seed_t RndCnstKeymgrCdi = {
    256'h161FED72_416DFD29_3DE3A18A_8837B0DD_4CB694DD_540451D7_69D28E1D_9E76007B
  };

  // Compile-time random bits for generation seed when no destination selected
  parameter keymgr_pkg::seed_t RndCnstKeymgrNoneSeed = {
    256'h7A9E0F6E_3D591A7F_D8C7BA26_4AF78F28_AEE0D28E_4D638D95_D1806E87_0336CD96
  };

  ////////////////////////////////////////////
  // csrng
  ////////////////////////////////////////////
  // Compile-time random bits for csrng state group diversification value
  parameter csrng_pkg::cs_keymgr_div_t RndCnstCsrngCsKeymgrDivNonProduction = {
    128'h1D2049F3_32011CAB_7D512B69_B6B766DC,
    256'h84760801_C9AAE19E_8A6DD42F_94A9A15F_A77F118B_21BA52C5_D59D755F_58D2D862
  };

  // Compile-time random bits for csrng state group diversification value
  parameter csrng_pkg::cs_keymgr_div_t RndCnstCsrngCsKeymgrDivProduction = {
    128'h44D2DC25_8CA12CC7_0B776B16_DD95013B,
    256'h9569BD77_059093ED_3CE77AEA_86FFD82C_B1CDEE3F_CD6039C7_C0402496_5B7C1E1C
  };

  ////////////////////////////////////////////
  // sram_ctrl_main
  ////////////////////////////////////////////
  // Compile-time random reset value for SRAM scrambling key.
  parameter otp_ctrl_pkg::sram_key_t RndCnstSramCtrlMainSramKey = {
    128'h07548A9B_F5956E74_82848DE7_D401512A
  };

  // Compile-time random reset value for SRAM scrambling nonce.
  parameter otp_ctrl_pkg::sram_nonce_t RndCnstSramCtrlMainSramNonce = {
    128'h2573043A_8E0AD9B1_56D761AD_532F38F0
  };

  // // Compile-time random bits for initial LFSR seed
  // parameter sram_ctrl_pkg::lfsr_seed_t RndCnstSramCtrlMainLfsrSeed = {
  //   32'h767AFF4B
  // };

  // // Compile-time random permutation for LFSR output
  // parameter sram_ctrl_pkg::lfsr_perm_t RndCnstSramCtrlMainLfsrPerm = {
  //   160'h6CD8E170_15D40914_D8A70990_BFF77996_28F1F957
  // };

  ////////////////////////////////////////////
  // rom_ctrl
  ////////////////////////////////////////////
  // Fixed nonce used for address / data scrambling
  parameter bit [63:0] RndCnstRomCtrlScrNonce = {
    64'h755CF00B_D7432C3F
  };

  // Randomised constant used as a scrambling key for ROM data
  parameter bit [127:0] RndCnstRomCtrlScrKey = {
    128'h8CD4E7EF_F1B9EC59_CE812447_C5714595
  };

  ////////////////////////////////////////////
  // rv_core_ibex
  ////////////////////////////////////////////
  // Default seed of the PRNG used for random instructions.
  // parameter ibex_pkg::lfsr_seed_t RndCnstRvCoreIbexLfsrSeed = {
  //   32'hF17463DB
  // };

  // // Permutation applied to the LFSR of the PRNG used for random instructions.
  // parameter ibex_pkg::lfsr_perm_t RndCnstRvCoreIbexLfsrPerm = {
  //   160'h7D3352C5_76E13E90_EFC895C1_36094776_203E9B4D
  // };

  // // Default icache scrambling key
  // parameter logic [ibex_pkg::SCRAMBLE_KEY_W-1:0] RndCnstRvCoreIbexIbexKeyDefault = {
  //   128'hC10D8DD7_F82D1584_4E53A6AF_23823858
  // };

  // // Default icache scrambling nonce
  // parameter logic [ibex_pkg::SCRAMBLE_NONCE_W-1:0] RndCnstRvCoreIbexIbexNonceDefault = {
  //   64'h2F4520C3_2D5E0D6D
  // };

endpackage : top_earlgrey_rnd_cnst_rot_pkg



`include "prim_assert.sv"

module rot_top #(
  // parameters for hmac
  // parameters for kmac
  parameter bit KmacEnMasking = 1,
  parameter bit KmacSwKeyMasked = 0,
  parameter int SecKmacCmdDelay = 0,
  parameter bit SecKmacIdleAcceptSwMsg = 0,
  // parameters for keymgr
  parameter bit KeymgrKmacEnMasking = 1,
  // parameters for rom_ctrl
  parameter RomCtrlBootRomInitFile = "/nfs/home/zhangdongrong/Desktop/tmp/Nanhu-V3-main/src/main/resources/TLROT/test.vmem",
  parameter bit SecRomCtrlDisableScrambling = 1'b0,
  // parameters for csrng
  parameter aes_pkg::sbox_impl_e CsrngSBoxImpl = aes_pkg::SBoxImplCanright,
  // parameters for entropy_src
  parameter int EntropySrcEsFifoDepth = 4,
  parameter bit EntropySrcStub = 0,
  // parameters for edn0
  // parameters for otbn
  parameter bit OtbnStub = 0,
  parameter otbn_pkg::regfile_e OtbnRegFile = otbn_pkg::RegFileFF,
  parameter bit SecOtbnMuteUrnd = 0,
  parameter bit SecOtbnSkipUrndReseedAtStart = 0,
  // alert
  parameter logic [14-1:0] AlertAsyncOn = {14{1'b1}}
) (
    input clk_i,
    input rst_ni,
    input rst_shadowed_ni,
    input clk_edn_i,
    input rst_edn_ni,
    input scan_mode,

    // Bus Interface
    input  tlul_pkg::tl_h2d_t tl_i,
    output tlul_pkg::tl_d2h_t tl_o,

    // Interrupt
    output logic intr_hmac_hmac_done_o,
    output logic intr_hmac_fifo_empty_o,
    output logic intr_hmac_hmac_err_o,
    output logic intr_kmac_kmac_done_o,
    output logic intr_kmac_fifo_empty_o,
    output logic intr_kmac_kmac_err_o,
    output logic intr_keymgr_op_done_o,
    output logic intr_csrng_cs_cmd_req_done_o,
    output logic intr_csrng_cs_entropy_req_o,
    output logic intr_csrng_cs_hw_inst_exc_o,
    output logic intr_csrng_cs_fatal_err_o,
    output logic intr_entropy_src_es_entropy_valid_o,
    output logic intr_entropy_src_es_health_test_failed_o,
    output logic intr_entropy_src_es_observe_fifo_ready_o,
    output logic intr_entropy_src_es_fatal_err_o,
    output logic intr_edn0_edn_cmd_req_done_o,
    output logic intr_edn0_edn_fatal_err_o,
    // output logic intr_otbn_done,

    // key output
    // output keymgr_pkg::hw_key_req_t       keymgr_aes_key,
    // output keymgr_pkg::hw_key_req_t       keymgr_kmac_key,
    // output keymgr_pkg::otbn_key_req_t       keymgr_otbn_key,
    input [255:0] key0,
    input logic key_valid,

    // entropy src
    output entropy_src_pkg::entropy_src_rng_req_t       es_rng_req_o,
    input entropy_src_pkg::entropy_src_rng_rsp_t       es_rng_rsp_i,
    // input prim_mubi_pkg::mubi8_t       entropy_src_otp_en_entropy_src_fw_read,
    // input prim_mubi_pkg::mubi8_t       entropy_src_otp_en_entropy_src_fw_over,
    output logic       es_rng_fips_o, 
    // input tlul_pkg::tl_h2d_t       entropy_src_tl_req,
    // output tlul_pkg::tl_d2h_t       entropy_src_tl_rsp,

    // rom
    // input kmac_pkg::app_rsp_t kmac_app_rsp_rom,
    // output kmac_pkg::app_req_t kmac_app_req_rom,
    output rom_ctrl_pkg::pwrmgr_data_t       rom_ctrl_pwrmgr_data,
    // input prim_rom_pkg::rom_cfg_t       ast_rom_cfg,
    input tlul_pkg::tl_h2d_t64 rom_ctrl_rom_tl_req,
    output tlul_pkg::tl_d2h_t64 rom_ctrl_rom_tl_rsp

    // kmac
    // output kmac_pkg::app_rsp_t kmac_app_rsp_lc,
    // input kmac_pkg::app_req_t kmac_app_req_lc,
    // output prim_mubi_pkg::mubi4_t  clkmgr_aon_idle_rot,

    //csrng
    // input csrng_pkg::csrng_req_t  rot_top_csrng_csrng_cmd_req,
    // output csrng_pkg::csrng_rsp_t  rot_top_csrng_csrng_cmd_rsp,
    // input csrng_pkg::csrng_req_t [1:0] csrng_csrng_cmd_req,
    // output csrng_pkg::csrng_rsp_t [1:0]  csrng_csrng_cmd_rsp,
    // input prim_mubi_pkg::mubi8_t       csrng_otp_en_csrng_sw_app_read,
    // input lc_ctrl_pkg::lc_tx_t lc_ctrl_lc_hw_debug_en,
    // input tlul_pkg::tl_h2d_t       csrng_tl_req,
    // output tlul_pkg::tl_d2h_t       csrng_tl_rsp,

    //edn0
    // output edn_pkg::edn_req_t edn0_edn_req_rot,
    // input edn_pkg::edn_rsp_t edn0_edn_rsp_rot,
    // input edn_pkg::edn_req_t [7:0] edn0_edn_req,
    // output edn_pkg::edn_rsp_t [7:0] edn0_edn_rsp,
    // input tlul_pkg::tl_h2d_t       edn0_tl_req,
    // output tlul_pkg::tl_d2h_t       edn0_tl_rsp,

    //otbn
    // input prim_ram_1p_pkg::ram_1p_cfg_t       ast_ram_1p_cfg,
    // output otp_ctrl_pkg::otbn_otp_key_req_t       otp_ctrl_otbn_otp_key_req,
    // input otp_ctrl_pkg::otbn_otp_key_rsp_t       otp_ctrl_otbn_otp_key_rsp,
    // input lc_ctrl_pkg::lc_tx_t       flash_ctrl_rma_ack,
    // output lc_ctrl_pkg::lc_tx_t       otbn_lc_rma_ack,

    // alerts NAlerts = 14
    // input  prim_alert_pkg::alert_rx_t [14-1:0] alert_rx_i,
    // output prim_alert_pkg::alert_tx_t [14-1:0] alert_tx_o
);

  import tlul_pkg::*;
  import top_pkg::*;
  // Compile-time random constants
  import top_earlgrey_rnd_cnst_rot_pkg::*;

  //local parameter
  

  // Signals
  //tlul signle
  tlul_pkg::tl_h2d_t       hmac_tl_req;
  tlul_pkg::tl_d2h_t       hmac_tl_rsp;
  tlul_pkg::tl_h2d_t       kmac_tl_req;
  tlul_pkg::tl_d2h_t       kmac_tl_rsp;
  tlul_pkg::tl_h2d_t       entropy_src_tl_req;
  tlul_pkg::tl_d2h_t       entropy_src_tl_rsp;
  tlul_pkg::tl_h2d_t       csrng_tl_req;
  tlul_pkg::tl_d2h_t       csrng_tl_rsp;
  tlul_pkg::tl_h2d_t       edn0_tl_req;
  tlul_pkg::tl_d2h_t       edn0_tl_rsp;
  tlul_pkg::tl_h2d_t       keymgr_tl_req;
  tlul_pkg::tl_d2h_t       keymgr_tl_rsp;
  // tlul_pkg::tl_h2d_t       rom_ctrl_rom_tl_req;
  // tlul_pkg::tl_d2h_t       rom_ctrl_rom_tl_rsp;
  tlul_pkg::tl_h2d_t       rom_ctrl_regs_tl_req;
  tlul_pkg::tl_d2h_t       rom_ctrl_regs_tl_rsp;
  tlul_pkg::tl_h2d_t       otbn_tl_req;
  tlul_pkg::tl_d2h_t       otbn_tl_rsp;
  tlul_pkg::tl_h2d_t       sm3_tl_req;
  tlul_pkg::tl_d2h_t       sm3_tl_rsp;
  tlul_pkg::tl_h2d_t       sm4_tl_req;
  tlul_pkg::tl_d2h_t       sm4_tl_rsp;
  tlul_pkg::tl_h2d_t       rs_encode_tl_req;
  tlul_pkg::tl_d2h_t       rs_encode_tl_rsp;
  tlul_pkg::tl_h2d_t       rs_decode_tl_req;
  tlul_pkg::tl_d2h_t       rs_decode_tl_rsp;
  tlul_pkg::tl_h2d_t       puf_tl_req;
  tlul_pkg::tl_d2h_t       puf_tl_rsp;
  tlul_pkg::tl_h2d_t       puf2_tl_req;
  tlul_pkg::tl_d2h_t       puf2_tl_rsp;


  // Alert list
  localparam NAlerts = 14;
  prim_alert_pkg::alert_tx_t [NAlerts-1:0]  alert_tx_o;
  // prim_alert_pkg::alert_rx_t [NAlerts-1:0]  alert_rx;
  localparam prim_alert_pkg::alert_rx_t [NAlerts-1:0] alert_rx_i = {NAlerts{prim_alert_pkg::ALERT_RX_DEFAULT}};

  
  // Interrupt source list
  // logic [16:0]  intr_vector;
  // logic  unused_intr_vector;
  // logic intr_hmac_hmac_done;
  // logic intr_hmac_fifo_empty;
  // logic intr_hmac_hmac_err;
  // logic intr_kmac_kmac_done;
  // logic intr_kmac_fifo_empty;
  // logic intr_kmac_kmac_err;
  // logic intr_keymgr_op_done;
  // logic intr_csrng_cs_cmd_req_done;
  // logic intr_csrng_cs_entropy_req;
  // logic intr_csrng_cs_hw_inst_exc;
  // logic intr_csrng_cs_fatal_err;
  // logic intr_entropy_src_es_entropy_valid;
  // logic intr_entropy_src_es_health_test_failed;
  // logic intr_entropy_src_es_observe_fifo_ready;
  // logic intr_entropy_src_es_fatal_err;
  // logic intr_edn0_edn_cmd_req_done;
  // logic intr_edn0_edn_fatal_err;
  logic intr_otbn_done;

  // define inter-module signal
  prim_mubi_pkg::mubi4_t [2:0] clkmgr_aon_idle;
  logic unused_clkmgr_aon_idle;
  assign unused_clkmgr_aon_idle = ^ clkmgr_aon_idle;

  // localparam  kmac_pkg::lc_tx_t       lc_ctrl_lc_escalate_en = kmac_pkg::LC_TX_DEFAULT;
  localparam  lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_escalate_en = lc_ctrl_pkg::Off;

  //Keymgr
  // edn_pkg::edn_req_t [1:0] edn0_edn_req;
  // edn_pkg::edn_rsp_t [1:0] edn0_edn_rsp;
  otp_ctrl_pkg::otp_keymgr_key_t       otp_ctrl_otp_keymgr_key;
  // otp_ctrl_pkg::otp_device_id_t       keymgr_otp_device_id;
  // localparam otp_ctrl_pkg::otp_keymgr_key_t otp_ctrl_otp_keymgr_key = otp_ctrl_pkg::OTP_KEYMGR_KEY_DEFAULT;
  assign otp_ctrl_otp_keymgr_key.key_share1 = otp_ctrl_pkg::OTP_KEYMGR_KEY_DEFAULT.key_share1;
  assign otp_ctrl_otp_keymgr_key.key_share0 = key0;
  assign otp_ctrl_otp_keymgr_key.valid = key_valid;
  localparam otp_ctrl_pkg::otp_device_id_t keymgr_otp_device_id = 256'h48ecf6c738f0f108a5b08620695ffd4d48ecf6c738f0f108a5b08620695ffd4d;
  keymgr_pkg::hw_key_req_t       keymgr_aes_key;
  logic unused_keymgr_aes_key;
  assign unused_keymgr_aes_key = ^ keymgr_aes_key;
  keymgr_pkg::hw_key_req_t       keymgr_kmac_key;
  keymgr_pkg::otbn_key_req_t       keymgr_otbn_key;
  kmac_pkg::app_req_t [2:0] kmac_app_req;
  // assign kmac_app_req[1] = kmac_pkg::APP_REQ_DEFAULT;
  kmac_pkg::app_rsp_t [2:0] kmac_app_rsp;
  // assign kmac_app_rsp[1] = kmac_pkg::APP_RSP_DEFAULT;
  logic       kmac_en_masking;
  // flash_ctrl_pkg::keymgr_flash_t       flash_ctrl_keymgr;
  // localparam keymgr_pkg::keymgr_flash_t flash_ctrl_keymgr = keymgr_pkg::KEYMGR_FLASH_DEFAULT;
  localparam flash_ctrl_pkg::keymgr_flash_t flash_ctrl_keymgr = flash_ctrl_pkg::KEYMGR_FLASH_DEFAULT;

  // lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_keymgr_en;
  // lc_ctrl_pkg::lc_keymgr_div_t       lc_ctrl_lc_keymgr_div;
  localparam lc_ctrl_pkg::lc_tx_t lc_ctrl_lc_keymgr_en = lc_ctrl_pkg::On;
  localparam lc_ctrl_pkg::lc_keymgr_div_t lc_ctrl_lc_keymgr_div = 128'h48aaf6c738f0f108a5b08620695ffd4d;
  rom_ctrl_pkg::keymgr_data_t       rom_ctrl_keymgr_data;
  // localparam rom_ctrl_pkg::keymgr_data_t rom_ctrl_keymgr_data = rom_ctrl_pkg::ROM_KEYMGR_DATA_DEFAULT;

  //ROM
  // prim_rom_pkg::rom_cfg_t       ast_rom_cfg;
  localparam prim_rom_pkg::rom_cfg_t       ast_rom_cfg = prim_rom_pkg::ROM_CFG_DEFAULT;
  // rom_ctrl_pkg::pwrmgr_data_t       rom_ctrl_pwrmgr_data;
  // logic       unused_rom_ctrl_pwrmgr_data;
  // assign unused_rom_ctrl_pwrmgr_data = ^ rom_ctrl_pwrmgr_data;
  // rom_ctrl_pkg::keymgr_data_t       rom_ctrl_keymgr_data;

  //csrng
  csrng_pkg::csrng_req_t [1:0]  csrng_csrng_cmd_req;
  assign csrng_csrng_cmd_req[1] = '0;
  csrng_pkg::csrng_rsp_t [1:0] csrng_csrng_cmd_rsp;
  // prim_mubi_pkg::mubi8_t       csrng_otp_en_csrng_sw_app_read;
  localparam  MuBi8False = 8'h69;
  localparam prim_mubi_pkg::mubi8_t       csrng_otp_en_csrng_sw_app_read = prim_mubi_pkg::mubi8_t'(MuBi8False);
  // lc_ctrl_pkg::lc_tx_t       lc_ctrl_lc_hw_debug_en;
  localparam lc_ctrl_pkg::lc_tx_t lc_ctrl_lc_hw_debug_en = lc_ctrl_pkg::On;

    // EDN0
  edn_pkg::edn_req_t [7:0] edn0_edn_req_intr;
  edn_pkg::edn_rsp_t [7:0] edn0_edn_rsp_intr;

  //entropy src
  entropy_src_pkg::entropy_src_hw_if_req_t       csrng_entropy_src_hw_if_req;
  entropy_src_pkg::entropy_src_hw_if_rsp_t       csrng_entropy_src_hw_if_rsp;
  entropy_src_pkg::cs_aes_halt_req_t       csrng_cs_aes_halt_req;
  entropy_src_pkg::cs_aes_halt_rsp_t       csrng_cs_aes_halt_rsp;
  // entropy_src_pkg::entropy_src_rng_req_t       es_rng_req_o;
  entropy_src_pkg::entropy_src_rng_rsp_t       es_rng_rsp_i_puf;
  // localparam entropy_src_pkg::entropy_src_rng_rsp_t       es_rng_rsp_i = entropy_src_pkg::ENTROPY_SRC_RNG_RSP_DEFAULT; 
  // prim_mubi_pkg::mubi8_t       entropy_src_otp_en_entropy_src_fw_read;
  // prim_mubi_pkg::mubi8_t       entropy_src_otp_en_entropy_src_fw_over;
  localparam prim_mubi_pkg::mubi8_t       entropy_src_otp_en_entropy_src_fw_read = prim_mubi_pkg::mubi8_t'(MuBi8False);
  localparam prim_mubi_pkg::mubi8_t       entropy_src_otp_en_entropy_src_fw_over = prim_mubi_pkg::mubi8_t'(MuBi8False);
  // logic       es_rng_fips_o;

  // otbn
  localparam prim_ram_1p_pkg::ram_1p_cfg_t       ast_ram_1p_cfg = prim_ram_1p_pkg::RAM_1P_CFG_DEFAULT;
  otp_ctrl_pkg::otbn_otp_key_req_t       otp_ctrl_otbn_otp_key_req;
  otp_ctrl_pkg::otbn_otp_key_rsp_t       otp_ctrl_otbn_otp_key_rsp;
  localparam lc_ctrl_pkg::lc_tx_t       flash_ctrl_rma_ack = lc_ctrl_pkg::LC_TX_DEFAULT;
  lc_ctrl_pkg::lc_tx_t       otbn_lc_rma_ack;

  // puf
  logic [3:0] rng4bit;
  logic rng4bit_done;
  logic rng_mode;

  // sinterrupt assignments
  // assign intr_vector = {
  //   intr_hmac_hmac_done,
  //   intr_hmac_fifo_empty,
  //   intr_hmac_hmac_err,
  //   intr_kmac_kmac_done,
  //   intr_kmac_fifo_empty,
  //   intr_kmac_kmac_err,
  //   intr_keymgr_op_done,
  //   intr_edn0_edn_cmd_req_done,
  //   intr_edn0_edn_fatal_err,
  //   intr_entropy_src_es_fatal_err, 
  //   intr_entropy_src_es_observe_fifo_ready, 
  //   intr_entropy_src_es_health_test_failed, 
  //   intr_entropy_src_es_entropy_valid, 
  //   intr_csrng_cs_fatal_err, 
  //   intr_csrng_cs_hw_inst_exc, 
  //   intr_csrng_cs_entropy_req, 
  //   intr_csrng_cs_cmd_req_done
  // };

  // assign unused_intr_vector = ^ intr_vector;

  assign kmac_app_req[2] = kmac_pkg::APP_REQ_DEFAULT;
  
  // assign kmac_app_rsp_lc = kmac_app_rsp[2]; 

  // assign csrng_csrng_cmd_req[1] = rot_top_csrng_csrng_cmd_req;
  // assign rot_top_csrng_csrng_cmd_rsp = csrng_csrng_cmd_rsp[1];

  assign edn0_edn_req_intr[1] = '0;
  assign edn0_edn_req_intr[2] = '0;
  assign edn0_edn_req_intr[4] = '0;
  // assign edn0_edn_req_intr[5] = edn0_edn_req[5];
  // assign edn0_edn_req_intr[6] = edn0_edn_req[6];
  assign edn0_edn_req_intr[7] = '0;

  // assign edn0_edn_rsp[1] = edn0_edn_rsp_intr[1];
  // assign edn0_edn_rsp[2] = edn0_edn_rsp_intr[2];
  // assign edn0_edn_rsp[4] = edn0_edn_rsp_intr[4];
  // // assign edn0_edn_rsp[5] = edn0_edn_rsp_intr[5];
  // // assign edn0_edn_rsp[6] = edn0_edn_rsp_intr[6];
  // assign edn0_edn_rsp[7] = edn0_edn_rsp_intr[7];

  hmac #(
    .AlertAsyncOn(1'b1)
  ) u_hmac (

      // Interrupt
      .intr_hmac_done_o  (intr_hmac_hmac_done_o),
      .intr_fifo_empty_o (intr_hmac_fifo_empty_o),
      .intr_hmac_err_o   (intr_hmac_hmac_err_o),
      // [0]: fatal_fault
      .alert_tx_o  ( alert_tx_o[0:0] ),
      .alert_rx_i  ( alert_rx_i[0:0] ),

      // Inter-module signals
      .idle_o(clkmgr_aon_idle[0]),
      .tl_i(hmac_tl_req),
      .tl_o(hmac_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .rst_ni
  );
  
  kmac #(
    .AlertAsyncOn(2'b11),
    .EnMasking(KmacEnMasking),
    .SwKeyMasked(KmacSwKeyMasked),
    .SecCmdDelay(SecKmacCmdDelay),
    .SecIdleAcceptSwMsg(SecKmacIdleAcceptSwMsg),
    .RndCnstLfsrSeed(RndCnstKmacLfsrSeed),
    .RndCnstLfsrPerm(RndCnstKmacLfsrPerm),
    .RndCnstLfsrFwdPerm(RndCnstKmacLfsrFwdPerm),
    .RndCnstMsgPerm(RndCnstKmacMsgPerm)
  ) u_kmac (

      // Interrupt
      .intr_kmac_done_o  (intr_kmac_kmac_done_o),
      .intr_fifo_empty_o (intr_kmac_fifo_empty_o),
      .intr_kmac_err_o   (intr_kmac_kmac_err_o),
      // [1]: recov_operation_err
      // [2]: fatal_fault_err
      .alert_tx_o  ( alert_tx_o[2:1] ),
      .alert_rx_i  ( alert_rx_i[2:1] ),

      // Inter-module signals
      .keymgr_key_i(keymgr_kmac_key),
      .app_i(kmac_app_req),
      .app_o(kmac_app_rsp),
      .entropy_o(edn0_edn_req_intr[3]),
      .entropy_i(edn0_edn_rsp_intr[3]),
      // .entropy_o(edn0_edn_req_rot),
      // .entropy_i(edn0_edn_rsp_rot),
      .idle_o(clkmgr_aon_idle[1]),
      // .idle_o(clkmgr_aon_idle_rot),
      .en_masking_o(kmac_en_masking),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .tl_i(kmac_tl_req),
      .tl_o(kmac_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .clk_edn_i,
      .rst_shadowed_ni,
      .rst_ni,
      .rst_edn_ni
  );
  
  keymgr #(
    .AlertAsyncOn(2'b11),
    .KmacEnMasking(KeymgrKmacEnMasking),
    .RndCnstLfsrSeed(RndCnstKeymgrLfsrSeed),
    .RndCnstLfsrPerm(RndCnstKeymgrLfsrPerm),
    .RndCnstRandPerm(RndCnstKeymgrRandPerm),
    .RndCnstRevisionSeed(RndCnstKeymgrRevisionSeed),
    .RndCnstCreatorIdentitySeed(RndCnstKeymgrCreatorIdentitySeed),
    .RndCnstOwnerIntIdentitySeed(RndCnstKeymgrOwnerIntIdentitySeed),
    .RndCnstOwnerIdentitySeed(RndCnstKeymgrOwnerIdentitySeed),
    .RndCnstSoftOutputSeed(RndCnstKeymgrSoftOutputSeed),
    .RndCnstHardOutputSeed(RndCnstKeymgrHardOutputSeed),
    .RndCnstAesSeed(RndCnstKeymgrAesSeed),
    .RndCnstKmacSeed(RndCnstKeymgrKmacSeed),
    .RndCnstOtbnSeed(RndCnstKeymgrOtbnSeed),
    .RndCnstCdi(RndCnstKeymgrCdi),
    .RndCnstNoneSeed(RndCnstKeymgrNoneSeed)
  ) u_keymgr (

      // Interrupt
      .intr_op_done_o (intr_keymgr_op_done_o),
      // [3]: recov_operation_err
      // [4]: fatal_fault_err
      .alert_tx_o  ( alert_tx_o[4:3] ),
      .alert_rx_i  ( alert_rx_i[4:3] ),

      // Inter-module signals
      .edn_o(edn0_edn_req_intr[0]),
      .edn_i(edn0_edn_rsp_intr[0]),
      .aes_key_o(keymgr_aes_key),
      .kmac_key_o(keymgr_kmac_key),
      .otbn_key_o(keymgr_otbn_key),
      .kmac_data_o(kmac_app_req[0]),
      .kmac_data_i(kmac_app_rsp[0]),
      .otp_key_i(otp_ctrl_otp_keymgr_key),
      .otp_device_id_i(keymgr_otp_device_id),
      .flash_i(flash_ctrl_keymgr),
      .lc_keymgr_en_i(lc_ctrl_lc_keymgr_en),
      .lc_keymgr_div_i(lc_ctrl_lc_keymgr_div),
      .rom_digest_i(rom_ctrl_keymgr_data),
      .kmac_en_masking_i(kmac_en_masking),
      .tl_i(keymgr_tl_req),
      .tl_o(keymgr_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .clk_edn_i,
      .rst_shadowed_ni,
      .rst_ni,
      .rst_edn_ni
  );

  rom_ctrl #(
    .AlertAsyncOn(1'b1),
    .BootRomInitFile(RomCtrlBootRomInitFile),
    .RndCnstScrNonce(RndCnstRomCtrlScrNonce),
    .RndCnstScrKey(RndCnstRomCtrlScrKey),
    .SecDisableScrambling(SecRomCtrlDisableScrambling)
  ) u_rom_ctrl (
      // [5]: fatal
      .alert_tx_o  ( alert_tx_o[5:5] ),
      .alert_rx_i  ( alert_rx_i[5:5] ),

      // Inter-module signals
      .rom_cfg_i(ast_rom_cfg),
      .pwrmgr_data_o(rom_ctrl_pwrmgr_data),
      .keymgr_data_o(rom_ctrl_keymgr_data),
      .kmac_data_o(kmac_app_req[1]),
      .kmac_data_i(kmac_app_rsp[1]),
      // .kmac_data_o(kmac_app_req_rom),
      // .kmac_data_i(kmac_app_rsp_rom),
      .regs_tl_i(rom_ctrl_regs_tl_req),
      .regs_tl_o(rom_ctrl_regs_tl_rsp),
      .rom_tl_i(rom_ctrl_rom_tl_req),
      .rom_tl_o(rom_ctrl_rom_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .rst_ni
  );

  edn #(
    .AlertAsyncOn(2'b11),
    .NumEndPoints(8)
  ) u_edn0 (

      // Interrupt
      .intr_edn_cmd_req_done_o (intr_edn0_edn_cmd_req_done_o),
      .intr_edn_fatal_err_o    (intr_edn0_edn_fatal_err_o),
      // [6]: recov_alert
      // [7]: fatal_alert
      .alert_tx_o  ( alert_tx_o[7:6] ),
      .alert_rx_i  ( alert_rx_i[7:6] ),

      // Inter-module signals
      .csrng_cmd_o(csrng_csrng_cmd_req[0]),
      .csrng_cmd_i(csrng_csrng_cmd_rsp[0]),
      .edn_i(edn0_edn_req_intr),
      .edn_o(edn0_edn_rsp_intr),
      .tl_i(edn0_tl_req),
      .tl_o(edn0_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .rst_ni
  );

  csrng #(
    .AlertAsyncOn(2'b11),
    .RndCnstCsKeymgrDivNonProduction(RndCnstCsrngCsKeymgrDivNonProduction),
    .RndCnstCsKeymgrDivProduction(RndCnstCsrngCsKeymgrDivProduction),
    .SBoxImpl(CsrngSBoxImpl),
    .NHwApps(2)
  ) u_csrng (

      // Interrupt
      .intr_cs_cmd_req_done_o (intr_csrng_cs_cmd_req_done_o),
      .intr_cs_entropy_req_o  (intr_csrng_cs_entropy_req_o),
      .intr_cs_hw_inst_exc_o  (intr_csrng_cs_hw_inst_exc_o),
      .intr_cs_fatal_err_o    (intr_csrng_cs_fatal_err_o),
      // [8]: recov_alert
      // [9]: fatal_alert
      .alert_tx_o  ( alert_tx_o[9:8] ),
      .alert_rx_i  ( alert_rx_i[9:8] ),

      // Inter-module signals
      .csrng_cmd_i(csrng_csrng_cmd_req),
      .csrng_cmd_o(csrng_csrng_cmd_rsp),
      .entropy_src_hw_if_o(csrng_entropy_src_hw_if_req),
      .entropy_src_hw_if_i(csrng_entropy_src_hw_if_rsp),
      .cs_aes_halt_i(csrng_cs_aes_halt_req),
      .cs_aes_halt_o(csrng_cs_aes_halt_rsp),
      .otp_en_csrng_sw_app_read_i(csrng_otp_en_csrng_sw_app_read),
      .lc_hw_debug_en_i(lc_ctrl_lc_hw_debug_en),
      .tl_i(csrng_tl_req),
      .tl_o(csrng_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .rst_ni
  );

  always_comb begin
    if (!rng_mode) begin  // puf in rng mode
      es_rng_rsp_i_puf.rng_valid = rng4bit_done;
      es_rng_rsp_i_puf.rng_b = rng4bit; 
    end else begin
      // puf in puf mode, rng from lfsr
      es_rng_rsp_i_puf = es_rng_rsp_i;
    end
  end

  entropy_src #(
    .AlertAsyncOn(2'b11),
    .EsFifoDepth(EntropySrcEsFifoDepth),
    .Stub(EntropySrcStub)
  ) u_entropy_src (

      // Interrupt
      .intr_es_entropy_valid_o      (intr_entropy_src_es_entropy_valid_o),
      .intr_es_health_test_failed_o (intr_entropy_src_es_health_test_failed_o),
      .intr_es_observe_fifo_ready_o (intr_entropy_src_es_observe_fifo_ready_o),
      .intr_es_fatal_err_o          (intr_entropy_src_es_fatal_err_o),
      // [10]: recov_alert
      // [11]: fatal_alert
      .alert_tx_o  ( alert_tx_o[11:10] ),
      .alert_rx_i  ( alert_rx_i[11:10] ),

      // Inter-module signals
      .entropy_src_hw_if_i(csrng_entropy_src_hw_if_req),
      .entropy_src_hw_if_o(csrng_entropy_src_hw_if_rsp),
      .cs_aes_halt_o(csrng_cs_aes_halt_req),
      .cs_aes_halt_i(csrng_cs_aes_halt_rsp),
      .entropy_src_rng_o(es_rng_req_o),
      .entropy_src_rng_i(es_rng_rsp_i_puf),
      .entropy_src_xht_o(),
      .entropy_src_xht_i(entropy_src_pkg::ENTROPY_SRC_XHT_RSP_DEFAULT),
      .otp_en_entropy_src_fw_read_i(entropy_src_otp_en_entropy_src_fw_read),
      .otp_en_entropy_src_fw_over_i(entropy_src_otp_en_entropy_src_fw_over),
      .rng_fips_o(es_rng_fips_o),
      .tl_i(entropy_src_tl_req),
      .tl_o(entropy_src_tl_rsp),

      // Clock and reset connections
      .clk_i,
      .rst_ni
  );

  otbn #(
    .AlertAsyncOn(2'b11),
    .Stub(OtbnStub),
    .RegFile(OtbnRegFile),
    .RndCnstUrndPrngSeed(RndCnstOtbnUrndPrngSeed),
    .SecMuteUrnd(SecOtbnMuteUrnd),
    .SecSkipUrndReseedAtStart(SecOtbnSkipUrndReseedAtStart),
    .RndCnstOtbnKey(RndCnstOtbnOtbnKey),
    .RndCnstOtbnNonce(RndCnstOtbnOtbnNonce)
  ) u_otbn (

      // Interrupt
      .intr_done_o (intr_otbn_done),
      // [12]: fatal
      // [13]: recov
      .alert_tx_o  ( alert_tx_o[13:12] ),
      .alert_rx_i  ( alert_rx_i[13:12] ),

      // Inter-module signals
      .otbn_otp_key_o(otp_ctrl_otbn_otp_key_req),
      .otbn_otp_key_i(otp_ctrl_otbn_otp_key_rsp),
      .edn_rnd_o(edn0_edn_req_intr[5]),
      .edn_rnd_i(edn0_edn_rsp_intr[5]),
      .edn_urnd_o(edn0_edn_req_intr[6]),
      .edn_urnd_i(edn0_edn_rsp_intr[6]),
      .idle_o(clkmgr_aon_idle[2]),
      .ram_cfg_i(ast_ram_1p_cfg),
      .lc_escalate_en_i(lc_ctrl_lc_escalate_en),
      .lc_rma_req_i(flash_ctrl_rma_ack),
      .lc_rma_ack_o(otbn_lc_rma_ack),
      .keymgr_key_i(keymgr_otbn_key),
      .tl_i(otbn_tl_req),
      .tl_o(otbn_tl_rsp),

      // Clock and reset connections
      .clk_i (clk_i),
      .clk_edn_i (clk_edn_i),
      .clk_otp_i (clk_i),
      .rst_ni (rst_ni),
      .rst_edn_ni (rst_edn_ni),
      .rst_otp_ni (rst_ni)
  );

  otbn_otp_controller u_otbn_otp_ctrl (
    .clk(clk_i),
    .rst_n(rst_ni),
    .req(otp_ctrl_otbn_otp_key_req),
    .rsp(otp_ctrl_otbn_otp_key_rsp)
  );

  sm3 u_sm3 (

      // Inter-module signals
      .tl_i(sm3_tl_req),
      .tl_o(sm3_tl_rsp),

      // Clock and reset connections
      .clk_i (clk_i),
      .rst_ni (rst_ni)
  );
  sm4 u_sm4 (

      // Inter-module signals
      .tl_i(sm4_tl_req),
      .tl_o(sm4_tl_rsp),

      // Clock and reset connections
      .clk_i (clk_i),
      .rst_ni (rst_ni)
  );

  rs_encode u_rs_encode (

      // Inter-module signals
      .tl_i(rs_encode_tl_req),
      .tl_o(rs_encode_tl_rsp),
      .scan_mode(scan_mode),

      // Clock and reset connections
      .clk_i (clk_i),
      .rst_ni (rst_ni)
  );
  rs_decode u_rs_decode (

      // Inter-module signals
      .tl_i(rs_decode_tl_req),
      .tl_o(rs_decode_tl_rsp),
      .scan_mode(scan_mode),

      // Clock and reset connections
      .clk_i (clk_i),
      .rst_ni (rst_ni)
  );
  puf u_puf (

      // Inter-module signals
      .tl_i(puf_tl_req),
      .tl_o(puf_tl_rsp),

      .rng4bit                 ( rng4bit ),
      .rng4bit_done            ( rng4bit_done ),
      .rng_mode                ( rng_mode ),
      .es_rng_req              ( es_rng_req_o ),

      // Clock and reset connections
      .clk_i (clk_i),
      .rst_ni (rst_ni)
  );

  puf u_puf2 (

      // Inter-module signals
      .tl_i(puf2_tl_req),
      .tl_o(puf2_tl_rsp),

      .rng4bit                 (  ),
      .rng4bit_done            (  ),
      .rng_mode                (  ),
      .es_rng_req              ( '0 ),

      // Clock and reset connections
      .clk_i (clk_i),
      .rst_ni (rst_ni)
  );

  xbar_main_rot u_xbar_main (
    .clk_i,
    .rst_ni,

    // port: tl_rv_core_ibex__corei
    .tl_host_i(tl_i),
    .tl_host_o(tl_o),

    // // port: tl_rom_ctrl__rom
    // .tl_rom_ctrl__rom_o(rom_ctrl_rom_tl_req),
    // .tl_rom_ctrl__rom_i(rom_ctrl_rom_tl_rsp),

    // port: tl_rom_ctrl__regs
    .tl_rom_ctrl__regs_o(rom_ctrl_regs_tl_req),
    .tl_rom_ctrl__regs_i(rom_ctrl_regs_tl_rsp),

    // port: tl_hmac
    .tl_hmac_o(hmac_tl_req),
    .tl_hmac_i(hmac_tl_rsp),

    // port: tl_kmac
    .tl_kmac_o(kmac_tl_req),
    .tl_kmac_i(kmac_tl_rsp),

    // port: tl_keymgr
    .tl_keymgr_o(keymgr_tl_req),
    .tl_keymgr_i(keymgr_tl_rsp),

    // port: tl_entropy_src
    .tl_entropy_src_o(entropy_src_tl_req),
    .tl_entropy_src_i(entropy_src_tl_rsp),

    // // port: tl_csrng
    .tl_csrng_o(csrng_tl_req),
    .tl_csrng_i(csrng_tl_rsp),

    // port: tl_edn0
    .tl_edn0_o(edn0_tl_req),
    .tl_edn0_i(edn0_tl_rsp),
    
    // port: tl_otbn
    .tl_otbn_o(otbn_tl_req),
    .tl_otbn_i(otbn_tl_rsp),

    // port: tl_sm3
    .tl_sm3_o(sm3_tl_req),
    .tl_sm3_i(sm3_tl_rsp),

    // port: tl_sm4
    .tl_sm4_o(sm4_tl_req),
    .tl_sm4_i(sm4_tl_rsp),

     // port: tl_rs_encode
    .tl_rs_encode_o(rs_encode_tl_req),
    .tl_rs_encode_i(rs_encode_tl_rsp),

    // port: tl_rs_decode
    .tl_rs_decode_o(rs_decode_tl_req),
    .tl_rs_decode_i(rs_decode_tl_rsp),

    // port: tl_puf
    .tl_puf_o(puf_tl_req),
    .tl_puf_i(puf_tl_rsp),

    // port: tl_puf2
    .tl_puf2_o(puf2_tl_req),
    .tl_puf2_i(puf2_tl_rsp)

  );
    

endmodule



module otbn_otp_controller (
  input  logic               clk,    // Clock input
  input  logic               rst_n,  // Active low reset
  input otp_ctrl_pkg::otbn_otp_key_req_t       req,
  output otp_ctrl_pkg::otbn_otp_key_rsp_t       rsp
);

// LFSR signals
//reg [127:0] lfsr_key;
//reg [63:0]  lfsr_nonce;

// Use a simple LFSR polynomial, e.g., x^128 + x^7 + x^2 + x + 1 for key
// and x^64 + x^4 + x^3 + x + 1 for nonce.
// These are not necessarily maximal length polynomials.
//wire lfsr_key_feedback = lfsr_key[127] ^ lfsr_key[7] ^ lfsr_key[2] ^ lfsr_key[1];
//wire lfsr_nonce_feedback = lfsr_nonce[63] ^ lfsr_nonce[4] ^ lfsr_nonce[3] ^ lfsr_nonce[1];

// Ack generation logic
reg ack_pulse;

// Generate a single-cycle pulse for ack
always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        ack_pulse      <= 1'b0;
  end else begin
        ack_pulse <= req.req && !ack_pulse; // Generate pulse on rising edge of req
  end
end

//assign rsp.key = lfsr_key;
//assign rsp.nonce = lfsr_nonce;

// LFSR and output logic
always_ff @(posedge clk or negedge rst_n) begin
  if (!rst_n) begin
    // Reset condition
    rsp.ack        <= 1'b0;
//    rsp.key        <= {128{1'b0}}; // Initialize with a non-zero random value
//    rsp.nonce      <= {64{1'b0}};  // Initialize with a non-zero random value
    rsp.seed_valid <= 1'b1;
    rsp.key       <= 128'h4235171482c225f79289b32181a0163a; // Initialize LFSR with a non-zero value
    rsp.nonce     <= 64'h760355d3447063d1;  // Initialize LFSR with a non-zero value
  //end else if (req.req)  begin
    // Update LFSRs with feedback
  //  lfsr_key   <= {lfsr_key[126:0], lfsr_key_feedback};
   // lfsr_nonce <= {lfsr_nonce[62:0], lfsr_nonce_feedback};
  end else if (ack_pulse) begin
      // Update key and nonce with new random values on ack pulse
    //lfsr_key   <= {lfsr_key[126:0], lfsr_key_feedback};
    //lfsr_nonce <= {lfsr_nonce[62:0], lfsr_nonce_feedback};
      rsp.key <= rsp.key + 1'b1;
      rsp.nonce <= rsp.nonce + 1'b1;
      rsp.ack <= ack_pulse;
  end else begin
    // Update the ack signal with the pulse
    rsp.ack <= ack_pulse;
  end
end

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// xbar_main module generated by `tlgen.py` tool
// all reset signals should be generated from one reset signal to not make any deadlock
//
// Interconnect

//   -> s1n_57
//     -> sm1_28
//       -> rom_ctrl.rom
//     -> sm1_33
//       -> rom_ctrl.regs
//     -> sm1_50
//       -> hmac
//     -> sm1_53
//       -> keymgr
//     -> sm1_54
//       -> kmac
//     -> sm1_46
//       -> entropy_src
//     -> sm1_47
//       -> csrng
//     -> sm1_48
//       -> edn0
//     -> sm1_52
//       -> otbn
//     -> sm1_60
//       -> sm3
//     -> sm1_61
//       -> sm4
//     -> sm1_65
//       -> rs_encode
//     -> sm1_66
//       -> rs_decode
//     -> sm1_67
//       -> puf
//     -> sm1_68
//       -> puf

module xbar_main_rot (
  input clk_i,
  input rst_ni,
  

  // Host interfaces
  input  tlul_pkg::tl_h2d_t tl_host_i,
  output tlul_pkg::tl_d2h_t tl_host_o,
  

  // Device interfaces
  // output tlul_pkg::tl_h2d_t tl_rom_ctrl__rom_o,
  // input  tlul_pkg::tl_d2h_t tl_rom_ctrl__rom_i,
  output tlul_pkg::tl_h2d_t tl_rom_ctrl__regs_o,
  input  tlul_pkg::tl_d2h_t tl_rom_ctrl__regs_i,
  output tlul_pkg::tl_h2d_t tl_hmac_o,
  input  tlul_pkg::tl_d2h_t tl_hmac_i,
  output tlul_pkg::tl_h2d_t tl_kmac_o,
  input  tlul_pkg::tl_d2h_t tl_kmac_i,
  output tlul_pkg::tl_h2d_t tl_keymgr_o,
  input  tlul_pkg::tl_d2h_t tl_keymgr_i,
  output tlul_pkg::tl_h2d_t tl_entropy_src_o,
  input  tlul_pkg::tl_d2h_t tl_entropy_src_i,
  output tlul_pkg::tl_h2d_t tl_csrng_o,
  input  tlul_pkg::tl_d2h_t tl_csrng_i,
  output tlul_pkg::tl_h2d_t tl_edn0_o,
  input  tlul_pkg::tl_d2h_t tl_edn0_i,
  output tlul_pkg::tl_h2d_t tl_otbn_o,
  input  tlul_pkg::tl_d2h_t tl_otbn_i,
  output tlul_pkg::tl_h2d_t tl_sm3_o,
  input  tlul_pkg::tl_d2h_t tl_sm3_i,
  output tlul_pkg::tl_h2d_t tl_sm4_o,
  input  tlul_pkg::tl_d2h_t tl_sm4_i,
  output tlul_pkg::tl_h2d_t tl_rs_encode_o,
  input  tlul_pkg::tl_d2h_t tl_rs_encode_i,
  output tlul_pkg::tl_h2d_t tl_rs_decode_o,
  input  tlul_pkg::tl_d2h_t tl_rs_decode_i,
  output tlul_pkg::tl_h2d_t tl_puf_o,
  input  tlul_pkg::tl_d2h_t tl_puf_i,
  output tlul_pkg::tl_h2d_t tl_puf2_o,
  input  tlul_pkg::tl_d2h_t tl_puf2_i
);

  import tlul_pkg::*;
  import tl_main_rot_pkg::*;

  // scanmode_i is currently not used, but provisioned for future use
  // this assignment prevents lint warnings
//   logic unused_scanmode;
//   assign unused_scanmode = ^scanmode_i;


  // Create steering signal


  // tl_h2d_t tl_sm1_28_us_h2d [1];
  // tl_d2h_t tl_sm1_28_us_d2h [1];

  // tl_h2d_t tl_sm1_28_ds_h2d ;
  // tl_d2h_t tl_sm1_28_ds_d2h ;


  tl_h2d_t tl_s1n_32_us_h2d ;
  tl_h2d_t tl_s1n_32_us_h2d_mask ;
  tl_d2h_t tl_s1n_32_us_d2h ;


  tl_h2d_t tl_s1n_32_ds_h2d [14];
  tl_d2h_t tl_s1n_32_ds_d2h [14];

  // Create steering signal
  logic [3:0] dev_sel_s1n_32;


  tl_h2d_t tl_sm1_33_us_h2d [1];
  tl_d2h_t tl_sm1_33_us_d2h [1];

  tl_h2d_t tl_sm1_33_ds_h2d ;
  tl_d2h_t tl_sm1_33_ds_d2h ;


  tl_h2d_t tl_sm1_50_us_h2d [1];
  tl_d2h_t tl_sm1_50_us_d2h [1];

  tl_h2d_t tl_sm1_50_ds_h2d ;
  tl_d2h_t tl_sm1_50_ds_d2h ;


  tl_h2d_t tl_sm1_53_us_h2d [1];
  tl_d2h_t tl_sm1_53_us_d2h [1];

  tl_h2d_t tl_sm1_53_ds_h2d ;
  tl_d2h_t tl_sm1_53_ds_d2h ;


  tl_h2d_t tl_sm1_54_us_h2d [1];
  tl_d2h_t tl_sm1_54_us_d2h [1];

  tl_h2d_t tl_sm1_54_ds_h2d ;
  tl_d2h_t tl_sm1_54_ds_d2h ;

  tl_h2d_t tl_sm1_46_us_h2d [1];
  tl_d2h_t tl_sm1_46_us_d2h [1];

  tl_h2d_t tl_sm1_46_ds_h2d ;
  tl_d2h_t tl_sm1_46_ds_d2h ;


  tl_h2d_t tl_sm1_47_us_h2d [1];
  tl_d2h_t tl_sm1_47_us_d2h [1];

  tl_h2d_t tl_sm1_47_ds_h2d ;
  tl_d2h_t tl_sm1_47_ds_d2h ;


  tl_h2d_t tl_sm1_48_us_h2d [1];
  tl_d2h_t tl_sm1_48_us_d2h [1];

  tl_h2d_t tl_sm1_48_ds_h2d ;
  tl_d2h_t tl_sm1_48_ds_d2h ;

  tl_h2d_t tl_sm1_52_us_h2d [1];
  tl_d2h_t tl_sm1_52_us_d2h [1];

  tl_h2d_t tl_sm1_52_ds_h2d ;
  tl_d2h_t tl_sm1_52_ds_d2h ;

  tl_h2d_t tl_sm1_60_us_h2d [1];
  tl_d2h_t tl_sm1_60_us_d2h [1];

  tl_h2d_t tl_sm1_60_ds_h2d ;
  tl_d2h_t tl_sm1_60_ds_d2h ;


  tl_h2d_t tl_sm1_61_us_h2d [1];
  tl_d2h_t tl_sm1_61_us_d2h [1];

  tl_h2d_t tl_sm1_61_ds_h2d ;
  tl_d2h_t tl_sm1_61_ds_d2h ;

  tl_h2d_t tl_sm1_65_us_h2d [1];
  tl_d2h_t tl_sm1_65_us_d2h [1];

  tl_h2d_t tl_sm1_65_ds_h2d ;
  tl_d2h_t tl_sm1_65_ds_d2h ;


  tl_h2d_t tl_sm1_66_us_h2d [1];
  tl_d2h_t tl_sm1_66_us_d2h [1];

  tl_h2d_t tl_sm1_66_ds_h2d ;
  tl_d2h_t tl_sm1_66_ds_d2h ;


  tl_h2d_t tl_sm1_67_us_h2d [1];
  tl_d2h_t tl_sm1_67_us_d2h [1];

  tl_h2d_t tl_sm1_67_ds_h2d ;
  tl_d2h_t tl_sm1_67_ds_d2h ;

  tl_h2d_t tl_sm1_68_us_h2d [1];
  tl_d2h_t tl_sm1_68_us_d2h [1];

  tl_h2d_t tl_sm1_68_ds_h2d ;
  tl_d2h_t tl_sm1_68_ds_d2h ;



  // Create steering signal
  
  // assign tl_sm1_28_us_h2d[0] = tl_s1n_32_ds_h2d[0];
  // assign tl_s1n_32_ds_d2h[0] = tl_sm1_28_us_d2h[0];

  assign tl_sm1_33_us_h2d[0] = tl_s1n_32_ds_h2d[1];
  assign tl_s1n_32_ds_d2h[1] = tl_sm1_33_us_d2h[0];

  assign tl_sm1_50_us_h2d[0] = tl_s1n_32_ds_h2d[2];
  assign tl_s1n_32_ds_d2h[2] = tl_sm1_50_us_d2h[0];

  assign tl_sm1_53_us_h2d[0] = tl_s1n_32_ds_h2d[3];
  assign tl_s1n_32_ds_d2h[3] = tl_sm1_53_us_d2h[0];

  assign tl_sm1_54_us_h2d[0] = tl_s1n_32_ds_h2d[4];
  assign tl_s1n_32_ds_d2h[4] = tl_sm1_54_us_d2h[0];

  assign tl_sm1_46_us_h2d[0] = tl_s1n_32_ds_h2d[5];
  assign tl_s1n_32_ds_d2h[5] = tl_sm1_46_us_d2h[0];

  assign tl_sm1_47_us_h2d[0] = tl_s1n_32_ds_h2d[6];
  assign tl_s1n_32_ds_d2h[6] = tl_sm1_47_us_d2h[0];

  assign tl_sm1_48_us_h2d[0] = tl_s1n_32_ds_h2d[7];
  assign tl_s1n_32_ds_d2h[7] = tl_sm1_48_us_d2h[0];

  assign tl_sm1_52_us_h2d[0] = tl_s1n_32_ds_h2d[8];
  assign tl_s1n_32_ds_d2h[8] = tl_sm1_52_us_d2h[0];

  assign tl_sm1_60_us_h2d[0] = tl_s1n_32_ds_h2d[9];
  assign tl_s1n_32_ds_d2h[9] = tl_sm1_60_us_d2h[0];

  assign tl_sm1_61_us_h2d[0] = tl_s1n_32_ds_h2d[10];
  assign tl_s1n_32_ds_d2h[10] = tl_sm1_61_us_d2h[0];

  assign tl_sm1_65_us_h2d[0] = tl_s1n_32_ds_h2d[11];
  assign tl_s1n_32_ds_d2h[11] = tl_sm1_65_us_d2h[0];

  assign tl_sm1_66_us_h2d[0] = tl_s1n_32_ds_h2d[12];
  assign tl_s1n_32_ds_d2h[12] = tl_sm1_66_us_d2h[0];

  assign tl_sm1_67_us_h2d[0] = tl_s1n_32_ds_h2d[0];
  assign tl_s1n_32_ds_d2h[0] = tl_sm1_67_us_d2h[0];

  assign tl_sm1_68_us_h2d[0] = tl_s1n_32_ds_h2d[13];
  assign tl_s1n_32_ds_d2h[13] = tl_sm1_68_us_d2h[0];


  assign tl_s1n_32_us_h2d = tl_host_i;
  assign tl_host_o = tl_s1n_32_us_d2h;


  // assign tl_rom_ctrl__rom_o = tl_sm1_28_ds_h2d;
  // assign tl_sm1_28_ds_d2h = tl_rom_ctrl__rom_i;

  assign tl_rom_ctrl__regs_o = tl_sm1_33_ds_h2d;
  assign tl_sm1_33_ds_d2h = tl_rom_ctrl__regs_i;

  assign tl_hmac_o = tl_sm1_50_ds_h2d;
  assign tl_sm1_50_ds_d2h = tl_hmac_i;

  assign tl_keymgr_o = tl_sm1_53_ds_h2d;
  assign tl_sm1_53_ds_d2h = tl_keymgr_i;

  assign tl_kmac_o = tl_sm1_54_ds_h2d;
  assign tl_sm1_54_ds_d2h = tl_kmac_i;

  assign tl_entropy_src_o = tl_sm1_46_ds_h2d;
  assign tl_sm1_46_ds_d2h = tl_entropy_src_i;

  assign tl_csrng_o = tl_sm1_47_ds_h2d;
  assign tl_sm1_47_ds_d2h = tl_csrng_i;

  assign tl_edn0_o = tl_sm1_48_ds_h2d;
  assign tl_sm1_48_ds_d2h = tl_edn0_i;

  assign tl_otbn_o = tl_sm1_52_ds_h2d;
  assign tl_sm1_52_ds_d2h = tl_otbn_i;

  assign tl_sm3_o = tl_sm1_60_ds_h2d;
  assign tl_sm1_60_ds_d2h = tl_sm3_i;

  assign tl_sm4_o = tl_sm1_61_ds_h2d;
  assign tl_sm1_61_ds_d2h = tl_sm4_i;

  assign tl_rs_encode_o = tl_sm1_65_ds_h2d;
  assign tl_sm1_65_ds_d2h = tl_rs_encode_i;

  assign tl_rs_decode_o = tl_sm1_66_ds_h2d;
  assign tl_sm1_66_ds_d2h = tl_rs_decode_i;

  assign tl_puf_o = tl_sm1_67_ds_h2d;
  assign tl_sm1_67_ds_d2h = tl_puf_i;

  assign tl_puf2_o = tl_sm1_68_ds_h2d;
  assign tl_sm1_68_ds_d2h = tl_puf2_i;

  

  always_comb begin
    // default steering to generate error response if address is not within the range
    dev_sel_s1n_32 = 4'd14;
    tl_s1n_32_us_h2d_mask = tl_s1n_32_us_h2d;
    // if ((tl_s1n_32_us_h2d.a_address &
    //      ~(ADDR_MASK_ROM_CTRL__ROM_ROT)) == ADDR_SPACE_ROM_CTRL__ROM_ROT) begin
    //   dev_sel_s1n_32 = 4'd0;
    //   tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_ROM_CTRL__ROM_ROT;

    // end else 
    if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_ROM_CTRL__REGS_ROT)) == ADDR_SPACE_ROM_CTRL__REGS_ROT) begin
      dev_sel_s1n_32 = 4'd1;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_ROM_CTRL__REGS_ROT;
    
    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_HMAC_ROT)) == ADDR_SPACE_HMAC_ROT) begin
      dev_sel_s1n_32 = 4'd2;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_HMAC_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_KEYMGR_ROT)) == ADDR_SPACE_KEYMGR_ROT) begin
      dev_sel_s1n_32 = 4'd3;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_KEYMGR_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_KMAC_ROT)) == ADDR_SPACE_KMAC_ROT) begin
      dev_sel_s1n_32 = 4'd4;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_KMAC_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_ENTROPY_SRC_ROT)) == ADDR_SPACE_ENTROPY_SRC_ROT) begin
      dev_sel_s1n_32 = 4'd5;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_ENTROPY_SRC_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_CSRNG_ROT)) == ADDR_SPACE_CSRNG_ROT) begin
      dev_sel_s1n_32 = 4'd6;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_CSRNG_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_EDN0_ROT)) == ADDR_SPACE_EDN0_ROT) begin
      dev_sel_s1n_32 = 4'd7;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_EDN0_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_OTBN_ROT)) == ADDR_SPACE_OTBN_ROT) begin
      dev_sel_s1n_32 = 4'd8;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_OTBN_ROT;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_SM3)) == ADDR_SPACE_SM3) begin
      dev_sel_s1n_32 = 5'd9;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_SM3;

    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_SM4)) == ADDR_SPACE_SM4) begin
      dev_sel_s1n_32 = 5'd10;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_SM4;
    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_RS_ENCODE)) == ADDR_SPACE_RS_ENCODE) begin
      dev_sel_s1n_32 = 5'd11;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_RS_ENCODE;
    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_RS_DECODE)) == ADDR_SPACE_RS_DECODE) begin
      dev_sel_s1n_32 = 5'd12;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_RS_DECODE;
    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_PUF)) == ADDR_SPACE_PUF) begin
      dev_sel_s1n_32 = 5'd0;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_PUF;
    end else if ((tl_s1n_32_us_h2d.a_address &
                  ~(ADDR_MASK_PUF2)) == ADDR_SPACE_PUF2) begin
      dev_sel_s1n_32 = 5'd13;
      tl_s1n_32_us_h2d_mask.a_address = tl_s1n_32_us_h2d.a_address & ADDR_MASK_PUF2;
    end
  end


  // Instantiation phase
 
  // tlul_socket_m1 #(
  //   .HReqDepth (12'h0),
  //   .HRspDepth (12'h0),
  //   .DRspPass  (1'b0),
  //   .M         (1)
  // ) u_sm1_28 (
  //   .clk_i        (clk_i),
  //   .rst_ni       (rst_ni),
  //   .tl_h_i       (tl_sm1_28_us_h2d),
  //   .tl_h_o       (tl_sm1_28_us_d2h),
  //   .tl_d_o       (tl_sm1_28_ds_h2d),
  //   .tl_d_i       (tl_sm1_28_ds_d2h)
  // );
  
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_33 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_33_us_h2d),
    .tl_h_o       (tl_sm1_33_us_d2h),
    .tl_d_o       (tl_sm1_33_ds_h2d),
    .tl_d_i       (tl_sm1_33_ds_d2h)
  );
  
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_50 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_50_us_h2d),
    .tl_h_o       (tl_sm1_50_us_d2h),
    .tl_d_o       (tl_sm1_50_ds_h2d),
    .tl_d_i       (tl_sm1_50_ds_d2h)
  );
  
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_53 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_53_us_h2d),
    .tl_h_o       (tl_sm1_53_us_d2h),
    .tl_d_o       (tl_sm1_53_ds_h2d),
    .tl_d_i       (tl_sm1_53_ds_d2h)
  );

  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_54 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_54_us_h2d),
    .tl_h_o       (tl_sm1_54_us_d2h),
    .tl_d_o       (tl_sm1_54_ds_h2d),
    .tl_d_i       (tl_sm1_54_ds_d2h)
  );
  
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_46 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_46_us_h2d),
    .tl_h_o       (tl_sm1_46_us_d2h),
    .tl_d_o       (tl_sm1_46_ds_h2d),
    .tl_d_i       (tl_sm1_46_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_47 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_47_us_h2d),
    .tl_h_o       (tl_sm1_47_us_d2h),
    .tl_d_o       (tl_sm1_47_ds_h2d),
    .tl_d_i       (tl_sm1_47_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_48 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_48_us_h2d),
    .tl_h_o       (tl_sm1_48_us_d2h),
    .tl_d_o       (tl_sm1_48_ds_h2d),
    .tl_d_i       (tl_sm1_48_ds_d2h)
  );

  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_52 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_52_us_h2d),
    .tl_h_o       (tl_sm1_52_us_d2h),
    .tl_d_o       (tl_sm1_52_ds_h2d),
    .tl_d_i       (tl_sm1_52_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_60 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_60_us_h2d),
    .tl_h_o       (tl_sm1_60_us_d2h),
    .tl_d_o       (tl_sm1_60_ds_h2d),
    .tl_d_i       (tl_sm1_60_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_61 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_61_us_h2d),
    .tl_h_o       (tl_sm1_61_us_d2h),
    .tl_d_o       (tl_sm1_61_ds_h2d),
    .tl_d_i       (tl_sm1_61_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_65 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_65_us_h2d),
    .tl_h_o       (tl_sm1_65_us_d2h),
    .tl_d_o       (tl_sm1_65_ds_h2d),
    .tl_d_i       (tl_sm1_65_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_66 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_66_us_h2d),
    .tl_h_o       (tl_sm1_66_us_d2h),
    .tl_d_o       (tl_sm1_66_ds_h2d),
    .tl_d_i       (tl_sm1_66_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_67 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_67_us_h2d),
    .tl_h_o       (tl_sm1_67_us_d2h),
    .tl_d_o       (tl_sm1_67_ds_h2d),
    .tl_d_i       (tl_sm1_67_ds_d2h)
  );
  tlul_socket_m1 #(
    .HReqDepth (8'h0),
    .HRspDepth (8'h0),
    .DReqPass  (1'b0),
    .DRspPass  (1'b0),
    .M         (1)
  ) u_sm1_68 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_sm1_68_us_h2d),
    .tl_h_o       (tl_sm1_68_us_d2h),
    .tl_d_o       (tl_sm1_68_ds_h2d),
    .tl_d_i       (tl_sm1_68_ds_d2h)
  );

  tlul_socket_1n #(
    .HReqDepth (4'h0),
    .HRspDepth (4'h0),
    .DReqDepth (56'h0),
    .DRspDepth (56'h0),
    .N         (14)
  ) u_s1n_32 (
    .clk_i        (clk_i),
    .rst_ni       (rst_ni),
    .tl_h_i       (tl_s1n_32_us_h2d_mask),
    .tl_h_o       (tl_s1n_32_us_d2h),
    .tl_d_o       (tl_s1n_32_ds_h2d),
    .tl_d_i       (tl_s1n_32_ds_d2h),
    .dev_select_i (dev_sel_s1n_32)
  );
 

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//############################################################################
// *Name: ast_pulse_symc
// *Module Description: AST Pulse Synchronizer
//
// Synchronizes a pulse from source clock domain (clk_src) to destination
// clock domain (clk_dst). The source pulse can have any length of the
// source clock cycle.
// The destination pulse has the length of one destination clock cycle.
// Consecutive pulses need to be spaced appropriately apart from each other
// depending on the clock frequency ratio of the two clock domains.
//############################################################################

`include "prim_assert.sv"

module ast_pulse_sync (
  input scan_mode_i,
  // source clock domain
  input clk_src_i,
  input rst_src_ni,
  input src_pulse_i,
  output logic src_pulse_en_o,
  output logic src_busy_o,
  // destination clock domain
  input clk_dst_i,
  input rst_dst_ni,
  output logic dst_pulse_o
);

// Reset all flops by both resets
////////////////////////////////////////
logic rst_src_n, rst_dst_da_n;
logic rst_dst_n, rst_src_da_n;

prim_flop_2sync #(
  .Width ( 1 ),
  .ResetValue ( 1'b0 )
) u_rst_dst_da (
  .clk_i ( clk_src_i),
  .rst_ni ( rst_dst_ni ),
  .d_i ( 1'b1 ),
  .q_o ( rst_dst_da_n )
);

prim_flop_2sync #(
  .Width ( 1 ),
  .ResetValue ( 1'b0 )
) u_rst_src_da (
  .clk_i ( clk_dst_i),
  .rst_ni ( rst_src_ni ),
  .d_i ( 1'b1 ),
  .q_o ( rst_src_da_n )
);

assign rst_src_n = scan_mode_i ? rst_src_ni : rst_src_ni && rst_dst_da_n;
assign rst_dst_n = scan_mode_i ? rst_dst_ni : rst_dst_ni && rst_src_da_n;


// Pulse Rising Edge Detect & Block
///////////////////////////////////////
logic src_pulse_d;

always_ff @( posedge clk_src_i, negedge rst_src_n ) begin
  if ( !rst_src_n ) begin
    src_pulse_d <= 1'b0;
  end else begin
    src_pulse_d <= src_pulse_i;
  end
end

assign src_pulse_en_o = src_pulse_i & !src_pulse_d & !src_busy_o;


// Pulse Transformation
///////////////////////////////////////
logic src_req;

// Convert src_pulse_en to a level signal
always_ff @( posedge clk_src_i, negedge rst_src_n ) begin
 if ( !rst_src_n ) begin
   src_req <= 1'b0;
  end else begin
   src_req <= (src_pulse_en_o ^ src_req);
  end
end


// SRC_REQ Synchronizer to DST
///////////////////////////////////////
logic dst_req;

prim_flop_2sync #(
  .Width ( 1 ),
  .ResetValue ( 1'b0 )
) u_dst_req (
  .clk_i ( clk_dst_i ),
  .rst_ni ( rst_dst_n ),
  .d_i ( src_req ),
  .q_o ( dst_req )
);


// DST_REQ Synchronizer to SRC for ACK
///////////////////////////////////////
logic src_ack;

prim_flop_2sync #(
  .Width ( 1 ),
  .ResetValue ( 1'b0 )
) u_sync2_ack (
  .clk_i ( clk_src_i ),
  .rst_ni ( rst_src_n ),
  .d_i ( dst_req ),
  .q_o ( src_ack )
);

// Source is BUSY when REQ not equel to ACK
assign src_busy_o = (src_req ^ src_ack);


// Pulse Reconstruction
///////////////////////////////////////
logic dst_req_d;

always_ff @( posedge clk_dst_i, negedge rst_dst_n ) begin
  if ( !rst_dst_n ) begin
    dst_req_d <= 1'b0;
  end else begin
    dst_req_d <= dst_req;
  end
end

assign dst_pulse_o = (dst_req ^ dst_req_d);


////////////////////
// Assertions
////////////////////

// A new PULSE can only be introduced when source is not BUSY.
`ASSERT(NewPulseWhenSrcBusy, $rose(src_pulse_i) |-> !src_busy_o, clk_src_i, !rst_src_n)

`ASSERT(DstPulseCheck_A, dst_pulse_o |=> !dst_pulse_o, clk_dst_i, !rst_dst_n)

endmodule : ast_pulse_sync


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// -------- W A R N I N G: A U T O - G E N E R A T E D  C O D E !! -------- //
// PLEASE DO NOT HAND-EDIT THIS FILE. IT HAS BEEN AUTO-GENERATED.
//
//############################################################################
// *Name: rng
// *Module Description:  Random (bit/s) Generator (Pseudo Model)
//############################################################################

`include "prim_assert.sv"

module rng #(
  parameter int EntropyStreams = 4
) (
  input clk_i,                                // Non-Jittery Clock (TLUL)
  input rst_ni,                               // Non-Jittery Reset (TLUL)
  input clk_ast_rng_i,                        // Jittery Clock (RNG)
  input rst_ast_rng_ni,                       // Jittery Reset (RNG)
  input rng_en_i,                             // RNG Enable
  input rng_fips_i,                           // RNG FIPS Enable
  input scan_mode_i,                          // Scan Mode
  output logic [EntropyStreams-1:0] rng_b_o,  // RNG Bus/Bits Output
  output logic rng_val_o                      // RNG Bus/Bits Valid
);

///////////////////////////////////////
// RNG Bus using LFSR
///////////////////////////////////////
logic rst_n;
logic[EntropyStreams-1:0] lfsr_val;

assign rst_n = scan_mode_i ? rst_ni : rst_ni && rng_en_i;

// These LFSR parameters have been generated with
// $ ./util/design/gen-lfsr-seed.py --width 64 --seed 15513 --prefix "Rng"
localparam int RngLfsrWidth = 64;
typedef logic [RngLfsrWidth-1:0] rng_lfsr_seed_t;
typedef logic [RngLfsrWidth-1:0][$clog2(RngLfsrWidth)-1:0] rng_lfsr_perm_t;
localparam rng_lfsr_seed_t RndCnstRngLfsrSeedDefault = 64'h1d033d20eed3b14;
localparam rng_lfsr_perm_t RndCnstRngLfsrPermDefault = {
  128'h98c2c94ab5e40420ed73f6c7396cd9e1,
  256'h58c6d7435ddb2ed1f22400c53a5aaa796ef7785e120628fbabc87f0b3928550f
};

prim_lfsr #(
  .LfsrDw ( RngLfsrWidth ),
  .EntropyDw ( 1 ),
  .StateOutDw ( EntropyStreams ),
  .DefaultSeed ( RndCnstRngLfsrSeedDefault ),
  .StatePermEn ( 1'b1 ),
  .StatePerm ( RndCnstRngLfsrPermDefault ),
  .ExtSeedSVA ( 1'b0 )  // ext seed is unused
) u_rng_lfsr (
  .clk_i ( clk_i ),
  .rst_ni ( rst_n ),
  .lfsr_en_i ( rng_en_i ),
  .seed_en_i ( 1'b0 ),
  .seed_i ( '0 ),
  .entropy_i ( 1'b0 ),
  .state_o ( lfsr_val )
);

logic srate_rng_val;
logic [12-1:0] srate_cnt, srate_value;
logic [EntropyStreams-1:0] rng_b;

`ifndef SYNTHESIS
logic [12-1:0] dv_srate_value;
// 4-bit rng_b needs at least 5 clocks. While the limit for these min and max values is 5:500, the
// default is set to a shorter window of 32:128 to avoid large runtimes.
logic [12-1:0] rng_srate_value_min = 12'd32;
logic [12-1:0] rng_srate_value_max = 12'd128;

initial begin : rng_plusargs
  void'($value$plusargs("rng_srate_value_min=%0d", rng_srate_value_min));
  void'($value$plusargs("rng_srate_value_max=%0d", rng_srate_value_max));
  `ASSERT_I(DvRngSrateMinCheck, rng_srate_value_min inside {[5:500]})
  `ASSERT_I(DvRngSrateMaxCheck, rng_srate_value_max inside {[5:500]})
  `ASSERT_I(DvRngSrateBoundsCheck, rng_srate_value_max >= rng_srate_value_min)
  dv_srate_value = 12'($urandom_range(int'(rng_srate_value_min), int'(rng_srate_value_max)));
  void'($value$plusargs("rng_srate_value=%0d", dv_srate_value));
  `ASSERT_I(DvSrateValueCheck, dv_srate_value inside {[5:500]})
end

assign srate_value = dv_srate_value;
`else
assign srate_value = 12'd120;
`endif

logic src_busy;

always_ff @( posedge clk_i, negedge rst_n ) begin
  if ( !rst_n ) begin
    srate_cnt     <= 12'h000;
    srate_rng_val <= 1'b0;
  end else if ( (srate_cnt == srate_value) && src_busy ) begin
    srate_rng_val <= 1'b0;
  end else if ( srate_cnt == srate_value ) begin
    srate_cnt     <= 12'h000;
    srate_rng_val <= 1'b1;
  end else begin
    srate_cnt     <= srate_cnt + 1'b1;
    srate_rng_val <= 1'b0;
  end
end


////////////////////////////////////////
// Sychronize Bus & Valid to RNG Clock
////////////////////////////////////////
logic sync_rng_val, srate_rng_val_en;

ast_pulse_sync u_rng_val_pulse_sync (
  .scan_mode_i ( scan_mode_i ),
  // source clock domain
  .clk_src_i ( clk_i ),
  .rst_src_ni ( rst_n ),
  .src_pulse_i ( srate_rng_val ),
  .src_pulse_en_o ( srate_rng_val_en ),
  .src_busy_o ( src_busy ),
  // destination clock domain
  .clk_dst_i ( clk_ast_rng_i ),
  .rst_dst_ni ( rst_ast_rng_ni ),
  .dst_pulse_o ( sync_rng_val )
);

// Sanple & Hold the rng_b value until the sync completes
always_ff @( posedge clk_i, negedge rst_n ) begin
  if ( !rst_n ) begin
    rng_b <= {EntropyStreams{1'b0}};
  end else if ( srate_rng_val_en ) begin
    rng_b <= lfsr_val[EntropyStreams-1:0];
  end
end

//Sync to RNG clock domain
always_ff @( posedge clk_ast_rng_i, negedge rst_ast_rng_ni ) begin
  if (!rst_ast_rng_ni ) begin
    rng_b_o <= {EntropyStreams{1'b0}};
    rng_val_o <= 1'b0;
  end else if ( sync_rng_val ) begin
    rng_b_o <= rng_b[EntropyStreams-1:0];
    rng_val_o <= 1'b1;
  end else begin
    rng_val_o <= 1'b0;
  end
end


///////////////////////
// Unused Signals
///////////////////////
logic unused_sigs;
assign unused_sigs = ^{
                        rng_fips_i  // Used in ASIC implementation
                      };

endmodule : rng


// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:     SHU
// Engineer:    lf
// 
// Create Date: 2020/04/26 16:24:02
// Design Name: 
// Module Name: adder_32b
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//              32 位 加法器 性能分析用
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_32b(
    input   [31:0]      A,
    input   [31:0]      B,
    output  [31:0]      R   
    );
    wire    [32:0]      R_tmp;         
    assign      R_tmp   = A + B;
    assign      R       = R_tmp[31:0];
endmodule


// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:     SHU
// Engineer:    lf
// 
// Create Date: 2020/04/26 16:24:02
// Design Name: 
// Module Name: csa_adder_3i_32b
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//              32 位 3 输入 CSA 加法器，不考虑进位 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module csa_adder_3i_32b(
    input   [31:0]      A,
    input   [31:0]      B,
    input   [31:0]      C,
    output  [31:0]      R   
    );

    wire [31:0]     S;
    wire [31:0]     Ca;
    wire [33:0]     R_tmp;

    //3-2 CSA
    assign  S = A ^ B ^ C;
    assign  Ca = (A & B) | (A & C) | (B & C);
    
    //加法器
    assign  R_tmp = {Ca,{1'b0}} + S;

    //输出端口,取低位，不考虑进位
    assign  R = R_tmp[31:0];
endmodule


// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Company:     SHU
// Engineer:    lf
// 
// Create Date: 2020/04/26 16:24:02
// Design Name: 
// Module Name: sm3_adder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//              SM3 32 位 3 输入 加法器，
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sm3_adder(
    input   [31:0]      A,
    input   [31:0]      B,
    input   [31:0]      C,
    output  [31:0]      R   
    );

    `ifdef SM3_CMPRSS_CSA_ADD
        //使用CSA加法器
        csa_adder_3i_32b U_csa_adder_3i_32b(
            .A(A),
            .B(B),
            .C(C),
            .R(R)  
        );
    `else
        //使用两级加法器
        wire [31:0]     tmp;
        adder_32b U_adder_0(
            .A(A),
            .B(B),
            .R(tmp) 
        );
        adder_32b U_adder_1(
            .A(tmp),
            .B(C),
            .R(R) 
        );

    `endif
    
endmodule


// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/28
// Design Name: sm3
// Module Name: sm3_cmprss_ceil_comb
// Description:
//      SM3 单轮迭代压缩模块 由组合逻辑构成
//      
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_cmprss_ceil_comb(
    input                   cmprss_round_sm_16_i,
    input [31:0]            tj_i,

    input [31:0]            reg_a_i,
    input [31:0]            reg_b_i,
    input [31:0]            reg_c_i,
    input [31:0]            reg_d_i,
    input [31:0]            reg_e_i,
    input [31:0]            reg_f_i,
    input [31:0]            reg_g_i,
    input [31:0]            reg_h_i,

    input [31:0]            wj_i,
    input [31:0]            wjj_i,

    output [31:0]           reg_a_o,
    output [31:0]           reg_b_o,
    output [31:0]           reg_c_o,
    output [31:0]           reg_d_o,
    output [31:0]           reg_e_o,
    output [31:0]           reg_f_o,
    output [31:0]           reg_g_o,
    output [31:0]           reg_h_o
    );


//wire
wire [31:0]	tmp_for_ss1_0	;
wire [31:0]	tmp_for_ss1_2	;
wire [31:0]	ss1				;
wire [31:0]	ss2				;
wire [31:0]	tmp_for_tt1_0	;
wire [31:0]	tmp_for_tt1_1	;
wire [31:0]	tt1				;
wire [31:0]	tmp_for_tt2_0	;
wire [31:0]	tmp_for_tt2_1	;
wire [31:0]	tt2				;
wire [31:0]	tt2_after_p0	;

wire [31:0]	TJ				=	tj_i;

//加法器0
`ifdef SM3_CMPRSS_DIRECT_ADD
    assign  tmp_for_ss1_0	=	{reg_a_i[31-12:0], reg_a_i[31:31-12+1]} + reg_e_i;
    assign  tmp_for_ss1_2	=	tmp_for_ss1_0 + TJ;
`else
    sm3_adder U_ss1(
        .A({reg_a_i[31-12:0], reg_a_i[31:31-12+1]}),
        .B(reg_e_i),
        .C(TJ),
        .R(tmp_for_ss1_2) 
    );
`endif

assign      ss1				=	{tmp_for_ss1_2[31 - 7 : 0], tmp_for_ss1_2[31 : 31 - 7 + 1]};
assign  	ss2				=	ss1 ^ {reg_a_i[31 - 12 : 0], reg_a_i[31 : 31 - 12 + 1]};

//加法器1
assign  	tmp_for_tt1_0	=	cmprss_round_sm_16_i? reg_a_i ^ reg_b_i ^ reg_c_i : (reg_a_i & reg_b_i | reg_a_i & reg_c_i | reg_b_i & reg_c_i);
`ifdef SM3_CMPRSS_DIRECT_ADD
    assign  	tmp_for_tt1_1	=	reg_d_i + ss2 + wjj_i;
    assign  	tt1				=	tmp_for_tt1_0 + tmp_for_tt1_1;
`else
    //tmp_for_tt1_1 = reg_d_i + tmp_for_tt1_0 + wjj_i
    sm3_adder U_tmp_for_tt1_1(
        .A(reg_d_i),
        .B(tmp_for_tt1_0),
        .C(wjj_i),
        .R(tmp_for_tt1_1) 
    );
    //tt1 = ss2 + tmp_for_tt1_1
    adder_32b U_tt1(
        .A(ss2),
        .B(tmp_for_tt1_1),
        .R(tt1) 
    );
`endif

//加法器2
assign  	tmp_for_tt2_0	=	cmprss_round_sm_16_i? reg_e_i ^ reg_f_i ^ reg_g_i : (reg_e_i & reg_f_i | ~reg_e_i & reg_g_i);
`ifdef SM3_CMPRSS_DIRECT_ADD
    assign  	tmp_for_tt2_1	=	reg_h_i + ss1 + wj_i;
    assign  	tt2				=	tmp_for_tt2_0 + tmp_for_tt2_1;
`else
    //tmp_for_tt2_1 = reg_h_i + tmp_for_tt2_0 + wj_i
    sm3_adder U_tmp_for_tt2_1(
        .A(reg_h_i),
        .B(tmp_for_tt2_0),
        .C(wj_i),
        .R(tmp_for_tt2_1) 
    );
    //tt2 = ss1 + tmp_for_tt2_1
    adder_32b U_tt2(
        .A(ss1),
        .B(tmp_for_tt2_1),
        .R(tt2) 
    );
`endif

assign  	tt2_after_p0	=	tt2 ^ {tt2[31-9:0], tt2[31:31-9+1]} ^ {tt2[31-17:0], tt2[31:31-17+1]};

assign  reg_a_o             =   tt1;
assign  reg_b_o             =   reg_a_i;
assign  reg_c_o             =   {reg_b_i[31 - 9 : 0], reg_b_i[31 : 31 - 9 + 1]};
assign  reg_d_o             =   reg_c_i;
assign  reg_e_o             =   tt2_after_p0;
assign  reg_f_o             =   reg_e_i;
assign  reg_g_o             =   {reg_f_i[31 - 19 : 0], reg_f_i[31 : 31 - 19 + 1]};
assign  reg_h_o             =   reg_g_i;

endmodule


// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/27 
// Design Name: sm3
// Module Name: sm3_cmprss_core
// Description:
//      SM3 迭代压缩模块-SM3 迭代压缩核心单元
//      输入位宽：INPT_DW1 定义，支持32/64bit
//      输出位宽：与输入位宽对应
//      特性：在 64bit 位宽下，采用二度展开结构（暂未）
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_cmprss_core (
    input                       clk,
    input                       rst_n,

    input  [`INPT_DW1:0]        expnd_inpt_wj_i,                    
    input  [`INPT_DW1:0]        expnd_inpt_wjj_i,                    
    input                       expnd_inpt_lst_i,                  
    input                       expnd_inpt_vld_i,    

    output [255:0]              cmprss_otpt_res_o,
    output                      cmprss_otpt_vld_o
);

//每时钟输入的数据字数量 32bit位宽：1 64bit位宽：2
`ifdef SM3_INPT_DW_32
    localparam [1:0]            INPT_WORD_NUM               =   2'd1;
`elsif SM3_INPT_DW_64
    localparam [1:0]            INPT_WORD_NUM               =   2'd2;
`endif

localparam  [6:0]           CMPRSS_RND_NUM = 7'd64;

//A-H 字寄存器
reg		[31 : 0]	reg_a;
reg		[31 : 0]	reg_b;
reg		[31 : 0]	reg_c;
reg		[31 : 0]	reg_d;
reg		[31 : 0]	reg_e;
reg		[31 : 0]	reg_f;
reg		[31 : 0]	reg_g;
reg		[31 : 0]	reg_h;
reg		[31 : 0]	reg_tj;
reg		[5  : 0]	reg_cmprss_round;

reg                 cmprss_round_sm_16;

//结果寄存器
reg                 sm3_res_valid;
reg                 sm3_res_valid_r1;
reg  [255:0]        sm3_res;

reg                 cmprss_blk_res_finish;

//A-H 字运算中间值
wire	[31 : 0]	reg_a_new;
wire	[31 : 0]	reg_b_new;
wire	[31 : 0]	reg_c_new;
wire	[31 : 0]	reg_d_new;
wire	[31 : 0]	reg_e_new;
wire	[31 : 0]	reg_f_new;
wire	[31 : 0]	reg_g_new;
wire	[31 : 0]	reg_h_new;

`ifdef SM3_INPT_DW_64
    wire	[31 : 0]	reg_a_mid;
    wire	[31 : 0]	reg_b_mid;
    wire	[31 : 0]	reg_c_mid;
    wire	[31 : 0]	reg_d_mid;
    wire	[31 : 0]	reg_e_mid;
    wire	[31 : 0]	reg_f_mid;
    wire	[31 : 0]	reg_g_mid;
    wire	[31 : 0]	reg_h_mid;

    //两轮运算的 tj 值
    wire	[31 : 0]	reg_tj_rnd_odd;
    wire	[31 : 0]	reg_tj_rnd_even;
`endif

//块迭代标志
wire                cmprss_new_round_valid;
wire                cmprss_blk_start;  
wire                cmprss_blk_finish; 

//对输入的 wj 值打拍或者分离
reg                 sm3_wj_wjj_vld_r;
reg                 sm3_wj_wjj_lst_r;

`ifdef SM3_INPT_DW_32
    reg     [31:0]      wj_rnd_r;
    reg     [31:0]      wjj_rnd_r;
`elsif SM3_INPT_DW_64
    reg     [31:0]      wj_rnd_odd_r;
    reg     [31:0]      wjj_rnd_odd_r;
    reg     [31:0]      wj_rnd_even_r;
    reg     [31:0]      wjj_rnd_even_r;
`endif

//输入每数据块所属数据字计数
reg     [5:0]       inpt_wrd_of_blk_cntr;
wire                inpt_wrd_of_blk_cntr_add;
wire                inpt_wrd_of_blk_cntr_clr;

//管理tj寄存器
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        reg_tj          <=  32'h79cc4519;
    end else if (cmprss_blk_res_finish) begin
        reg_tj          <=  32'h79cc4519;
    end
    else if(sm3_wj_wjj_vld_r)begin
        if(reg_cmprss_round == 6'd16 - INPT_WORD_NUM)
            reg_tj          <=  32'h9d8a7a87;
        
        else begin
            `ifdef SM3_INPT_DW_32
                reg_tj          <=  {reg_tj[30:0],reg_tj[31]};
            `elsif SM3_INPT_DW_64 //每次循环左移两位
                reg_tj          <=  {reg_tj[29:0],reg_tj[31:30]};
            `endif
        end
    end
end

`ifdef SM3_INPT_DW_64
    //两轮运算的 tj 值
    assign  	reg_tj_rnd_odd      =   {reg_tj[30:0],reg_tj[31]};
    assign  	reg_tj_rnd_even     =   reg_tj;
`endif

//对输入的 wj 值打拍或者分离
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        sm3_wj_wjj_vld_r    <=   1'b0;
        sm3_wj_wjj_lst_r    <=   1'b0;        
    end
    else begin
        sm3_wj_wjj_vld_r    <=   expnd_inpt_vld_i;
        sm3_wj_wjj_lst_r    <=   expnd_inpt_lst_i;       
    end
end

`ifdef SM3_INPT_DW_32
    always @(posedge clk or negedge rst_n) begin
        if(~rst_n) begin
            wj_rnd_r        <=   32'd0;
            wjj_rnd_r       <=   32'd0;       
        end
        else begin
            wj_rnd_r        <=   expnd_inpt_wj_i;
            wjj_rnd_r       <=   expnd_inpt_wjj_i;     
        end
    end
    
`elsif SM3_INPT_DW_64
    always @(posedge clk or negedge rst_n) begin
        if(~rst_n) begin
            wj_rnd_odd_r    <=   32'd0;
            wjj_rnd_odd_r   <=   32'd0;       
            wj_rnd_even_r   <=   32'd0;       
            wjj_rnd_even_r  <=   32'd0;       
        end
        else begin
            {wj_rnd_even_r,wj_rnd_odd_r}    <=   expnd_inpt_wj_i;
            {wjj_rnd_even_r,wjj_rnd_odd_r}  <=   expnd_inpt_wjj_i;    
        end
    end
    
`endif

//标记最后一块
assign              cmprss_new_round_valid  =   sm3_wj_wjj_vld_r;  
assign              cmprss_blk_finish       =   inpt_wrd_of_blk_cntr_clr;  

//块运算完成信号 
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        cmprss_blk_res_finish   <=  1'b0;
    end
    else begin
        cmprss_blk_res_finish   <=  inpt_wrd_of_blk_cntr_clr;
    end
end

//输入每数据块所属数据字计数
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        inpt_wrd_of_blk_cntr              <= 6'b0;
    end else if(inpt_wrd_of_blk_cntr_add)begin
        inpt_wrd_of_blk_cntr              <= inpt_wrd_of_blk_cntr + INPT_WORD_NUM;
    end else if(inpt_wrd_of_blk_cntr_clr)begin
        inpt_wrd_of_blk_cntr              <= 6'b0;
    end
end
assign                  inpt_wrd_of_blk_cntr_add  = sm3_wj_wjj_vld_r;
assign                  inpt_wrd_of_blk_cntr_clr  = sm3_wj_wjj_vld_r 
                                                && inpt_wrd_of_blk_cntr == (CMPRSS_RND_NUM - INPT_WORD_NUM);

//压缩迭代轮计数
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        reg_cmprss_round        <=  6'd0;
    end
    else if(cmprss_blk_finish)begin
        reg_cmprss_round        <=  6'd0;
    end
    else if(cmprss_new_round_valid)begin
        reg_cmprss_round        <=  reg_cmprss_round + INPT_WORD_NUM;
    end
end

//产生16轮内标记
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        cmprss_round_sm_16      <= 1'b0;
    end else begin
        cmprss_round_sm_16      <= reg_cmprss_round <  6'd16 - INPT_WORD_NUM; //标识当前小于
    end
end

//寄存器组初值装填与迭代
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        reg_a	<=	32'h7380166f;//0;
		reg_b	<=	32'h4914b2b9;//0;
		reg_c	<=	32'h172442d7;//0;
		reg_d	<=	32'hda8a0600;//0;
		reg_e	<=	32'ha96f30bc;//0;
		reg_f	<=	32'h163138aa;//0;
		reg_g	<=	32'he38dee4d;//0;
		reg_h	<=	32'hb0fb0e4e;//0;
    end else if (sm3_res_valid_r1) begin
        reg_a	<=	32'h7380166f;//0;
		reg_b	<=	32'h4914b2b9;//0;
		reg_c	<=	32'h172442d7;//0;
		reg_d	<=	32'hda8a0600;//0;
		reg_e	<=	32'ha96f30bc;//0;
		reg_f	<=	32'h163138aa;//0;
		reg_g	<=	32'he38dee4d;//0;
		reg_h	<=	32'hb0fb0e4e;//0;
    end
    else if(cmprss_new_round_valid)begin
        reg_a	<=	reg_a_new;
		reg_b	<=	reg_b_new;
		reg_c	<=	reg_c_new;
		reg_d	<=	reg_d_new;
		reg_e	<=	reg_e_new;
		reg_f	<=	reg_f_new;
		reg_g	<=	reg_g_new;
		reg_h	<=	reg_h_new;
    end
    else if(cmprss_blk_res_finish)begin
        reg_a	<=	reg_a ^ sm3_res[255-:32];
		reg_b	<=	reg_b ^ sm3_res[223-:32];
		reg_c	<=	reg_c ^ sm3_res[191-:32];
		reg_d	<=	reg_d ^ sm3_res[159-:32];
		reg_e	<=	reg_e ^ sm3_res[127-:32];
		reg_f	<=	reg_f ^ sm3_res[95 -:32];
		reg_g	<=	reg_g ^ sm3_res[63 -:32];
		reg_h	<=	reg_h ^ sm3_res[31 -:32];
    end
end

//消息所属块均计算完毕，输出计算结果
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        sm3_res_valid           <=  1'b0;
        sm3_res_valid_r1        <=  1'b0;
    end
    else begin
        sm3_res_valid           <=  sm3_wj_wjj_lst_r;
        sm3_res_valid_r1        <=  sm3_res_valid;
    end
end

always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        sm3_res                 <=  {32'h7380166f, 32'h4914b2b9, 32'h172442d7, 32'hda8a0600, 32'ha96f30bc, 32'h163138aa, 32'he38dee4d, 32'hb0fb0e4e};
    end else if (sm3_res_valid_r1) begin
        sm3_res                 <=  {32'h7380166f, 32'h4914b2b9, 32'h172442d7, 32'hda8a0600, 32'ha96f30bc, 32'h163138aa, 32'he38dee4d, 32'hb0fb0e4e};        
    end
    else if(cmprss_blk_res_finish)begin
        sm3_res                 <=  {reg_a,reg_b,reg_c,reg_d,reg_e,reg_f,reg_g,reg_h} ^ sm3_res;
    end
end

`ifdef SM3_INPT_DW_32
    sm3_cmprss_ceil_comb U_sm3_cmprss_ceil_comb
    (
        .cmprss_round_sm_16_i   (cmprss_round_sm_16),
        .tj_i                   (reg_tj),
        .reg_a_i                (reg_a),
        .reg_b_i                (reg_b),
        .reg_c_i                (reg_c),
        .reg_d_i                (reg_d),
        .reg_e_i                (reg_e),
        .reg_f_i                (reg_f),
        .reg_g_i                (reg_g),
        .reg_h_i                (reg_h),
        .wj_i                   (wj_rnd_r),
        .wjj_i                  (wjj_rnd_r),
        .reg_a_o                (reg_a_new),
        .reg_b_o                (reg_b_new),
        .reg_c_o                (reg_c_new),
        .reg_d_o                (reg_d_new),
        .reg_e_o                (reg_e_new),
        .reg_f_o                (reg_f_new),
        .reg_g_o                (reg_g_new),
        .reg_h_o                (reg_h_new)
    );

`elsif SM3_INPT_DW_64
    sm3_cmprss_ceil_comb U_sm3_cmprss_ceil_comb
    (
        .cmprss_round_sm_16_i   (cmprss_round_sm_16),
        .tj_i                   (reg_tj_rnd_even),
        .reg_a_i                (reg_a),
        .reg_b_i                (reg_b),
        .reg_c_i                (reg_c),
        .reg_d_i                (reg_d),
        .reg_e_i                (reg_e),
        .reg_f_i                (reg_f),
        .reg_g_i                (reg_g),
        .reg_h_i                (reg_h),
        .wj_i                   (wj_rnd_even_r),
        .wjj_i                  (wjj_rnd_even_r),
        .reg_a_o                (reg_a_mid),
        .reg_b_o                (reg_b_mid),
        .reg_c_o                (reg_c_mid),
        .reg_d_o                (reg_d_mid),
        .reg_e_o                (reg_e_mid),
        .reg_f_o                (reg_f_mid),
        .reg_g_o                (reg_g_mid),
        .reg_h_o                (reg_h_mid)
    );

    sm3_cmprss_ceil_comb U_sm3_cmprss_ceil_comb_1
    (
        .cmprss_round_sm_16_i   (cmprss_round_sm_16),
        .tj_i                   (reg_tj_rnd_odd),
        .reg_a_i                (reg_a_mid),
        .reg_b_i                (reg_b_mid),
        .reg_c_i                (reg_c_mid),
        .reg_d_i                (reg_d_mid),
        .reg_e_i                (reg_e_mid),
        .reg_f_i                (reg_f_mid),
        .reg_g_i                (reg_g_mid),
        .reg_h_i                (reg_h_mid),
        .wj_i                   (wj_rnd_odd_r),
        .wjj_i                  (wjj_rnd_odd_r),
        .reg_a_o                (reg_a_new),
        .reg_b_o                (reg_b_new),
        .reg_c_o                (reg_c_new),
        .reg_d_o                (reg_d_new),
        .reg_e_o                (reg_e_new),
        .reg_f_o                (reg_f_new),
        .reg_g_o                (reg_g_new),
        .reg_h_o                (reg_h_new)
    );
`endif

//输出控制
assign                      cmprss_otpt_vld_o     =   sm3_res_valid_r1;
assign                      cmprss_otpt_res_o     =   sm3_res;

`ifdef SM3_CMPRS_SIM_DBG
    `ifdef SM3_CMPRS_SIM_FILE_LOG
        integer file;
        initial begin:inital_file
            
            file = $fopen("wj.txt","w");
        end
    `endif

    generate
        if(1) begin
            always@(*) begin		
                if(cmprss_otpt_vld_o)
                begin
                    `ifdef SM3_CMPRS_SIM_FILE_LOG
                        $fdisplay(file,"LOG: res : %64h",cmprss_otpt_res_o);
                    `else
                        $display("LOG: res : %64h",cmprss_otpt_res_o);
                    `endif
                    
                end
            end
        end
    endgenerate
`endif

endmodule

// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/26 
// Design Name: sm3
// Module Name: sm3_cmprss_core_wrapper
// Description:
//      sm3_cmprss_core 的 SV 封装
//          封装 sm3_if 总线接口，类型为 CMPRSS
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_cmprss_core_wrapper (
    sm3_if.CMPRSS sm3if
);

sm3_cmprss_core U_sm3_cmprss_core(
    .clk                        (sm3if.clk                    ),
    .rst_n                      (sm3if.rst_n                  ),

    .expnd_inpt_wj_i            ( sm3if.expnd_otpt_wj                  ),
    .expnd_inpt_wjj_i           ( sm3if.expnd_otpt_wjj                  ),
    .expnd_inpt_lst_i           ( sm3if.expnd_otpt_lst                  ),
    .expnd_inpt_vld_i           ( sm3if.expnd_otpt_vld                  ),

    .cmprss_otpt_res_o          ( sm3if.cmprss_otpt_res               ),
    .cmprss_otpt_vld_o          ( sm3if.cmprss_otpt_vld               )
);   
    
endmodule

// `timescale 1ns / 1ps
// `include "./inc/sm3_cfg.v"
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/29 
// Design Name: sm3
// Module Name: sm3_core_top
// Description:
//      SM3 顶层模块，例化下层的 SM3 填充、扩展以及迭代压缩三个模块
//      输入位宽：INPT_DW1 定义，支持32/64
//      输出位宽：与输入位宽一致
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_core_top (

    input                       clk,
    input                       rst_n,
    input [`INPT_DW1:0]         msg_inpt_d,
    input [`INPT_BYTE_DW1:0]    msg_inpt_vld_byte,
    input                       msg_inpt_vld,
    input                       msg_inpt_lst,
    
    output                      msg_inpt_rdy,

    output[255:0]               cmprss_otpt_res,
    output                      cmprss_otpt_vld,
    output                      msg_inpt_rdy_re,
    output                      cmprss_vld_re,
    output[7:0]                 cmprss_res_re
);

//interface
sm3_if int_if();
wire msg_inpt_lst_real;

assign msg_inpt_lst_real = msg_inpt_lst & msg_inpt_vld;
assign msg_inpt_rdy_re = 1'b1;
assign cmprss_vld_re = cmprss_otpt_vld;
assign cmprss_res_re = {8{cmprss_otpt_vld}};

sm3_pad_core U_sm3_pad_core(

    .clk                    (clk                    ),
    .rst_n                  (rst_n                  ),

    .msg_inpt_d_i           (msg_inpt_d             ),
    .msg_inpt_vld_byte_i    (msg_inpt_vld_byte      ),
    .msg_inpt_vld_i         (msg_inpt_vld           ),
    .msg_inpt_lst_i         (msg_inpt_lst_real      ),

    .msg_inpt_rdy_o         (msg_inpt_rdy           ),

    .pad_otpt_ena_i         (int_if.pad_otpt_ena        ),

    .pad_otpt_d_o           (int_if.pad_otpt_d             ),
    .pad_otpt_lst_o         (int_if.pad_otpt_lst           ),
    .pad_otpt_vld_o         (int_if.pad_otpt_vld           )
); 

sm3_expnd_core U_sm3_expnd_core(
    
    .clk                    (clk                    ),
    .rst_n                  (rst_n                  ),


    .pad_inpt_d_i               ( int_if.pad_otpt_d                    ),
    .pad_inpt_vld_i             ( int_if.pad_otpt_vld                  ),
    .pad_inpt_lst_i             ( int_if.pad_otpt_lst                  ),

    .pad_inpt_rdy_o             ( int_if.pad_otpt_ena                  ),
    .expnd_otpt_wj_o            ( int_if.expnd_otpt_wj                 ),
    .expnd_otpt_wjj_o           ( int_if.expnd_otpt_wjj                ),
    .expnd_otpt_lst_o           ( int_if.expnd_otpt_lst                ),
    .expnd_otpt_vld_o           ( int_if.expnd_otpt_vld                )
);   

sm3_cmprss_core U_sm3_cmprss_core(
    .clk                    (clk                    ),
    .rst_n                  (rst_n                  ),


    .expnd_inpt_wj_i            ( int_if.expnd_otpt_wj                  ),
    .expnd_inpt_wjj_i           ( int_if.expnd_otpt_wjj                  ),
    .expnd_inpt_lst_i           ( int_if.expnd_otpt_lst                  ),
    .expnd_inpt_vld_i           ( int_if.expnd_otpt_vld                  ),

    .cmprss_otpt_res_o          ( cmprss_otpt_res               ),
    .cmprss_otpt_vld_o          ( cmprss_otpt_vld               )

);  
    
endmodule

// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/26 
// Design Name: sm3
// Module Name: sm3_expnd_core
// Description:
//      SM3 扩展模块-SM3 扩展核心单元
//      输入位宽：INPT_DW1 定义，支持32/64bit
//      输出位宽：与输入位宽对应
//      特性：预载寄存器（68->65clk(32b)/66->65clk(64b)）,目前仅支持32bit，默认开启
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_expnd_core (
    input                       clk,
    input                       rst_n,

    input   [`INPT_DW1:0]       pad_inpt_d_i,
    input                       pad_inpt_vld_i,
    input                       pad_inpt_lst_i,

    output                      pad_inpt_rdy_o,

    output  [`INPT_DW1:0]       expnd_otpt_wj_o,                    
    output  [`INPT_DW1:0]       expnd_otpt_wjj_o,                    
    output                      expnd_otpt_lst_o,                  
    output                      expnd_otpt_vld_o                    
);

//每时钟输入的数据字数量 32bit位宽：1 64bit位宽：2
`ifdef SM3_INPT_DW_32
    localparam [1:0]            INPT_WORD_NUM               =   2'd1;
`elsif SM3_INPT_DW_64
    localparam [1:0]            INPT_WORD_NUM               =   2'd2;
`endif

localparam                  WORD_INPT_NUM       = 512 / 32;//16
localparam [5:0]            WORD_EXPND_ROUND    = 52;//(68 - 16)

`ifdef SM3_EXPND_PRE_LOAD_REG
    localparam              PRE_BUFF_N = 4;
`endif

//字扩展电路
wire [31:0]             word_wj_expand;
wire [31:0]             word_wjj_otpt;
wire [31:0]             word_wj_expand_tmp_1;
wire [31:0]             word_wj_expand_tmp_2;

//字扩展电路（64bit）
`ifdef SM3_INPT_DW_64
    wire [31:0]             word_wj_expand_w1;
    wire [31:0]             word_wjj_otpt_w1;
    wire [31:0]             word_wj_expand_tmp_1_w1;
    wire [31:0]             word_wj_expand_tmp_2_w1;
`endif

wire                    word_exp_push_reg_ena;  //字拓展，并压入寄存器组使能

//寄存器组 reg
reg [31:0]              word_buff [15:0];   //16字缓冲区  缓存16个32位字
wire                    word_buff_shft_ena;  
wire[31:0]              word_buff_new_push; //寄存器组，新入组变量

//64bit 新增的一个扩展字
`ifdef SM3_INPT_DW_64
    wire[31:0]              word_buff_new_push_w1;
`endif

//预缓冲区
`ifdef SM3_EXPND_PRE_LOAD_REG
    reg [31:0]              word_buff_nb_pre [3:0];//4字 下一字预缓存区
    wire                    word_buff_rpd_shft_ena;  
    wire                    word_buff_nb_pre_shft_ena;  
`endif

//预缓冲区数据数量计数
`ifdef SM3_EXPND_PRE_LOAD_REG
    reg [1:0]               word_buff_nb_pre_cntr;
    wire                    word_buff_nb_pre_cntr_add;
    wire                    word_buff_nb_pre_cntr_clr; 
`endif

//原始字输入计数
reg [3:0]               msg_blk_word_inpt_cntr;  
wire                    msg_blk_word_inpt_cntr_add;
wire                    msg_blk_word_inpt_cntr_clr;

//字扩展输出计数，指本数据块中扩展电路的扩展字输出数量
reg [5:0]               msg_blk_word_exp_cntr;  
wire                    msg_blk_word_exp_cntr_add;
wire                    msg_blk_word_exp_cntr_clr;

//消息扩展主状态机
`define STT_W 8
`define STT_W1 `STT_W - 1

reg [`STT_W1:0]   state;
reg [`STT_W1:0]   nxt_state;

localparam IDLE                     = `STT_W'h1;
localparam INPT_ORGN_5W             = `STT_W'h2;//输入5个原始字w0-w4到寄存器组中
localparam INPT_OTPT                = `STT_W'h4;//输入剩下的11个原始字w5-w15，并输出11对扩展字
localparam EXP_OTPT                 = `STT_W'h8;//扩展并输出扩展字,直至扩展得到第48个扩展字w63
localparam EXP_OTPT_PRE_INPT        = `STT_W'h10;//当w64生成后，开始预接收下一消息块前3个消息字 wn0-wn2，消息字写入预存储寄存器
localparam EXP_OTPT_FIN             = `STT_W'h20;//扩展以及输出结束（输出最后一对扩展字）,接收下一消息块的第4个消息字 wn3,判断预存储器中数据数量
localparam WAT_PRE_INPT_FIN         = `STT_W'h40;//若预存储器数据数量>0 但 <4,等待预寄存器存储完成 4 字
localparam RPD_SHFT                 = `STT_W'h80;//快速移位原始数据,128b位宽的形式，包括预存储寄存器

//SM3填充消息输入反压逻辑
wire                    pad_inpt_d_inpt_rdy;

//消息最后一块标记信号
reg                     msg_lst_blk_flg;
wire                    msg_lst_blk_flg_ena;
wire                    msg_lst_blk_flg_clr;

//SM3填充消息输入反压逻辑，仅在 EXP_OTPT 状态下仅进行扩展，不提供输入
assign                  pad_inpt_d_inpt_rdy = (  state == IDLE 
                                        ||    state == INPT_ORGN_5W
                                        ||    (state == INPT_OTPT && ~(nxt_state   ==  EXP_OTPT))//提前一个周期置低输入有效信号     
                                        ||    state == EXP_OTPT_PRE_INPT     
                                        ||    state == EXP_OTPT_FIN        
                                        ||    state == WAT_PRE_INPT_FIN    
                                        ||    state == RPD_SHFT            
                                        ) ;
  
//原始字输入计数
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        msg_blk_word_inpt_cntr              <= 4'b0;
    end else if(msg_blk_word_inpt_cntr_add)begin
        msg_blk_word_inpt_cntr              <= msg_blk_word_inpt_cntr + INPT_WORD_NUM;
    end else if(msg_blk_word_inpt_cntr_clr)begin
        msg_blk_word_inpt_cntr              <= 4'b0;
    end
end
assign                  msg_blk_word_inpt_cntr_add  = pad_inpt_vld_i; //计数输入消息字
assign                  msg_blk_word_inpt_cntr_clr  = 1'b0; //0-f 对应 16 个消息字，计数自清

//字扩展输出计数
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        msg_blk_word_exp_cntr              <= 6'b0;
    end else if(msg_blk_word_exp_cntr_clr)begin
        msg_blk_word_exp_cntr              <= 6'b0;
    end else if(msg_blk_word_exp_cntr_add)begin
        msg_blk_word_exp_cntr              <= msg_blk_word_exp_cntr + INPT_WORD_NUM;
    end
end
assign                  msg_blk_word_exp_cntr_add  = word_exp_push_reg_ena;//字扩展并移入寄存器使能
assign                  msg_blk_word_exp_cntr_clr  = msg_blk_word_exp_cntr == WORD_EXPND_ROUND;//完成所有扩展次数后清除计数器

`ifdef SM3_EXPND_PRE_LOAD_REG
    //预缓冲区数据数量计数
    always @(posedge clk or negedge rst_n) begin
        if(~rst_n) begin
            word_buff_nb_pre_cntr              <= 2'b0;
        end else if(word_buff_nb_pre_cntr_add)begin
            word_buff_nb_pre_cntr              <= word_buff_nb_pre_cntr + INPT_WORD_NUM;
        end else if(word_buff_nb_pre_cntr_clr)begin
            word_buff_nb_pre_cntr              <= 2'b0;
        end
    end
    assign                  word_buff_nb_pre_cntr_add  = (  state == EXP_OTPT_PRE_INPT 
                                                        ||  state == EXP_OTPT_FIN  
                                                        ||  state == WAT_PRE_INPT_FIN  
                                                        ) && pad_inpt_vld_i;//预输入状态下的外部数据输入有效
    assign                  word_buff_nb_pre_cntr_clr  = state == RPD_SHFT ;//预输入寄存器该状态下被移出
`endif

//消息最后一块标记信号
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        msg_lst_blk_flg              <= 1'b0;
    end else if(msg_lst_blk_flg_ena)begin
        msg_lst_blk_flg              <= 1'b1;
    end else if(msg_lst_blk_flg_clr)begin
        msg_lst_blk_flg              <= 1'b0;
    end
end

assign                  msg_lst_blk_flg_ena  = pad_inpt_lst_i;
assign                  msg_lst_blk_flg_clr  = expnd_otpt_lst_o;

//消息扩展主状态机
always @(*) begin
    case (state)
        IDLE: begin
            if(pad_inpt_vld_i)
                nxt_state   =   INPT_ORGN_5W;
            else
                nxt_state   =   IDLE;
        end
        INPT_ORGN_5W:begin
            if(msg_blk_word_inpt_cntr == 4'd4 && pad_inpt_vld_i) 
                nxt_state   =   INPT_OTPT;//输入前 5 个原始字后，开始一边输入，一边输出
            else
                nxt_state   =   INPT_ORGN_5W;
        end
        INPT_OTPT:begin
            if(msg_blk_word_inpt_cntr == (WORD_INPT_NUM - INPT_WORD_NUM) && pad_inpt_vld_i) 
                nxt_state   =   EXP_OTPT;//输入所有 16 个原始字后，开始向寄存器组输入扩展字
            else
                nxt_state   =   INPT_OTPT;
        end
        EXP_OTPT:begin
            if(msg_blk_word_exp_cntr == 6'd48) 
                nxt_state   =   EXP_OTPT_PRE_INPT; //在生成w63（第48个扩展字后）后，允许下一个块预输入 
            else
                nxt_state   =   EXP_OTPT;
        end
        EXP_OTPT_PRE_INPT:begin
            if(msg_blk_word_exp_cntr == (WORD_EXPND_ROUND - INPT_WORD_NUM)) 
                nxt_state   =   EXP_OTPT_FIN; //在生成51个扩展字后,转入最后一个扩展字 
            else
                nxt_state   =   EXP_OTPT_PRE_INPT;
        end
        EXP_OTPT_FIN:begin
            `ifdef SM3_EXPND_PRE_LOAD_REG
                if(word_buff_nb_pre_cntr == 2'd0 && ~pad_inpt_vld_i) 
                    nxt_state   =   IDLE; //扩展期间无预缓存字，转为idle，等待下次输入
                else if((word_buff_nb_pre_cntr == 3'd4 - INPT_WORD_NUM) && pad_inpt_vld_i)
                    nxt_state   =   RPD_SHFT;//4 个预缓存字，转入 RPD_SHFT
                else 
                    nxt_state   =   WAT_PRE_INPT_FIN;//存在预缓存字，转入 WAT_PRE_INPT_FIN，等待条件满足
            `else
                nxt_state   =   IDLE;
            `endif
        end
        WAT_PRE_INPT_FIN:begin
            `ifdef SM3_EXPND_PRE_LOAD_REG
                if((word_buff_nb_pre_cntr == 3'd4 - INPT_WORD_NUM) && pad_inpt_vld_i) 
                    nxt_state   =   RPD_SHFT; //4 个预缓存字，转入 RPD_SHFT
                else 
                    nxt_state   =   WAT_PRE_INPT_FIN;//存在预缓存字，转入WAT_PRE_INPT_FIN
            `else
                nxt_state   =   IDLE;
            `endif
        end
        RPD_SHFT:begin
            `ifdef SM3_EXPND_PRE_LOAD_REG
                if(pad_inpt_vld_i) 
                    nxt_state   =   INPT_OTPT; //5个原始字输入完毕，开始一边输入，一边输出
                else
                    nxt_state   =   RPD_SHFT;//等待第5个原始字
            `else
                nxt_state   =   IDLE;
            `endif
        end
        default: 
            nxt_state   =   IDLE;
    endcase
end

always @(posedge clk or negedge rst_n) begin
    if(~rst_n)
        state   <=  `STT_W'b1;
    else begin
        state   <=  nxt_state;
    end  
end

//扩展电路
assign                  word_wj_expand_tmp_1        =   word_buff[0] ^ word_buff[7] ^ {word_buff[13][16:0],word_buff[13][31:17]};
assign                  word_wj_expand_tmp_2        =   {word_wj_expand_tmp_1 ^ {word_wj_expand_tmp_1[16:0],word_wj_expand_tmp_1[31:17]} 
                                                                                ^ {word_wj_expand_tmp_1[8:0],word_wj_expand_tmp_1[31:9]}};

assign                  word_wj_expand              =   word_wj_expand_tmp_2 ^ word_buff[10] ^ {word_buff[3][24:0],word_buff[3][31:25]};

`ifdef SM3_INPT_DW_64
    assign                  word_wj_expand_tmp_1_w1        =   word_buff[1] ^ word_buff[8] ^ {word_buff[14][16:0],word_buff[14][31:17]};
    assign                  word_wj_expand_tmp_2_w1        =   {word_wj_expand_tmp_1_w1 ^ {word_wj_expand_tmp_1_w1[16:0],word_wj_expand_tmp_1_w1[31:17]} 
                                                                                    ^ {word_wj_expand_tmp_1_w1[8:0],word_wj_expand_tmp_1_w1[31:9]}};

    assign                  word_wj_expand_w1              =   word_wj_expand_tmp_2_w1 ^ word_buff[11] ^ {word_buff[4][24:0],word_buff[4][31:25]};
`endif

`ifdef SM3_INPT_DW_32
    assign                  word_wjj_otpt                 =   word_buff[11] ^ word_buff[15];
`elsif SM3_INPT_DW_64
    assign                  word_wjj_otpt                 =   word_buff[10] ^ word_buff[14];
    assign                  word_wjj_otpt_w1              =   word_buff[11] ^ word_buff[15];
`endif

    
//扩展电路输出至主寄存器使能
assign                  word_exp_push_reg_ena       =   (state == EXP_OTPT         
                                                    ||   state == EXP_OTPT_PRE_INPT
                                                    ||   state == EXP_OTPT_FIN     
                                                        );

// 根据当前扩展轮数，确定补充进缓冲区的数据类型：原始数据(0-15) 扩展数据(16-67) 0( >67)
assign                  word_buff_new_push          =   (state == IDLE
                                                    ||   state == INPT_ORGN_5W
                                                    ||   state == RPD_SHFT
                                                    ||   state == INPT_OTPT 
                                                    `ifdef SM3_INPT_DW_32
                                                        ) ? pad_inpt_d_i[31:0] : 
                                                    `elsif SM3_INPT_DW_64
                                                        ) ? pad_inpt_d_i[63:32] : 
                                                    `endif
                                                        word_exp_push_reg_ena ? word_wj_expand : 
                                                        32'd0;

`ifdef SM3_INPT_DW_64
    assign                  word_buff_new_push_w1   =   (state == IDLE
                                                    ||   state == INPT_ORGN_5W
                                                    ||   state == RPD_SHFT
                                                    ||   state == INPT_OTPT 
                                                        ) ? pad_inpt_d_i[31:0] : 
                                                        word_exp_push_reg_ena ? word_wj_expand_w1 : 
                                                        32'd0;
`endif

//消息缓冲区 push
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin : buff_init
        integer i;
        for ( i = 0 ; i < WORD_INPT_NUM; i = i + 1) begin:buff_init
            word_buff[i]                <=      32'd0;          
        end
    end
    else if(word_buff_shft_ena)begin : buff_shift // w0 <- w1; w1 <- w2;....w15 <- w_new
        integer i;
        `ifdef SM3_INPT_DW_32
            for ( i = WORD_INPT_NUM - 1 ; i > 0 ; i = i - 1) begin
                word_buff[i-1]                  <=      word_buff[i];    
            end
            word_buff[15]                   <=      word_buff_new_push;  
        `elsif SM3_INPT_DW_64
            for ( i = (WORD_INPT_NUM / INPT_WORD_NUM)- 1 ; i > 0 ; i = i - 1) begin
                word_buff[2*i-1]                    <=      word_buff[2*i+1];    
                word_buff[2*(i-1)]                  <=      word_buff[2*i];    
            end
            {word_buff[14],word_buff[15]}                   <=      {word_buff_new_push,word_buff_new_push_w1};    
        `endif
    end
    `ifdef SM3_EXPND_PRE_LOAD_REG
        else if(word_buff_rpd_shft_ena)begin : buff_rpd_shift //快速移位阶段
            `ifdef SM3_INPT_DW_32
                word_buff[15]                   <=      pad_inpt_d_i;      
                word_buff[14]                   <=      word_buff_nb_pre[3];      
                word_buff[13]                   <=      word_buff_nb_pre[2];      
                word_buff[12]                   <=      word_buff_nb_pre[1];      
                word_buff[11]                   <=      word_buff_nb_pre[0]; 
            `elsif SM3_INPT_DW_64
                {word_buff[14],word_buff[15]}   <=      pad_inpt_d_i;      
                word_buff[13]                   <=      word_buff_nb_pre[2];      
                word_buff[12]                   <=      word_buff_nb_pre[3];      
                word_buff[11]                   <=      word_buff_nb_pre[0];      
                word_buff[10]                   <=      word_buff_nb_pre[1];  
            `endif
                 
        end
    `endif
end

assign                  word_buff_shft_ena      =   (state == IDLE && pad_inpt_vld_i)
                                                ||  (state == INPT_ORGN_5W  && pad_inpt_vld_i)
                                                ||  (state == INPT_OTPT     && pad_inpt_vld_i)
                                                ||  state == EXP_OTPT 
                                                ||  state == EXP_OTPT_PRE_INPT 
                                                ||  state == EXP_OTPT_FIN 
                                                ;//寄存器组左移使能 20.5.13 fix

`ifdef SM3_EXPND_PRE_LOAD_REG
    assign                  word_buff_rpd_shft_ena  =   state == RPD_SHFT && pad_inpt_vld_i; //缓存区快速移位使能 

    //消息预缓冲区
    always @(posedge clk or negedge rst_n) begin
        if(~rst_n) begin : pre_buff_init
            integer i;
            for ( i = 0 ; i < PRE_BUFF_N; i = i + 1) begin : pre_buff_init
                word_buff_nb_pre[i]                <=      32'd0;          
            end
        end
        else if(word_buff_nb_pre_shft_ena)begin : pre_buff_shift // wnb0 <- wnb1....wnb3 <- input
            integer i;
            `ifdef SM3_INPT_DW_32
                for ( i = PRE_BUFF_N - 1 ; i > 0 ; i = i - 1) begin
                    word_buff_nb_pre[i-1]                  <=      word_buff_nb_pre[i];    
                end
                word_buff_nb_pre[PRE_BUFF_N - 1]                   <=      pad_inpt_d_i;    
            `elsif SM3_INPT_DW_64
                for ( i = (PRE_BUFF_N / INPT_WORD_NUM)- 1 ; i > 0 ; i = i - 1) begin
                    word_buff_nb_pre[2*i-1]                    <=      word_buff_nb_pre[2*i+1];    
                    word_buff_nb_pre[2*(i-1)]                  <=      word_buff_nb_pre[2*i];    
                end
                {word_buff_nb_pre[PRE_BUFF_N - 1], word_buff_nb_pre[PRE_BUFF_N - 2]}                  <=      pad_inpt_d_i;    
            `endif
        end
    end

    assign                  word_buff_nb_pre_shft_ena   =   (   state == EXP_OTPT_PRE_INPT
                                                            ||  state == EXP_OTPT_FIN 
                                                            ||  state == WAT_PRE_INPT_FIN 
                                                            ) && pad_inpt_vld_i;//预缓冲区移位使能
`endif

//输出控制
`ifdef SM3_INPT_DW_32
    assign                  expnd_otpt_wj_o                =  word_buff[11];// 从倒数第5个寄存器输出
    assign                  expnd_otpt_wjj_o               =  word_wjj_otpt;
`elsif SM3_INPT_DW_64
    assign                  expnd_otpt_wj_o                =  {word_buff[10],word_buff[11]};
    assign                  expnd_otpt_wjj_o               =  {word_wjj_otpt,word_wjj_otpt_w1};
`endif

assign                  expnd_otpt_vld_o        =  (state == INPT_OTPT && pad_inpt_vld_i) //20.5.13 fix   
                                                ||  state == EXP_OTPT         
                                                ||  state == EXP_OTPT_PRE_INPT
                                                ||  state == EXP_OTPT_FIN
                                                    ;
assign                  expnd_otpt_lst_o        =  msg_lst_blk_flg && state == EXP_OTPT_FIN;
assign                  pad_inpt_rdy_o           =  pad_inpt_d_inpt_rdy; //反压控制

//调试打印信息 debug log
`ifdef SM3_EXPND_SIM_DBG
    generate
        always@(posedge clk) begin
            if(expnd_otpt_vld_o)begin
                `ifdef SM3_INPT_DW_32
                    $display("LOG: EXPND WORD %8h | %8h", expnd_otpt_wj_o[31:0],expnd_otpt_wjj_o[31:0],);
                `elsif SM3_INPT_DW_64
                    $display("LOG: EXPND WORD wj[63:32]:%8h | wj[31:0]:%8h | wjj[63:32]:%8h | wjj[31:0]:%8h"  
                                                                    ,expnd_otpt_wj_o[63:32]
                                                                    ,expnd_otpt_wj_o[31:0]
                                                                    ,expnd_otpt_wjj_o[63:32]
                                                                    ,expnd_otpt_wjj_o[31:0]
                                                                    );
                `endif    
            end	
        end
    endgenerate
`endif
endmodule


// `timescale 1ns / 1ps
// `include "../inc/sm3_cfg"
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/22 
// Design Name: sm3
// Module Name: sm3_if
// Description:
//      SM3 总线定义
//          分为 pad/expnd/cmprss/monitor/top 类型
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
interface sm3_if;
logic                       clk;
logic                       rst_n;
logic [`INPT_DW1:0]         msg_inpt_d;
logic [`INPT_BYTE_DW1:0]    msg_inpt_vld_byte;
logic                       msg_inpt_vld;
logic                       msg_inpt_lst;
logic                       msg_inpt_rdy;
logic                       msg_inpt_rdy_re;

logic                       pad_otpt_ena;
logic [`INPT_DW1:0]         pad_otpt_d;
logic                       pad_otpt_lst;
logic                       pad_otpt_vld;

logic [`INPT_DW1:0]         expnd_otpt_wj; 
logic [`INPT_DW1:0]         expnd_otpt_wjj; 
logic                       expnd_otpt_lst;
logic                       expnd_otpt_vld; 

logic [255:0]               cmprss_otpt_res;
logic                       cmprss_otpt_vld;
logic                       cmprss_vld_re;
logic [7:0]                 cmprss_res_re;

modport PAD (
    input clk,rst_n,msg_inpt_d,msg_inpt_vld_byte,msg_inpt_vld,msg_inpt_lst,pad_otpt_ena,
    output msg_inpt_rdy,pad_otpt_d,pad_otpt_lst,pad_otpt_vld 
);

modport MONITOR (
    input clk,rst_n,msg_inpt_d,msg_inpt_vld_byte,msg_inpt_vld,msg_inpt_lst,pad_otpt_ena,
    msg_inpt_rdy,pad_otpt_d,pad_otpt_lst,pad_otpt_vld 
);

modport EXPND (
    input clk,rst_n,pad_otpt_d,pad_otpt_lst,pad_otpt_vld,
    output expnd_otpt_wj,expnd_otpt_wjj,expnd_otpt_lst,expnd_otpt_vld,pad_otpt_ena
);

modport CMPRSS (
    input clk,rst_n,expnd_otpt_wj,expnd_otpt_wjj,expnd_otpt_lst,expnd_otpt_vld,
    output cmprss_otpt_res,cmprss_otpt_vld
);

modport TOP (
    input clk,rst_n,msg_inpt_d,msg_inpt_vld_byte,msg_inpt_vld,msg_inpt_lst,
    output msg_inpt_rdy,cmprss_otpt_res,cmprss_otpt_vld,msg_inpt_rdy_re,cmprss_vld_re,cmprss_res_re
);

endinterface //sm3_if

// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/26 
// Design Name: sm3
// Module Name: sm3_expnd_core_wrapper
// Description:
//      sm3_expnd_core 的 SV 封装
//          封装 sm3_if 总线接口，类型为 EXPND
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_expnd_core_wrapper (
    sm3_if.EXPND sm3if
);

sm3_expnd_core U_sm3_expnd_core(
    .clk                        (sm3if.clk                    ),
    .rst_n                      (sm3if.rst_n                  ),

    .pad_inpt_d_i            ( sm3if.pad_otpt_d                    ),
    .pad_inpt_vld_i          ( sm3if.pad_otpt_vld                  ),
    .pad_inpt_lst_i          ( sm3if.pad_otpt_lst                  ),

    .pad_inpt_rdy_o          ( sm3if.pad_otpt_ena                  ),
    .expnd_otpt_wj_o         ( sm3if.expnd_otpt_wj                 ),
    .expnd_otpt_wjj_o        ( sm3if.expnd_otpt_wjj                ),
    .expnd_otpt_lst_o        ( sm3if.expnd_otpt_lst                ),
    .expnd_otpt_vld_o        ( sm3if.expnd_otpt_vld                )
);   
    
endmodule

// `timescale 1ns / 1ps
// `include "./inc/sm3_cfg.v"
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/19 
// Design Name: sm3
// Module Name: sm3_pad_core
// Description:
//      SM3 填充模块-SM3 填充核心单元
//      输入位宽：INPT_DW1 定义，支持32/64
//      输出位宽：与输入位宽一致
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_pad_core (
    input                       clk,
    input                       rst_n,

    input   [`INPT_DW1:0]       msg_inpt_d_i,
    input   [`INPT_BYTE_DW1:0]  msg_inpt_vld_byte_i,
    input                       msg_inpt_vld_i,
    input                       msg_inpt_lst_i,

    input                       pad_otpt_ena_i,

    output                      msg_inpt_rdy_o,

    output  [`INPT_DW1:0]       pad_otpt_d_o,                    
    output                      pad_otpt_lst_o,                  
    output                      pad_otpt_vld_o                    
);

localparam [15:0]           PAD_BLK_WD_NUM              =   16;
localparam [15:0]           PAD_BLK_BIT_LEN_WD_NUM      =   2;
localparam [15:0]           PAD_BLK_WD_NUM_INIT         =   PAD_BLK_WD_NUM - PAD_BLK_BIT_LEN_WD_NUM;
localparam [ 3:0]           PAD_BLK_WD_NUM_WTHT_LEN     =   PAD_BLK_WD_NUM - PAD_BLK_BIT_LEN_WD_NUM;

//每时钟输入的数据字数量 32bit位宽：1 64bit位宽：2
`ifdef SM3_INPT_DW_32
    localparam [1:0]            INPT_WORD_NUM               =   2'd1;
`elsif SM3_INPT_DW_64
    localparam [1:0]            INPT_WORD_NUM               =   2'd2;
`endif

//最后一个数据的填充图样
`ifdef SM3_INPT_DW_32
    reg  [31:0]             lst_data_pad_mask;
`elsif SM3_INPT_DW_64
    reg  [63:0]             lst_data_pad_mask;
`endif

//对输入数据打拍  beat inpt signals
reg     [`INPT_DW1:0]       msg_inpt_d_r1;
reg     [`INPT_BYTE_DW1:0]  msg_inpt_vld_byte_r1;
reg                         msg_inpt_vld_r1;
reg                         msg_inpt_lst_r1;

//输入字数统计 count inpt words(32bit)
reg [15:0]                  inpt_wd_cntr;
wire                        inpt_wd_cntr_add;
wire                        inpt_wd_cntr_clr;

//输入字节数统计 count inpt byte
wire[60:0]                  inpt_byte_cntr;

//填充字数统计 count padded words
reg [4:0]                   pad_00_wd_cntr;
wire                        pad_00_wd_cntr_inpt_updt; //随数据输入递减 dec with data inpt
wire                        pad_00_wd_cntr_pad_updt;  //随数据填充递减 dec with pad data
wire                        pad_00_wd_cntr_rld;       //对于新消息，装填计数器 reload cntr for new msg   

//输入比特长度 count inpt bit length
wire [63:0]                 inpt_bit_cntr;

//填充后数据输出使能
wire                        pad_otpt_ena;

//统计最后一个数据的有效字节数  cnt vld byte of the last inpt data
reg  [3:0]                  inpt_vld_byte_cnt;
reg  [3:0]                  inpt_vld_byte_cnt_lat;
wire                        inpt_vld_byte_cmplt;                                 

integer i;

//流程状态机
`define STT_W2 10
`define STT_W21 `STT_W2 - 1

reg [`STT_W21:0]   state;
reg [`STT_W21:0]   nxt_state;

localparam IDLE                     = `STT_W2'h1;
localparam INPT_DATA                = `STT_W2'h2;
localparam INPT_PAD_LST_DATA        = `STT_W2'h4;
localparam PAD_10_DATA              = `STT_W2'h8;
localparam PAD_00_DATA              = `STT_W2'h10;
localparam PAD_LEN_H                = `STT_W2'h20;
localparam PAD_LEN_L                = `STT_W2'h40;
localparam ADD_BLK_PAD_00           = `STT_W2'h80;
localparam PAD_00_WAT_NEW_BLK       = `STT_W2'h100;
localparam PAD_10_WAT_NEW_BLK       = `STT_W2'h200;

//对输入数据打拍  beat inpt signals
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        msg_inpt_d_r1               <=  `INPT_DW'b0;
        msg_inpt_vld_byte_r1        <=  'b0;
        msg_inpt_vld_r1             <=  1'b0;
        msg_inpt_lst_r1             <=  1'b0;
    end else begin
        msg_inpt_d_r1               <=  msg_inpt_d_i;
        msg_inpt_vld_byte_r1        <=  msg_inpt_vld_byte_i;
        msg_inpt_vld_r1             <=  msg_inpt_vld_i;
        msg_inpt_lst_r1             <=  msg_inpt_lst_i;
    end
end

//生成最后一个数据的填充图样
always @(*) begin
    `ifdef SM3_INPT_DW_32
        case (inpt_vld_byte_cnt)
            4'd0: lst_data_pad_mask      =   32'h8000_0000;
            4'd1: lst_data_pad_mask      =   32'h0080_0000;
            4'd2: lst_data_pad_mask      =   32'h0000_8000;
            4'd3: lst_data_pad_mask      =   32'h0000_0080;
            4'd4: lst_data_pad_mask      =   32'h0000_0000;
            default: lst_data_pad_mask      =   32'h8000_0000;
        endcase
    `elsif SM3_INPT_DW_64
        case (inpt_vld_byte_cnt)
            4'd0: lst_data_pad_mask      =   64'h8000_0000_0000_0000;
            4'd1: lst_data_pad_mask      =   64'h0080_0000_0000_0000;
            4'd2: lst_data_pad_mask      =   64'h0000_8000_0000_0000;
            4'd3: lst_data_pad_mask      =   64'h0000_0080_0000_0000;
            4'd4: lst_data_pad_mask      =   64'h0000_0000_8000_0000;
            4'd5: lst_data_pad_mask      =   64'h0000_0000_0080_0000;
            4'd6: lst_data_pad_mask      =   64'h0000_0000_0000_8000;
            4'd7: lst_data_pad_mask      =   64'h0000_0000_0000_0080;
            4'd8: lst_data_pad_mask      =   64'h0000_0000_0000_0000;
            default: lst_data_pad_mask      =   64'h8000_0000_0000_0000;
        endcase
    `endif
end


//统计最后一个数据的有效字节数 
always @(*) begin
    inpt_vld_byte_cnt = 4'b0;
    for(i = 0;i <= `INPT_BYTE_DW1;i=i+1) begin
        inpt_vld_byte_cnt = inpt_vld_byte_cnt + msg_inpt_vld_byte_r1[i];
    end
end

assign                  inpt_vld_byte_cmplt =   inpt_vld_byte_cnt == 4 * INPT_WORD_NUM;

//在last信号，锁存 inpt_vld_byte_cnt
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        inpt_vld_byte_cnt_lat   <=  4'd0;
    end
    else if(msg_inpt_lst_r1)begin
        inpt_vld_byte_cnt_lat   <=  inpt_vld_byte_cnt;
    end
end

//输入字数统计
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        inpt_wd_cntr              <= 16'b0;
    end else if(inpt_wd_cntr_add)begin
        inpt_wd_cntr              <= inpt_wd_cntr + INPT_WORD_NUM;
    end else if(inpt_wd_cntr_clr)begin
        inpt_wd_cntr              <= 16'b0;
    end
end
assign                  inpt_wd_cntr_add    = msg_inpt_vld_r1;
assign                  inpt_wd_cntr_clr    = pad_otpt_lst_o;

assign                  inpt_byte_cntr      =   {inpt_wd_cntr,2'd0} + inpt_vld_byte_cnt_lat - {INPT_WORD_NUM,2'd0};
assign                  inpt_bit_cntr       =   {inpt_byte_cntr,3'd0};

//填充字数统计
always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        pad_00_wd_cntr              <= PAD_BLK_WD_NUM_INIT;//16-2=14
    end else if(pad_00_wd_cntr_inpt_updt)begin
        pad_00_wd_cntr              <= pad_00_wd_cntr == INPT_WORD_NUM 
                                    ? PAD_BLK_WD_NUM 
                                    : pad_00_wd_cntr - INPT_WORD_NUM;
    end else if(pad_00_wd_cntr_rld)begin
        pad_00_wd_cntr              <= PAD_BLK_WD_NUM_INIT;
    end else if(pad_00_wd_cntr_pad_updt)begin
        pad_00_wd_cntr              <= pad_00_wd_cntr - INPT_WORD_NUM;
    end
end
assign                  pad_00_wd_cntr_inpt_updt    = msg_inpt_vld_r1;
assign                  pad_00_wd_cntr_pad_updt     = state == PAD_10_DATA || state == PAD_00_DATA || state == ADD_BLK_PAD_00;
assign                  pad_00_wd_cntr_rld          = pad_otpt_lst_o;

//实现流程状态机
always @(*) begin
    nxt_state   =   IDLE;
    case (state)
        IDLE: begin
            if(msg_inpt_vld_i && ~msg_inpt_lst_i)
                nxt_state   =   INPT_DATA;
            else if(msg_inpt_lst_i)//fix 数据周期为1的情况
                nxt_state   =   INPT_PAD_LST_DATA;
            else
                nxt_state   =   IDLE;
        end
        INPT_DATA: begin //直接输出输入数据，无需填充
            if(msg_inpt_lst_i)
                nxt_state   =   INPT_PAD_LST_DATA;
            else
                nxt_state   =   INPT_DATA;
        end
        INPT_PAD_LST_DATA: begin//根据最后一个输入数据的情况，确定填充策略
            if(inpt_vld_byte_cmplt) begin
                // if(inpt_wd_cntr[3:0] == 4'd0 && ~(inpt_wd_cntr == 16'd0))begin
                if(inpt_wd_cntr[3:0] == PAD_BLK_WD_NUM - INPT_WORD_NUM)begin
                    nxt_state   =   PAD_10_WAT_NEW_BLK;//填充以'1'为首的新块
                end else begin//本块中填1
                    nxt_state   =   PAD_10_DATA;
                end
            end
            else if(inpt_wd_cntr[3:0] == PAD_BLK_WD_NUM_WTHT_LEN - INPT_WORD_NUM)//14 - 1/2
                nxt_state   =   PAD_LEN_H;
            else if(inpt_wd_cntr[3:0] < PAD_BLK_WD_NUM_WTHT_LEN - INPT_WORD_NUM)
                nxt_state   =   PAD_00_DATA;
            else if(inpt_wd_cntr[3:0] > PAD_BLK_WD_NUM_WTHT_LEN - INPT_WORD_NUM)
                `ifdef SM3_INPT_DW_32
                    if(inpt_wd_cntr[3:0] == PAD_BLK_WD_NUM_WTHT_LEN)
                        nxt_state   =   ADD_BLK_PAD_00;//（32位专用）为当前块填充最后一个全0双字
                    else
                        nxt_state   =   PAD_00_WAT_NEW_BLK;
                `elsif SM3_INPT_DW_64
                    nxt_state   =   PAD_00_WAT_NEW_BLK;
                `endif
        end
        PAD_10_DATA: begin//填充由1个1和若干个0组成的数据
            if(inpt_wd_cntr[3:0] < PAD_BLK_WD_NUM_WTHT_LEN - INPT_WORD_NUM)//14-2(64b)
                nxt_state   =   PAD_00_DATA;//直接填0
            else if(inpt_wd_cntr[3:0] == PAD_BLK_WD_NUM_WTHT_LEN - INPT_WORD_NUM)
                nxt_state   =   PAD_LEN_H;//填充长度
            else begin //>PAD_BLK_WD_NUM_WTHT_LEN - INPT_WORD_NUM
                `ifdef SM3_INPT_DW_32
                    if(inpt_wd_cntr[3:0] == PAD_BLK_WD_NUM_WTHT_LEN)
                        nxt_state   =   ADD_BLK_PAD_00;//（32位专用）为当前块填充最后一个全0双字
                    else
                        nxt_state   =   PAD_00_WAT_NEW_BLK;
                `elsif SM3_INPT_DW_64
                    nxt_state   =   PAD_00_WAT_NEW_BLK;
                `endif
            end
        end
        ADD_BLK_PAD_00:begin//在新增的填充块之前补一个0字（32位专用）
            nxt_state   =   PAD_00_WAT_NEW_BLK;
        end
        PAD_00_WAT_NEW_BLK: 
            if(~pad_otpt_ena_i) //等待上一块处理完毕后 开始新的一块输出
                nxt_state   =   PAD_00_WAT_NEW_BLK;
            else
                nxt_state   =   PAD_00_DATA;
        PAD_10_WAT_NEW_BLK: //与 PAD_00_WAT_NEW_BLK 状态的区别在于，新块跳转 PAD_10_DATA 添加 10 
            if(~pad_otpt_ena_i) 
                nxt_state   =   PAD_10_WAT_NEW_BLK;
            else
                nxt_state   =   PAD_10_DATA;
        PAD_00_DATA: //填充全 0 数据
            if(pad_00_wd_cntr == INPT_WORD_NUM)
                nxt_state   =   PAD_LEN_H;
            else
                nxt_state   =   PAD_00_DATA;
        PAD_LEN_H: //填充比特长度的高32位/填充整个比特长度
        `ifdef SM3_INPT_DW_32
            nxt_state   =   PAD_LEN_L;
        `elsif SM3_INPT_DW_64
            nxt_state   =   IDLE;
        `endif
        PAD_LEN_L: 
            nxt_state   =   IDLE;
        default: 
            nxt_state   =   IDLE;
    endcase
end

always @(posedge clk or negedge rst_n) begin
    if(~rst_n)
        state   <=  `STT_W2'b1;
    else begin
        state   <=  nxt_state;
    end  
end



assign                      pad_otpt_ena    =     state == PAD_10_DATA          
                                            ||    state == PAD_00_DATA          
                                            ||    state == PAD_LEN_H          
                                            ||    state == PAD_LEN_L          
                                            ||    state == ADD_BLK_PAD_00 ;                                                             
//输出控制
`ifdef SM3_INPT_DW_32
    assign                      pad_otpt_d_o    =   state == PAD_10_DATA ? 32'h8000_0000:
                                                    state == INPT_PAD_LST_DATA? msg_inpt_d_r1 | lst_data_pad_mask:
                                                    state == PAD_00_DATA || state == ADD_BLK_PAD_00? 32'h0:
                                                    state == PAD_LEN_H ? inpt_bit_cntr[63-:32]: 
                                                    state == PAD_LEN_L ? inpt_bit_cntr[31-:32]:
                                                    msg_inpt_d_r1;
    assign                      pad_otpt_lst_o      =   state == PAD_LEN_L;
`elsif SM3_INPT_DW_64
    assign                      pad_otpt_d_o    =   state == PAD_10_DATA ? 64'h8000_0000_0000_0000:
                                                    state == INPT_PAD_LST_DATA? msg_inpt_d_r1 | lst_data_pad_mask:
                                                    state == PAD_00_DATA || state == ADD_BLK_PAD_00? 64'h0:
                                                    state == PAD_LEN_H ? inpt_bit_cntr: 
                                                    msg_inpt_d_r1;
    assign                      pad_otpt_lst_o      =   state == PAD_LEN_H;
`endif

assign                      pad_otpt_vld_o      =   msg_inpt_vld_r1 || pad_otpt_ena;
assign                      msg_inpt_rdy_o      =   pad_otpt_ena_i && (state == IDLE || state == INPT_DATA);

endmodule

// `timescale 1ns / 1ps
`include "sm3_cfg.sv"
//////////////////////////////////////////////////////////////////////////////////
// Author:        ljgibbs / lf_gibbs@163.com
// Create Date: 2020/07/22 
// Design Name: sm3
// Module Name: sm3_pad_core_wrapper
// Description:
//      sm3_pad_core 的 SV 封装
//          封装 sm3_if 总线接口，类型为 PAD
// Dependencies: 
//      inc/sm3_cfg.v
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////////
module sm3_pad_core_wrapper (
    sm3_if.PAD sm3if
);

sm3_pad_core U_sm3_pad_core(
    .clk                    (sm3if.clk                    ),
    .rst_n                  (sm3if.rst_n                  ),

    .msg_inpt_d_i           (sm3if.msg_inpt_d             ),
    .msg_inpt_vld_byte_i    (sm3if.msg_inpt_vld_byte      ),
    .msg_inpt_vld_i         (sm3if.msg_inpt_vld           ),
    .msg_inpt_lst_i         (sm3if.msg_inpt_lst           ),

    .pad_otpt_ena_i         (sm3if.pad_otpt_ena           ),

    .msg_inpt_rdy_o         (sm3if.msg_inpt_rdy           ),

    .pad_otpt_d_o           (sm3if.pad_otpt_d             ),
    .pad_otpt_lst_o         (sm3if.pad_otpt_lst           ),
    .pad_otpt_vld_o         (sm3if.pad_otpt_vld           )
);   
    
endmodule

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package sm3_reg_pkg;

  // Param list
  parameter int ResultData = 8;

  // Address widths within the block
  parameter int BlockAw = 6;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } msg_inpt_lst;
    struct packed {
      logic        q;
      logic        qe;
    } msg_inpt_vld_byte_0;
    struct packed {
      logic        q;
      logic        qe;
    } msg_inpt_vld_byte_1;
    struct packed {
      logic        q;
      logic        qe;
    } msg_inpt_vld_byte_2;
    struct packed {
      logic        q;
      logic        qe;
    } msg_inpt_vld_byte_3;
  } sm3_reg2hw_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } cmprss_otpt_vld;
    struct packed {
      logic        q;
    } msg_inpt_rdy;
  } sm3_reg2hw_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } sm3_reg2hw_message_in_reg_t;

  typedef struct packed {
    logic [31:0] q;
  } sm3_reg2hw_result_out_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } msg_inpt_lst;
    struct packed {
      logic        d;
      logic        de;
    } msg_inpt_vld_byte_0;
    struct packed {
      logic        d;
      logic        de;
    } msg_inpt_vld_byte_1;
    struct packed {
      logic        d;
      logic        de;
    } msg_inpt_vld_byte_2;
    struct packed {
      logic        d;
      logic        de;
    } msg_inpt_vld_byte_3;
  } sm3_hw2reg_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } cmprss_otpt_vld;
    struct packed {
      logic        d;
      logic        de;
    } msg_inpt_rdy;
  } sm3_hw2reg_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } sm3_hw2reg_message_in_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } sm3_hw2reg_result_out_mreg_t;

  // Register -> HW type
  typedef struct packed {
    sm3_reg2hw_ctrl_signals_reg_t ctrl_signals; // [300:291]
    sm3_reg2hw_state_signals_reg_t state_signals; // [290:289]
    sm3_reg2hw_message_in_reg_t message_in; // [288:256]
    sm3_reg2hw_result_out_mreg_t [7:0] result_out; // [255:0]
  } sm3_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    sm3_hw2reg_ctrl_signals_reg_t ctrl_signals; // [310:301]
    sm3_hw2reg_state_signals_reg_t state_signals; // [300:297]
    sm3_hw2reg_message_in_reg_t message_in; // [296:264]
    sm3_hw2reg_result_out_mreg_t [7:0] result_out; // [263:0]
  } sm3_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] SM3_CTRL_SIGNALS_OFFSET = 6'h 0;
  parameter logic [BlockAw-1:0] SM3_STATE_SIGNALS_OFFSET = 6'h 4;
  parameter logic [BlockAw-1:0] SM3_MESSAGE_IN_OFFSET = 6'h 8;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_0_OFFSET = 6'h c;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_1_OFFSET = 6'h 10;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_2_OFFSET = 6'h 14;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_3_OFFSET = 6'h 18;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_4_OFFSET = 6'h 1c;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_5_OFFSET = 6'h 20;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_6_OFFSET = 6'h 24;
  parameter logic [BlockAw-1:0] SM3_RESULT_OUT_7_OFFSET = 6'h 28;

  // Register index
  typedef enum int {
    SM3_CTRL_SIGNALS,
    SM3_STATE_SIGNALS,
    SM3_MESSAGE_IN,
    SM3_RESULT_OUT_0,
    SM3_RESULT_OUT_1,
    SM3_RESULT_OUT_2,
    SM3_RESULT_OUT_3,
    SM3_RESULT_OUT_4,
    SM3_RESULT_OUT_5,
    SM3_RESULT_OUT_6,
    SM3_RESULT_OUT_7
  } sm3_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] SM3_PERMIT [11] = '{
    4'b 0001, // index[ 0] SM3_CTRL_SIGNALS
    4'b 0001, // index[ 1] SM3_STATE_SIGNALS
    4'b 1111, // index[ 2] SM3_MESSAGE_IN
    4'b 1111, // index[ 3] SM3_RESULT_OUT_0
    4'b 1111, // index[ 4] SM3_RESULT_OUT_1
    4'b 1111, // index[ 5] SM3_RESULT_OUT_2
    4'b 1111, // index[ 6] SM3_RESULT_OUT_3
    4'b 1111, // index[ 7] SM3_RESULT_OUT_4
    4'b 1111, // index[ 8] SM3_RESULT_OUT_5
    4'b 1111, // index[ 9] SM3_RESULT_OUT_6
    4'b 1111  // index[10] SM3_RESULT_OUT_7
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module sm3_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output sm3_reg_pkg::sm3_reg2hw_t reg2hw, // Write
  input  sm3_reg_pkg::sm3_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import sm3_reg_pkg::* ;

  localparam int AW = 6;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [10:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(11)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic ctrl_signals_we;
  logic ctrl_signals_msg_inpt_lst_qs;
  logic ctrl_signals_msg_inpt_lst_wd;
  logic ctrl_signals_msg_inpt_vld_byte_0_qs;
  logic ctrl_signals_msg_inpt_vld_byte_0_wd;
  logic ctrl_signals_msg_inpt_vld_byte_1_qs;
  logic ctrl_signals_msg_inpt_vld_byte_1_wd;
  logic ctrl_signals_msg_inpt_vld_byte_2_qs;
  logic ctrl_signals_msg_inpt_vld_byte_2_wd;
  logic ctrl_signals_msg_inpt_vld_byte_3_qs;
  logic ctrl_signals_msg_inpt_vld_byte_3_wd;
  logic state_signals_cmprss_otpt_vld_qs;
  logic state_signals_msg_inpt_rdy_qs;
  logic message_in_we;
  logic [31:0] message_in_qs;
  logic [31:0] message_in_wd;
  logic [31:0] result_out_0_qs;
  logic [31:0] result_out_1_qs;
  logic [31:0] result_out_2_qs;
  logic [31:0] result_out_3_qs;
  logic [31:0] result_out_4_qs;
  logic [31:0] result_out_5_qs;
  logic [31:0] result_out_6_qs;
  logic [31:0] result_out_7_qs;

  // Register instances
  // R[ctrl_signals]: V(False)
  logic ctrl_signals_qe;
  logic [4:0] ctrl_signals_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_ctrl_signals0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&ctrl_signals_flds_we),
    .q_o(ctrl_signals_qe)
  );
  //   F[msg_inpt_lst]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_msg_inpt_lst (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_msg_inpt_lst_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.msg_inpt_lst.de),
    .d      (hw2reg.ctrl_signals.msg_inpt_lst.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[0]),
    .q      (reg2hw.ctrl_signals.msg_inpt_lst.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_msg_inpt_lst_qs)
  );
  assign reg2hw.ctrl_signals.msg_inpt_lst.qe = ctrl_signals_qe;

  //   F[msg_inpt_vld_byte_0]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_msg_inpt_vld_byte_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_msg_inpt_vld_byte_0_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.msg_inpt_vld_byte_0.de),
    .d      (hw2reg.ctrl_signals.msg_inpt_vld_byte_0.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[1]),
    .q      (reg2hw.ctrl_signals.msg_inpt_vld_byte_0.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_msg_inpt_vld_byte_0_qs)
  );
  assign reg2hw.ctrl_signals.msg_inpt_vld_byte_0.qe = ctrl_signals_qe;

  //   F[msg_inpt_vld_byte_1]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_msg_inpt_vld_byte_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_msg_inpt_vld_byte_1_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.msg_inpt_vld_byte_1.de),
    .d      (hw2reg.ctrl_signals.msg_inpt_vld_byte_1.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[2]),
    .q      (reg2hw.ctrl_signals.msg_inpt_vld_byte_1.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_msg_inpt_vld_byte_1_qs)
  );
  assign reg2hw.ctrl_signals.msg_inpt_vld_byte_1.qe = ctrl_signals_qe;

  //   F[msg_inpt_vld_byte_2]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_msg_inpt_vld_byte_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_msg_inpt_vld_byte_2_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.msg_inpt_vld_byte_2.de),
    .d      (hw2reg.ctrl_signals.msg_inpt_vld_byte_2.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[3]),
    .q      (reg2hw.ctrl_signals.msg_inpt_vld_byte_2.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_msg_inpt_vld_byte_2_qs)
  );
  assign reg2hw.ctrl_signals.msg_inpt_vld_byte_2.qe = ctrl_signals_qe;

  //   F[msg_inpt_vld_byte_3]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_msg_inpt_vld_byte_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_msg_inpt_vld_byte_3_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.msg_inpt_vld_byte_3.de),
    .d      (hw2reg.ctrl_signals.msg_inpt_vld_byte_3.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[4]),
    .q      (reg2hw.ctrl_signals.msg_inpt_vld_byte_3.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_msg_inpt_vld_byte_3_qs)
  );
  assign reg2hw.ctrl_signals.msg_inpt_vld_byte_3.qe = ctrl_signals_qe;


  // R[state_signals]: V(False)
  //   F[cmprss_otpt_vld]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_cmprss_otpt_vld (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.cmprss_otpt_vld.de),
    .d      (hw2reg.state_signals.cmprss_otpt_vld.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.cmprss_otpt_vld.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_cmprss_otpt_vld_qs)
  );

  //   F[msg_inpt_rdy]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_msg_inpt_rdy (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.msg_inpt_rdy.de),
    .d      (hw2reg.state_signals.msg_inpt_rdy.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.msg_inpt_rdy.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_msg_inpt_rdy_qs)
  );


  // R[message_in]: V(False)
  logic message_in_qe;
  logic [0:0] message_in_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_message_in0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&message_in_flds_we),
    .q_o(message_in_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_message_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (message_in_we),
    .wd     (message_in_wd),

    // from internal hardware
    .de     (hw2reg.message_in.de),
    .d      (hw2reg.message_in.d),

    // to internal hardware
    .qe     (message_in_flds_we[0]),
    .q      (reg2hw.message_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (message_in_qs)
  );
  assign reg2hw.message_in.qe = message_in_qe;


  // Subregister 0 of Multireg result_out
  // R[result_out_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[0].de),
    .d      (hw2reg.result_out[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_0_qs)
  );


  // Subregister 1 of Multireg result_out
  // R[result_out_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[1].de),
    .d      (hw2reg.result_out[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_1_qs)
  );


  // Subregister 2 of Multireg result_out
  // R[result_out_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[2].de),
    .d      (hw2reg.result_out[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_2_qs)
  );


  // Subregister 3 of Multireg result_out
  // R[result_out_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[3].de),
    .d      (hw2reg.result_out[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_3_qs)
  );


  // Subregister 4 of Multireg result_out
  // R[result_out_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[4].de),
    .d      (hw2reg.result_out[4].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_4_qs)
  );


  // Subregister 5 of Multireg result_out
  // R[result_out_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[5].de),
    .d      (hw2reg.result_out[5].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_5_qs)
  );


  // Subregister 6 of Multireg result_out
  // R[result_out_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[6].de),
    .d      (hw2reg.result_out[6].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_6_qs)
  );


  // Subregister 7 of Multireg result_out
  // R[result_out_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[7].de),
    .d      (hw2reg.result_out[7].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_7_qs)
  );



  logic [10:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == SM3_CTRL_SIGNALS_OFFSET);
    addr_hit[ 1] = (reg_addr == SM3_STATE_SIGNALS_OFFSET);
    addr_hit[ 2] = (reg_addr == SM3_MESSAGE_IN_OFFSET);
    addr_hit[ 3] = (reg_addr == SM3_RESULT_OUT_0_OFFSET);
    addr_hit[ 4] = (reg_addr == SM3_RESULT_OUT_1_OFFSET);
    addr_hit[ 5] = (reg_addr == SM3_RESULT_OUT_2_OFFSET);
    addr_hit[ 6] = (reg_addr == SM3_RESULT_OUT_3_OFFSET);
    addr_hit[ 7] = (reg_addr == SM3_RESULT_OUT_4_OFFSET);
    addr_hit[ 8] = (reg_addr == SM3_RESULT_OUT_5_OFFSET);
    addr_hit[ 9] = (reg_addr == SM3_RESULT_OUT_6_OFFSET);
    addr_hit[10] = (reg_addr == SM3_RESULT_OUT_7_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(SM3_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(SM3_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(SM3_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(SM3_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(SM3_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(SM3_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(SM3_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(SM3_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(SM3_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(SM3_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(SM3_PERMIT[10] & ~reg_be)))));
  end

  // Generate write-enables
  assign ctrl_signals_we = addr_hit[0] & reg_we & !reg_error;

  assign ctrl_signals_msg_inpt_lst_wd = reg_wdata[0];

  assign ctrl_signals_msg_inpt_vld_byte_0_wd = reg_wdata[1];

  assign ctrl_signals_msg_inpt_vld_byte_1_wd = reg_wdata[2];

  assign ctrl_signals_msg_inpt_vld_byte_2_wd = reg_wdata[3];

  assign ctrl_signals_msg_inpt_vld_byte_3_wd = reg_wdata[4];
  assign message_in_we = addr_hit[2] & reg_we & !reg_error;

  assign message_in_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = ctrl_signals_we;
    reg_we_check[1] = 1'b0;
    reg_we_check[2] = message_in_we;
    reg_we_check[3] = 1'b0;
    reg_we_check[4] = 1'b0;
    reg_we_check[5] = 1'b0;
    reg_we_check[6] = 1'b0;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = 1'b0;
    reg_we_check[9] = 1'b0;
    reg_we_check[10] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = ctrl_signals_msg_inpt_lst_qs;
        reg_rdata_next[1] = ctrl_signals_msg_inpt_vld_byte_0_qs;
        reg_rdata_next[2] = ctrl_signals_msg_inpt_vld_byte_1_qs;
        reg_rdata_next[3] = ctrl_signals_msg_inpt_vld_byte_2_qs;
        reg_rdata_next[4] = ctrl_signals_msg_inpt_vld_byte_3_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = state_signals_cmprss_otpt_vld_qs;
        reg_rdata_next[1] = state_signals_msg_inpt_rdy_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = message_in_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = result_out_0_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = result_out_1_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = result_out_2_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = result_out_3_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = result_out_4_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = result_out_5_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = result_out_6_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = result_out_7_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


`include "prim_assert.sv"


module sm3
  import sm3_reg_pkg::*;
(
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  // Bus interface
  input  tlul_pkg::tl_h2d_t                         tl_i,
  output tlul_pkg::tl_d2h_t                         tl_o
);

  sm3_reg2hw_t               reg2hw;
  sm3_hw2reg_t               hw2reg;
  //wire                       ready_out;

  sm3_reg_top  u_sm3_reg_top (
    .clk_i                             ( clk_i           ),
    .rst_ni                            ( rst_ni          ),
    .tl_i                              ( tl_i            ),
    .hw2reg                            ( hw2reg          ),
    .devmode_i                         ( 1'b1            ),

    .tl_o                              ( tl_o            ),
    .reg2hw                            ( reg2hw          ),
    .intg_err_o                        (                 )
);

assign hw2reg.message_in.de = 1'd0;
assign hw2reg.ctrl_signals.msg_inpt_vld_byte_3.de = 1'd0;
assign hw2reg.ctrl_signals.msg_inpt_vld_byte_2.de = 1'd0;
assign hw2reg.ctrl_signals.msg_inpt_vld_byte_1.de = 1'd0;
assign hw2reg.ctrl_signals.msg_inpt_vld_byte_0.de = 1'd0;
assign hw2reg.ctrl_signals.msg_inpt_lst.de = 1'd0;


sm3_core_top  u_sm3_core_top (
    .clk                     ( clk_i  ),
    .rst_n                   ( rst_ni ),
    .msg_inpt_d              ( reg2hw.message_in.q ),
    .msg_inpt_vld_byte       ( {reg2hw.ctrl_signals.msg_inpt_vld_byte_3.q,reg2hw.ctrl_signals.msg_inpt_vld_byte_2.q,reg2hw.ctrl_signals.msg_inpt_vld_byte_1.q,reg2hw.ctrl_signals.msg_inpt_vld_byte_0.q} ),
    .msg_inpt_vld            ( reg2hw.message_in.qe ),
    .msg_inpt_lst            ( reg2hw.ctrl_signals.msg_inpt_lst.q ),

    .msg_inpt_rdy            ( hw2reg.state_signals.msg_inpt_rdy.d ),
    .cmprss_otpt_res         ( {hw2reg.result_out[7].d,hw2reg.result_out[6].d,hw2reg.result_out[5].d,hw2reg.result_out[4].d,hw2reg.result_out[3].d,hw2reg.result_out[2].d,hw2reg.result_out[1].d,hw2reg.result_out[0].d} ),
    .cmprss_otpt_vld         ( hw2reg.state_signals.cmprss_otpt_vld.d ),
    .msg_inpt_rdy_re         ( hw2reg.state_signals.msg_inpt_rdy.de ),
    .cmprss_vld_re           ( hw2reg.state_signals.cmprss_otpt_vld.de ),
    .cmprss_res_re           ( {hw2reg.result_out[7].de,hw2reg.result_out[6].de,hw2reg.result_out[5].de,hw2reg.result_out[4].de,hw2reg.result_out[3].de,hw2reg.result_out[2].de,hw2reg.result_out[1].de,hw2reg.result_out[0].de} )
);


endmodule


// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/09 21:11:26
// Design Name: 
// Module Name: get_cki
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module get_cki	
	(
		clk,
    	count_round_in,
		cki_out
	);
				
input   clk;
input	[4 :0]	count_round_in;
output	[31:0]	cki_out;

reg [31 : 0] cki_out;
    
always@(posedge clk)
	case(count_round_in)
		5'b0_0000:	cki_out	<=	32'h00070e15;
		5'b0_0001:	cki_out	<=	32'h1c232a31;
		5'b0_0010:	cki_out	<=	32'h383f464d;
		5'b0_0011:	cki_out	<=	32'h545b6269;
		5'b0_0100:	cki_out	<=	32'h70777e85;
		5'b0_0101:	cki_out	<=	32'h8c939aa1;
		5'b0_0110:	cki_out	<=	32'ha8afb6bd;
		5'b0_0111:	cki_out	<=	32'hc4cbd2d9;
		5'b0_1000:	cki_out	<=	32'he0e7eef5;
		5'b0_1001:	cki_out	<=	32'hfc030a11;
		5'b0_1010:	cki_out	<=	32'h181f262d;
		5'b0_1011:	cki_out	<=	32'h343b4249;
		5'b0_1100:	cki_out	<=	32'h50575e65;
		5'b0_1101:	cki_out	<=	32'h6c737a81;
		5'b0_1110:	cki_out	<=	32'h888f969d;
		5'b0_1111:	cki_out	<=	32'ha4abb2b9;
		5'b1_0000:	cki_out	<=	32'hc0c7ced5;
		5'b1_0001:	cki_out	<=	32'hdce3eaf1;
		5'b1_0010:	cki_out	<=	32'hf8ff060d;
		5'b1_0011:	cki_out	<=	32'h141b2229;
		5'b1_0100:	cki_out	<=	32'h30373e45;
		5'b1_0101:	cki_out	<=	32'h4c535a61;
		5'b1_0110:	cki_out	<=	32'h686f767d;
		5'b1_0111:	cki_out	<=	32'h848b9299;
		5'b1_1000:	cki_out	<=	32'ha0a7aeb5;
		5'b1_1001:	cki_out	<=	32'hbcc3cad1;
		5'b1_1010:	cki_out	<=	32'hd8dfe6ed;
		5'b1_1011:	cki_out	<=	32'hf4fb0209;
		5'b1_1100:	cki_out	<=	32'h10171e25;
		5'b1_1101:	cki_out	<=	32'h2c333a41;
		5'b1_1110:	cki_out	<=	32'h484f565d;
		5'b1_1111:	cki_out	<=	32'h646b7279;
		default:	cki_out	<=	32'h0;
	endcase

endmodule


// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/09 20:56:10
// Design Name: FPGA_SM4
// Module Name: key_expansion
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
//      KEY expansion of SM4 encryption algorithm
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module key_expansion
	(
        clk					,
        reset_n				,
        sm4_enable_in		,
        encdec_sel_in       ,
        enable_key_exp_in	,
        user_key_in			,
        user_key_valid_in	,
        key_exp_finished_out,
        rk00_out			,
        rk01_out			,
        rk02_out			,
        rk03_out			,
        rk04_out			,
        rk05_out			,
        rk06_out			,
        rk07_out			,
        rk08_out			,
        rk09_out			,
        rk10_out			,
        rk11_out			,
        rk12_out			,
        rk13_out			,
        rk14_out			,
        rk15_out			,
        rk16_out			,
        rk17_out			,
        rk18_out			,
        rk19_out			,
        rk20_out			,
        rk21_out			,
        rk22_out			,
        rk23_out			,
        rk24_out			,
        rk25_out			,
        rk26_out			,
        rk27_out			,
        rk28_out			,
        rk29_out			,
        rk30_out			,
        rk31_out			
);

input   clk                     ;
input   reset_n                 ;
input   sm4_enable_in           ;
input   encdec_sel_in           ;
input   enable_key_exp_in       ;
input   user_key_valid_in       ;
input   [127: 0]     user_key_in;

output  reg key_exp_finished_out;
output  reg [31 : 0] rk00_out;
output  reg [31 : 0] rk01_out;
output  reg [31 : 0] rk02_out;
output  reg [31 : 0] rk03_out;
output  reg [31 : 0] rk04_out;
output  reg [31 : 0] rk05_out;
output  reg [31 : 0] rk06_out;
output  reg [31 : 0] rk07_out;
output  reg [31 : 0] rk08_out;
output  reg [31 : 0] rk09_out;
output  reg [31 : 0] rk10_out;
output  reg [31 : 0] rk11_out;
output  reg [31 : 0] rk12_out;
output  reg [31 : 0] rk13_out;
output  reg [31 : 0] rk14_out;
output  reg [31 : 0] rk15_out;
output  reg [31 : 0] rk16_out;
output  reg [31 : 0] rk17_out;
output  reg [31 : 0] rk18_out;
output  reg [31 : 0] rk19_out;
output  reg [31 : 0] rk20_out;
output  reg [31 : 0] rk21_out;
output  reg [31 : 0] rk22_out;
output  reg [31 : 0] rk23_out;
output  reg [31 : 0] rk24_out;
output  reg [31 : 0] rk25_out;
output  reg [31 : 0] rk26_out;
output  reg [31 : 0] rk27_out;
output  reg [31 : 0] rk28_out;
output  reg [31 : 0] rk29_out;
output  reg [31 : 0] rk30_out;
output  reg [31 : 0] rk31_out;

reg     [127 : 0]   reg_user_key;
reg     [1   : 0]   current;
reg     [1   : 0]   next;
reg     [4   : 0]   count_round;
reg     [4   : 0]   reg_count_round;
wire    [4   : 0]   count_for_reg;
reg		[127 : 0]	reg_data_after_round;
reg     			reg_user_key_valid = 1'b0;
reg					reg_enable_key_exp;
wire    [31  : 0]  	cki;
wire	[127 : 0]	data_for_round;
wire	[127 : 0]	data_after_round;


always@(posedge clk)
if(!reset_n)
	reg_user_key_valid <= 1'b0;
else 
	reg_user_key_valid <= user_key_valid_in;
        
        
        
always@(posedge clk or negedge reset_n)
begin
	if(~reset_n)
    	reg_enable_key_exp <= 1'b0;
	else 
		reg_enable_key_exp <= enable_key_exp_in;
end

    
`define IDLE          2'b00
`define KEY_EXPANSION 2'b01

always@(posedge clk or negedge reset_n)
if(!reset_n)
	current	<=	`IDLE;
else if(sm4_enable_in)
	current	<=	next;
else
	current	<=	`IDLE;

always@(*) 
begin
	next = `IDLE;
	case(current)
		`IDLE:	
			if(enable_key_exp_in && ~reg_user_key_valid && user_key_valid_in )
				next = `KEY_EXPANSION;
			else
				next = `IDLE;
							
		`KEY_EXPANSION:
			if( reg_count_round == 5'd31)
				next =	`IDLE;
			else
				next =	`KEY_EXPANSION;
										
		default:	
				next =	`IDLE;
	endcase
end


always@(posedge clk or negedge reset_n)
if(!reset_n)
	count_round	<=	5'd0;
else if(next == `KEY_EXPANSION)
	count_round	<=	count_round	+	1'b1;
else 
	count_round <=	5'd0;


always@(posedge clk or negedge reset_n)
begin
    if(!reset_n)
        reg_count_round <= 5'd0;
    else
        reg_count_round <= count_round;
end

    
always@(posedge clk or negedge reset_n)
if(!reset_n)
	key_exp_finished_out <=	1'd0;
else if(~sm4_enable_in || ~enable_key_exp_in && reg_enable_key_exp)    
    key_exp_finished_out <=	1'd0;
else if(current == `KEY_EXPANSION && next == `IDLE)
	key_exp_finished_out <=	1'b1;

always@(posedge clk or negedge reset_n)
if(!reset_n)
	reg_user_key <= 128'h0;
else if(~reg_user_key_valid && user_key_valid_in)
	reg_user_key <= user_key_in;
	
	

assign	data_for_round = reg_count_round != 5'd0 ?	reg_data_after_round : reg_user_key; 


get_cki	u_get_cki
	(
        .clk(clk),
		.count_round_in(count_round),
		.cki_out(cki)
	);


one_round_for_key_exp	u_one_round	
	(	
		.count_round_in(reg_count_round),
		.data_in(data_for_round),
		.ck_parameter_in(cki),
		.result_out(data_after_round)
	);

    
always@(posedge clk or negedge reset_n)
if(!reset_n)
	reg_data_after_round <=	128'd0;
else if(current == `KEY_EXPANSION)
	reg_data_after_round <=	data_after_round;

    
assign count_for_reg = encdec_sel_in == 1'b0 ? reg_count_round : 5'b1_1111 -  reg_count_round;   
    
always@(posedge clk or negedge reset_n)
begin
if(!reset_n) begin
	rk00_out <=	32'd0;
	rk01_out <=	32'd0;
	rk02_out <=	32'd0;
	rk03_out <=	32'd0;
	rk04_out <=	32'd0;
	rk05_out <=	32'd0;
	rk06_out <=	32'd0;
	rk07_out <=	32'd0;
	rk08_out <=	32'd0;
	rk09_out <=	32'd0;
	rk10_out <=	32'd0;
	rk11_out <=	32'd0;
	rk12_out <=	32'd0;
	rk13_out <=	32'd0;
	rk14_out <=	32'd0;
	rk15_out <=	32'd0;
	rk16_out <=	32'd0;
	rk17_out <=	32'd0;
	rk18_out <=	32'd0;
	rk19_out <=	32'd0;
	rk20_out <=	32'd0;
	rk21_out <=	32'd0;
	rk22_out <=	32'd0;
	rk23_out <=	32'd0;
	rk24_out <=	32'd0;
	rk25_out <=	32'd0;
	rk26_out <=	32'd0;
	rk27_out <=	32'd0;
	rk28_out <=	32'd0;
	rk29_out <=	32'd0;
	rk30_out <=	32'd0;
	rk31_out <=	32'd0;
end
else begin
	rk00_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0000	?	data_after_round[31:0]	:	rk00_out;										
	rk01_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0001	?	data_after_round[31:0]	:	rk01_out;
	rk02_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0010	?	data_after_round[31:0]	:	rk02_out;
	rk03_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0011	?	data_after_round[31:0]	:	rk03_out;
	rk04_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0100	?	data_after_round[31:0]	:	rk04_out;
	rk05_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0101	?	data_after_round[31:0]	:	rk05_out;
	rk06_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0110	?	data_after_round[31:0]	:	rk06_out;
	rk07_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_0111	?	data_after_round[31:0]	:	rk07_out;
	rk08_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1000	?	data_after_round[31:0]	:	rk08_out;
	rk09_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1001	?	data_after_round[31:0]	:	rk09_out;
	rk10_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1010	?	data_after_round[31:0]	:	rk10_out;
	rk11_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1011	?	data_after_round[31:0]	:	rk11_out;
	rk12_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1100	?	data_after_round[31:0]	:	rk12_out;
	rk13_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1101	?	data_after_round[31:0]	:	rk13_out;
	rk14_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1110	?	data_after_round[31:0]	:	rk14_out;
	rk15_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b0_1111	?	data_after_round[31:0]	:	rk15_out;
	rk16_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0000	?	data_after_round[31:0]	:	rk16_out;
	rk17_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0001	?	data_after_round[31:0]	:	rk17_out;
	rk18_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0010	?	data_after_round[31:0]	:	rk18_out;
	rk19_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0011	?	data_after_round[31:0]	:	rk19_out;
	rk20_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0100	?	data_after_round[31:0]	:	rk20_out;
	rk21_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0101	?	data_after_round[31:0]	:	rk21_out;
	rk22_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0110	?	data_after_round[31:0]	:	rk22_out;
	rk23_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_0111	?	data_after_round[31:0]	:	rk23_out;
	rk24_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1000	?	data_after_round[31:0]	:	rk24_out;
	rk25_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1001	?	data_after_round[31:0]	:	rk25_out;
	rk26_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1010	?	data_after_round[31:0]	:	rk26_out;
	rk27_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1011	?	data_after_round[31:0]	:	rk27_out;
	rk28_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1100	?	data_after_round[31:0]	:	rk28_out;
	rk29_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1101	?	data_after_round[31:0]	:	rk29_out;
	rk30_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1110	?	data_after_round[31:0]	:	rk30_out;
	rk31_out <=	current == `KEY_EXPANSION && count_for_reg == 5'b1_1111	?	data_after_round[31:0]	:	rk31_out;
	end
end

endmodule







// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/10 10:20:34
// Design Name: 
// Module Name: one_round_for_encdec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module one_round_for_encdec(
		data_in,
		round_key_in,
		result_out
	);
input	[127:0]		data_in;
input	[31:0]		round_key_in;
output	[127:0]		result_out;

wire	[31:0]	word_0;
wire	[31:0]	word_1;
wire	[31:0]	word_2;
wire	[31:0]	word_3;
wire	[31:0]	tmp_0;
wire	[31:0]	tmp_1;
wire	[31:0]	data_for_transform;
wire	[31:0]	data_after_transform;

assign { word_0, word_1, word_2, word_3} = data_in;
			
assign	tmp_0				=	word_1 ^ word_2;
assign	tmp_1				=	word_3 ^ round_key_in;
assign	data_for_transform	=	tmp_0 ^ tmp_1;
assign	result_out			=	{word_1, word_2, word_3, data_after_transform ^ word_0}	;

transform_for_encdec u_transform	
	(
		.data_in(data_for_transform),
		.result_out(data_after_transform)
	);
	
endmodule	


// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/09 21:13:57
// Design Name: 
// Module Name: one_round_for_key_exp
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module one_round_for_key_exp
	(
		count_round_in,
		data_in,
		ck_parameter_in,
		result_out
	);

input	[127 : 0]	data_in;
input	[31  : 0]	ck_parameter_in;
input 	[4   : 0] 	count_round_in;

output	[127 : 0]	result_out;


localparam FK0	=	32'ha3b1bac6;
localparam FK1	=	32'h56aa3350;
localparam FK2	=	32'h677d9197;
localparam FK3	=	32'hb27022dc;

wire	[31:0]	word_0;
wire	[31:0]	word_1;
wire	[31:0]	word_2;
wire	[31:0]	word_3;
wire	[31:0]	tmp_0;
wire	[31:0]	tmp_1;
wire	[31:0]	data_for_xor;
wire	[31:0]	data_for_transform;
wire	[31:0]	data_after_transform_key;
wire	[31:0]	k0;
wire	[31:0]	k1;
wire	[31:0]	k2;
wire	[31:0]	k3;

assign	{	word_0,
			word_1,
			word_2,
			word_3}	=	data_in;

assign	k0					=	word_0^FK0;
assign	k1					=	word_1^FK1;
assign	k2					=	word_2^FK2;
assign	k3					=	word_3^FK3;
assign	data_for_xor		=	ck_parameter_in;
assign	tmp_0				=	count_round_in == 'd0 ? k1^k2 : word_1^word_2;
assign	tmp_1				=	count_round_in == 'd0 ? k3^data_for_xor	: word_3^data_for_xor;
assign	data_for_transform	=	tmp_0 ^ tmp_1;

assign	result_out			=	count_round_in == 'd0	?
								{k1, k2, k3, data_after_transform_key ^ k0}:
								{word_1, word_2, word_3, data_after_transform_key ^ word_0};

transform_for_key_exp	u_transform_key
	(
		.data_in(data_for_transform),
		.data_after_linear_key_out(data_after_transform_key)
	);

	
endmodule
						


module ready_valid (
    input wire clk,
    input wire ready_out,
    input wire encdec_enable_in,
    output reg valid_out
);

always @(posedge clk) begin
    if (ready_out == 1) begin
        valid_out <= 1; // 当ready_out信号为高电平时，A信号为高电平
    end
    else if (encdec_enable_in == 0) begin
        valid_out <= 0; // 当encdec_enable_in信号为低电平时，A信号为低电平
    end
end

endmodule

// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/09 21:25:02
// Design Name: 
// Module Name: sbox_replace
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module sbox_replace	
	(
		data_in,
		result_out														
	);

input	[7:0]	data_in;
output	[7:0]	result_out;

reg		[7:0]	result_out;

always@(*)
	case(data_in)
		8'h00:	result_out	=	8'hd6;
		8'h01:	result_out	=	8'h90;
		8'h02:	result_out	=	8'he9;
		8'h03:	result_out	=	8'hfe;
		8'h04:	result_out	=	8'hcc;
		8'h05:	result_out	=	8'he1;
		8'h06:	result_out	=	8'h3d;
		8'h07:	result_out	=	8'hb7;
		8'h08:	result_out	=	8'h16;
		8'h09:	result_out	=	8'hb6;
		8'h0a:	result_out	=	8'h14;
		8'h0b:	result_out	=	8'hc2;
		8'h0c:	result_out	=	8'h28;
		8'h0d:	result_out	=	8'hfb;
		8'h0e:	result_out	=	8'h2c;
		8'h0f:	result_out	=	8'h05;
		8'h10:	result_out	=	8'h2b;
		8'h11:	result_out	=	8'h67;
		8'h12:	result_out	=	8'h9a;
		8'h13:	result_out	=	8'h76;
		8'h14:	result_out	=	8'h2a;
		8'h15:	result_out	=	8'hbe;
		8'h16:	result_out	=	8'h04;
		8'h17:	result_out	=	8'hc3;
		8'h18:	result_out	=	8'haa;
		8'h19:	result_out	=	8'h44;
		8'h1a:	result_out	=	8'h13;
		8'h1b:	result_out	=	8'h26;
		8'h1c:	result_out	=	8'h49;
		8'h1d:	result_out	=	8'h86;
		8'h1e:	result_out	=	8'h06;
		8'h1f:	result_out	=	8'h99;
		8'h20:	result_out	=	8'h9c;
		8'h21:	result_out	=	8'h42;
		8'h22:	result_out	=	8'h50;
		8'h23:	result_out	=	8'hf4;
		8'h24:	result_out	=	8'h91;
		8'h25:	result_out	=	8'hef;
		8'h26:	result_out	=	8'h98;
		8'h27:	result_out	=	8'h7a;
		8'h28:	result_out	=	8'h33;
		8'h29:	result_out	=	8'h54;
		8'h2a:	result_out	=	8'h0b;
		8'h2b:	result_out	=	8'h43;
		8'h2c:	result_out	=	8'hed;
		8'h2d:	result_out	=	8'hcf;
		8'h2e:	result_out	=	8'hac;
		8'h2f:	result_out	=	8'h62;
		8'h30:	result_out	=	8'he4;
		8'h31:	result_out	=	8'hb3;
		8'h32:	result_out	=	8'h1c;
		8'h33:	result_out	=	8'ha9;
		8'h34:	result_out	=	8'hc9;
		8'h35:	result_out	=	8'h08;
		8'h36:	result_out	=	8'he8;
		8'h37:	result_out	=	8'h95;
		8'h38:	result_out	=	8'h80;
		8'h39:	result_out	=	8'hdf;
		8'h3a:	result_out	=	8'h94;
		8'h3b:	result_out	=	8'hfa;
		8'h3c:	result_out	=	8'h75;
		8'h3d:	result_out	=	8'h8f;
		8'h3e:	result_out	=	8'h3f;
		8'h3f:	result_out	=	8'ha6;
		8'h40:	result_out	=	8'h47;
		8'h41:	result_out	=	8'h07;
		8'h42:	result_out	=	8'ha7;
		8'h43:	result_out	=	8'hfc;
		8'h44:	result_out	=	8'hf3;
		8'h45:	result_out	=	8'h73;
		8'h46:	result_out	=	8'h17;
		8'h47:	result_out	=	8'hba;
		8'h48:	result_out	=	8'h83;
		8'h49:	result_out	=	8'h59;
		8'h4a:	result_out	=	8'h3c;
		8'h4b:	result_out	=	8'h19;
		8'h4c:	result_out	=	8'he6;
		8'h4d:	result_out	=	8'h85;
		8'h4e:	result_out	=	8'h4f;
		8'h4f:	result_out	=	8'ha8;
		8'h50:	result_out	=	8'h68;
		8'h51:	result_out	=	8'h6b;
		8'h52:	result_out	=	8'h81;
		8'h53:	result_out	=	8'hb2;
		8'h54:	result_out	=	8'h71;
		8'h55:	result_out	=	8'h64;
		8'h56:	result_out	=	8'hda;
		8'h57:	result_out	=	8'h8b;
		8'h58:	result_out	=	8'hf8;
		8'h59:	result_out	=	8'heb;
		8'h5a:	result_out	=	8'h0f;
		8'h5b:	result_out	=	8'h4b;
		8'h5c:	result_out	=	8'h70;
		8'h5d:	result_out	=	8'h56;
		8'h5e:	result_out	=	8'h9d;
		8'h5f:	result_out	=	8'h35;
		8'h60:	result_out	=	8'h1e;
		8'h61:	result_out	=	8'h24;
		8'h62:	result_out	=	8'h0e;
		8'h63:	result_out	=	8'h5e;
		8'h64:	result_out	=	8'h63;
		8'h65:	result_out	=	8'h58;
		8'h66:	result_out	=	8'hd1;
		8'h67:	result_out	=	8'ha2;
		8'h68:	result_out	=	8'h25;
		8'h69:	result_out	=	8'h22;
		8'h6a:	result_out	=	8'h7c;
		8'h6b:	result_out	=	8'h3b;
		8'h6c:	result_out	=	8'h01;
		8'h6d:	result_out	=	8'h21;
		8'h6e:	result_out	=	8'h78;
		8'h6f:	result_out	=	8'h87;
		8'h70:	result_out	=	8'hd4;
		8'h71:	result_out	=	8'h00;
		8'h72:	result_out	=	8'h46;
		8'h73:	result_out	=	8'h57;
		8'h74:	result_out	=	8'h9f;
		8'h75:	result_out	=	8'hd3;
		8'h76:	result_out	=	8'h27;
		8'h77:	result_out	=	8'h52;
		8'h78:	result_out	=	8'h4c;
		8'h79:	result_out	=	8'h36;
		8'h7a:	result_out	=	8'h02;
		8'h7b:	result_out	=	8'he7;
		8'h7c:	result_out	=	8'ha0;
		8'h7d:	result_out	=	8'hc4;
		8'h7e:	result_out	=	8'hc8;
		8'h7f:	result_out	=	8'h9e;
		8'h80:	result_out	=	8'hea;
		8'h81:	result_out	=	8'hbf;
		8'h82:	result_out	=	8'h8a;
		8'h83:	result_out	=	8'hd2;
		8'h84:	result_out	=	8'h40;
		8'h85:	result_out	=	8'hc7;
		8'h86:	result_out	=	8'h38;
		8'h87:	result_out	=	8'hb5;
		8'h88:	result_out	=	8'ha3;
		8'h89:	result_out	=	8'hf7;
		8'h8a:	result_out	=	8'hf2;
		8'h8b:	result_out	=	8'hce;
		8'h8c:	result_out	=	8'hf9;
		8'h8d:	result_out	=	8'h61;
		8'h8e:	result_out	=	8'h15;
		8'h8f:	result_out	=	8'ha1;
		8'h90:	result_out	=	8'he0;
		8'h91:	result_out	=	8'hae;
		8'h92:	result_out	=	8'h5d;
		8'h93:	result_out	=	8'ha4;
		8'h94:	result_out	=	8'h9b;
		8'h95:	result_out	=	8'h34;
		8'h96:	result_out	=	8'h1a;
		8'h97:	result_out	=	8'h55;
		8'h98:	result_out	=	8'had;
		8'h99:	result_out	=	8'h93;
		8'h9a:	result_out	=	8'h32;
		8'h9b:	result_out	=	8'h30;
		8'h9c:	result_out	=	8'hf5;
		8'h9d:	result_out	=	8'h8c;
		8'h9e:	result_out	=	8'hb1;
		8'h9f:	result_out	=	8'he3;
		8'ha0:	result_out	=	8'h1d;
		8'ha1:	result_out	=	8'hf6;
		8'ha2:	result_out	=	8'he2;
		8'ha3:	result_out	=	8'h2e;
		8'ha4:	result_out	=	8'h82;
		8'ha5:	result_out	=	8'h66;
		8'ha6:	result_out	=	8'hca;
		8'ha7:	result_out	=	8'h60;
		8'ha8:	result_out	=	8'hc0;
		8'ha9:	result_out	=	8'h29;
		8'haa:	result_out	=	8'h23;
		8'hab:	result_out	=	8'hab;
		8'hac:	result_out	=	8'h0d;
		8'had:	result_out	=	8'h53;
		8'hae:	result_out	=	8'h4e;
		8'haf:	result_out	=	8'h6f;
		8'hb0:	result_out	=	8'hd5;
		8'hb1:	result_out	=	8'hdb;
		8'hb2:	result_out	=	8'h37;
		8'hb3:	result_out	=	8'h45;
		8'hb4:	result_out	=	8'hde;
		8'hb5:	result_out	=	8'hfd;
		8'hb6:	result_out	=	8'h8e;
		8'hb7:	result_out	=	8'h2f;
		8'hb8:	result_out	=	8'h03;
		8'hb9:	result_out	=	8'hff;
		8'hba:	result_out	=	8'h6a;
		8'hbb:	result_out	=	8'h72;
		8'hbc:	result_out	=	8'h6d;
		8'hbd:	result_out	=	8'h6c;
		8'hbe:	result_out	=	8'h5b;
		8'hbf:	result_out	=	8'h51;
		8'hc0:	result_out	=	8'h8d;
		8'hc1:	result_out	=	8'h1b;
		8'hc2:	result_out	=	8'haf;
		8'hc3:	result_out	=	8'h92;
		8'hc4:	result_out	=	8'hbb;
		8'hc5:	result_out	=	8'hdd;
		8'hc6:	result_out	=	8'hbc;
		8'hc7:	result_out	=	8'h7f;
		8'hc8:	result_out	=	8'h11;
		8'hc9:	result_out	=	8'hd9;
		8'hca:	result_out	=	8'h5c;
		8'hcb:	result_out	=	8'h41;
		8'hcc:	result_out	=	8'h1f;
		8'hcd:	result_out	=	8'h10;
		8'hce:	result_out	=	8'h5a;
		8'hcf:	result_out	=	8'hd8;
		8'hd0:	result_out	=	8'h0a;
		8'hd1:	result_out	=	8'hc1;
		8'hd2:	result_out	=	8'h31;
		8'hd3:	result_out	=	8'h88;
		8'hd4:	result_out	=	8'ha5;
		8'hd5:	result_out	=	8'hcd;
		8'hd6:	result_out	=	8'h7b;
		8'hd7:	result_out	=	8'hbd;
		8'hd8:	result_out	=	8'h2d;
		8'hd9:	result_out	=	8'h74;
		8'hda:	result_out	=	8'hd0;
		8'hdb:	result_out	=	8'h12;
		8'hdc:	result_out	=	8'hb8;
		8'hdd:	result_out	=	8'he5;
		8'hde:	result_out	=	8'hb4;
		8'hdf:	result_out	=	8'hb0;
		8'he0:	result_out	=	8'h89;
		8'he1:	result_out	=	8'h69;
		8'he2:	result_out	=	8'h97;
		8'he3:	result_out	=	8'h4a;
		8'he4:	result_out	=	8'h0c;
		8'he5:	result_out	=	8'h96;
		8'he6:	result_out	=	8'h77;
		8'he7:	result_out	=	8'h7e;
		8'he8:	result_out	=	8'h65;
		8'he9:	result_out	=	8'hb9;
		8'hea:	result_out	=	8'hf1;
		8'heb:	result_out	=	8'h09;
		8'hec:	result_out	=	8'hc5;
		8'hed:	result_out	=	8'h6e;
		8'hee:	result_out	=	8'hc6;
		8'hef:	result_out	=	8'h84;
		8'hf0:	result_out	=	8'h18;
		8'hf1:	result_out	=	8'hf0;
		8'hf2:	result_out	=	8'h7d;
		8'hf3:	result_out	=	8'hec;
		8'hf4:	result_out	=	8'h3a;
		8'hf5:	result_out	=	8'hdc;
		8'hf6:	result_out	=	8'h4d;
		8'hf7:	result_out	=	8'h20;
		8'hf8:	result_out	=	8'h79;
		8'hf9:	result_out	=	8'hee;
		8'hfa:	result_out	=	8'h5f;
		8'hfb:	result_out	=	8'h3e;
		8'hfc:	result_out	=	8'hd7;
		8'hfd:	result_out	=	8'hcb;
		8'hfe:	result_out	=	8'h39;
		8'hff:	result_out	=	8'h48;
	endcase

endmodule


// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/10 10:37:43
// Design Name: 
// Module Name: sm4_encdec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module sm4_encdec(
    clk                 ,
    reset_n             ,
    sm4_enable_in       ,
    encdec_enable_in    ,
    key_exp_ready_in    ,
    valid_in            ,
    data_in             ,
    rk_00_in            ,
    rk_01_in            ,
    rk_02_in            ,
    rk_03_in            ,
    rk_04_in            ,
    rk_05_in            ,
    rk_06_in            ,
    rk_07_in            ,
    rk_08_in            ,
    rk_09_in            ,
    rk_10_in            ,
    rk_11_in            ,
    rk_12_in            ,
    rk_13_in            ,
    rk_14_in            ,
    rk_15_in            ,
    rk_16_in            ,
    rk_17_in            ,
    rk_18_in            ,
    rk_19_in            ,
    rk_20_in            ,
    rk_21_in            ,
    rk_22_in            ,
    rk_23_in            ,
    rk_24_in            ,
    rk_25_in            ,
    rk_26_in            ,
    rk_27_in            ,
    rk_28_in            ,
    rk_29_in            ,
    rk_30_in            ,
    rk_31_in            ,
    ready_out           ,
    result_out      
);
    input			 clk		        ;
    input			 reset_n	        ;
    input            sm4_enable_in      ;
    input            encdec_enable_in   ;
    input            key_exp_ready_in   ;
    input            valid_in           ;
    input   [127: 0] data_in            ;
    input   [31 : 0] rk_00_in           ;
    input   [31 : 0] rk_01_in           ;
    input   [31 : 0] rk_02_in           ;
    input   [31 : 0] rk_03_in           ;
    input   [31 : 0] rk_04_in           ;
    input   [31 : 0] rk_05_in           ;
    input   [31 : 0] rk_06_in           ;
    input   [31 : 0] rk_07_in           ;
    input   [31 : 0] rk_08_in           ;
    input   [31 : 0] rk_09_in           ;
    input   [31 : 0] rk_10_in           ;
    input   [31 : 0] rk_11_in           ;
    input   [31 : 0] rk_12_in           ;
    input   [31 : 0] rk_13_in           ;
    input   [31 : 0] rk_14_in           ;
    input   [31 : 0] rk_15_in           ;
    input   [31 : 0] rk_16_in           ;
    input   [31 : 0] rk_17_in           ;
    input   [31 : 0] rk_18_in           ;
    input   [31 : 0] rk_19_in           ;
    input   [31 : 0] rk_20_in           ;
    input   [31 : 0] rk_21_in           ;
    input   [31 : 0] rk_22_in           ;
    input   [31 : 0] rk_23_in           ;
    input   [31 : 0] rk_24_in           ;
    input   [31 : 0] rk_25_in           ;
    input   [31 : 0] rk_26_in           ;
    input   [31 : 0] rk_27_in           ;
    input   [31 : 0] rk_28_in           ;
    input   [31 : 0] rk_29_in           ;
    input   [31 : 0] rk_30_in           ;
    input   [31 : 0] rk_31_in           ;
    output  [127: 0] result_out         ;   
    output           ready_out          ;
    
    reg     [127 : 0] reg_result_00     ;
    reg     [127 : 0] reg_result_01     ;
    reg     [127 : 0] reg_result_02     ;
    reg     [127 : 0] reg_result_03     ;
    reg     [127 : 0] reg_result_04     ;
    reg     [127 : 0] reg_result_05     ;
    reg     [127 : 0] reg_result_06     ;
    reg     [127 : 0] reg_result_07     ;
    reg     [127 : 0] reg_result_08     ;
    reg     [127 : 0] reg_result_09     ;
    reg     [127 : 0] reg_result_10     ;
    reg     [127 : 0] reg_result_11     ;
    reg     [127 : 0] reg_result_12     ;
    reg     [127 : 0] reg_result_13     ;
    reg     [127 : 0] reg_result_14     ;
    reg     [127 : 0] reg_result_15     ;
    reg     [127 : 0] reg_result_16     ;
    reg     [127 : 0] reg_result_17     ;
    reg     [127 : 0] reg_result_18     ;
    reg     [127 : 0] reg_result_19     ;
    reg     [127 : 0] reg_result_20     ;
    reg     [127 : 0] reg_result_21     ;
    reg     [127 : 0] reg_result_22     ;
    reg     [127 : 0] reg_result_23     ;
    reg     [127 : 0] reg_result_24     ;
    reg     [127 : 0] reg_result_25     ;
    reg     [127 : 0] reg_result_26     ;
    reg     [127 : 0] reg_result_27     ;
    reg     [127 : 0] reg_result_28     ;
    reg     [127 : 0] reg_result_29     ;
    reg     [127 : 0] reg_result_30     ;
    reg     [127 : 0] result_out        ;
    reg     [31  : 0] reg_tmp           ;
    wire    [31  : 0] word_0            ;
    wire    [31  : 0] word_1            ;
    wire    [31  : 0] word_2            ;
    wire    [31  : 0] word_3            ;
    wire    [127 : 0] reversed_result_31;
    wire    [127 : 0] result_00         ;
    wire    [127 : 0] result_01         ;
    wire    [127 : 0] result_02         ;
    wire    [127 : 0] result_03         ;
    wire    [127 : 0] result_04         ;
    wire    [127 : 0] result_05         ;
    wire    [127 : 0] result_06         ;
    wire    [127 : 0] result_07         ;
    wire    [127 : 0] result_08         ;
    wire    [127 : 0] result_09         ;
    wire    [127 : 0] result_10         ;
    wire    [127 : 0] result_11         ;
    wire    [127 : 0] result_12         ;
    wire    [127 : 0] result_13         ;
    wire    [127 : 0] result_14         ;
    wire    [127 : 0] result_15         ;
    wire    [127 : 0] result_16         ;
    wire    [127 : 0] result_17         ;
    wire    [127 : 0] result_18         ;
    wire    [127 : 0] result_19         ;
    wire    [127 : 0] result_20         ;
    wire    [127 : 0] result_21         ;
    wire    [127 : 0] result_22         ;
    wire    [127 : 0] result_23         ;
    wire    [127 : 0] result_24         ;
    wire    [127 : 0] result_25         ;
    wire    [127 : 0] result_26         ;
    wire    [127 : 0] result_27         ;
    wire    [127 : 0] result_28         ;
    wire    [127 : 0] result_29         ;
    wire    [127 : 0] result_30         ;
    wire    [127 : 0] result_31         ;
    reg     [1   : 0] current           ;
    reg     [1   : 0] next              ;
    
    `define IDLE                2'b00
    `define WAITING_FOR_KEY     2'b01
    `define ENCRYPTION          2'b10
    
    always@(posedge clk or negedge reset_n)
    if(!reset_n)
        current <= `IDLE;
    else if(sm4_enable_in)
        current <= next;
        
    always@(*)        
        begin
            next = `IDLE;
            case(current)
                `IDLE :
                        if(sm4_enable_in && encdec_enable_in)
                            next = `WAITING_FOR_KEY;
                        else
                            next = `IDLE;
                `WAITING_FOR_KEY :
                        if(key_exp_ready_in)
                            next = `ENCRYPTION;
                        else
                            next = `WAITING_FOR_KEY;
                `ENCRYPTION :
                        if(!encdec_enable_in || !sm4_enable_in)
                            next = `IDLE;
                        else 
                            next = `ENCRYPTION;
                default :
                        next = `IDLE;
            endcase
        end
                
    always@(posedge clk or negedge reset_n)
    if(!reset_n)
        reg_tmp <= 32'b0;
    else if(current == `ENCRYPTION && valid_in)
        reg_tmp <= {reg_tmp[30 : 0], 1'b1};
    else
        reg_tmp <= {reg_tmp[30 : 0], 1'b0};


    assign ready_out = reg_tmp[31];
    
    one_round_for_encdec u_00 ( .data_in(data_in      ), .round_key_in(rk_00_in), .result_out(result_00) );
    one_round_for_encdec u_01 ( .data_in(reg_result_00), .round_key_in(rk_01_in), .result_out(result_01) );
    one_round_for_encdec u_02 ( .data_in(reg_result_01), .round_key_in(rk_02_in), .result_out(result_02) );
    one_round_for_encdec u_03 ( .data_in(reg_result_02), .round_key_in(rk_03_in), .result_out(result_03) );
    one_round_for_encdec u_04 ( .data_in(reg_result_03), .round_key_in(rk_04_in), .result_out(result_04) );
    one_round_for_encdec u_05 ( .data_in(reg_result_04), .round_key_in(rk_05_in), .result_out(result_05) );
    one_round_for_encdec u_06 ( .data_in(reg_result_05), .round_key_in(rk_06_in), .result_out(result_06) );
    one_round_for_encdec u_07 ( .data_in(reg_result_06), .round_key_in(rk_07_in), .result_out(result_07) );
    one_round_for_encdec u_08 ( .data_in(reg_result_07), .round_key_in(rk_08_in), .result_out(result_08) );
    one_round_for_encdec u_09 ( .data_in(reg_result_08), .round_key_in(rk_09_in), .result_out(result_09) );
    one_round_for_encdec u_10 ( .data_in(reg_result_09), .round_key_in(rk_10_in), .result_out(result_10) );
    one_round_for_encdec u_11 ( .data_in(reg_result_10), .round_key_in(rk_11_in), .result_out(result_11) );
    one_round_for_encdec u_12 ( .data_in(reg_result_11), .round_key_in(rk_12_in), .result_out(result_12) );
    one_round_for_encdec u_13 ( .data_in(reg_result_12), .round_key_in(rk_13_in), .result_out(result_13) );
    one_round_for_encdec u_14 ( .data_in(reg_result_13), .round_key_in(rk_14_in), .result_out(result_14) );
    one_round_for_encdec u_15 ( .data_in(reg_result_14), .round_key_in(rk_15_in), .result_out(result_15) );
    one_round_for_encdec u_16 ( .data_in(reg_result_15), .round_key_in(rk_16_in), .result_out(result_16) );
    one_round_for_encdec u_17 ( .data_in(reg_result_16), .round_key_in(rk_17_in), .result_out(result_17) );
    one_round_for_encdec u_18 ( .data_in(reg_result_17), .round_key_in(rk_18_in), .result_out(result_18) );
    one_round_for_encdec u_19 ( .data_in(reg_result_18), .round_key_in(rk_19_in), .result_out(result_19) );
    one_round_for_encdec u_20 ( .data_in(reg_result_19), .round_key_in(rk_20_in), .result_out(result_20) );
    one_round_for_encdec u_21 ( .data_in(reg_result_20), .round_key_in(rk_21_in), .result_out(result_21) );
    one_round_for_encdec u_22 ( .data_in(reg_result_21), .round_key_in(rk_22_in), .result_out(result_22) );
    one_round_for_encdec u_23 ( .data_in(reg_result_22), .round_key_in(rk_23_in), .result_out(result_23) );
    one_round_for_encdec u_24 ( .data_in(reg_result_23), .round_key_in(rk_24_in), .result_out(result_24) );
    one_round_for_encdec u_25 ( .data_in(reg_result_24), .round_key_in(rk_25_in), .result_out(result_25) );
    one_round_for_encdec u_26 ( .data_in(reg_result_25), .round_key_in(rk_26_in), .result_out(result_26) );
    one_round_for_encdec u_27 ( .data_in(reg_result_26), .round_key_in(rk_27_in), .result_out(result_27) );
    one_round_for_encdec u_28 ( .data_in(reg_result_27), .round_key_in(rk_28_in), .result_out(result_28) );
    one_round_for_encdec u_29 ( .data_in(reg_result_28), .round_key_in(rk_29_in), .result_out(result_29) );
    one_round_for_encdec u_30 ( .data_in(reg_result_29), .round_key_in(rk_30_in), .result_out(result_30) );
    one_round_for_encdec u_31 ( .data_in(reg_result_30), .round_key_in(rk_31_in), .result_out(result_31) );
    
    assign { word_0, word_1, word_2, word_3} = result_31;
    assign reversed_result_31 = {word_3, word_2, word_1, word_0};
    
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_00 <= 128'h0; else reg_result_00 <= result_00;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_01 <= 128'h0; else reg_result_01 <= result_01;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_02 <= 128'h0; else reg_result_02 <= result_02;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_03 <= 128'h0; else reg_result_03 <= result_03;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_04 <= 128'h0; else reg_result_04 <= result_04;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_05 <= 128'h0; else reg_result_05 <= result_05;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_06 <= 128'h0; else reg_result_06 <= result_06;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_07 <= 128'h0; else reg_result_07 <= result_07;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_08 <= 128'h0; else reg_result_08 <= result_08;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_09 <= 128'h0; else reg_result_09 <= result_09;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_10 <= 128'h0; else reg_result_10 <= result_10;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_11 <= 128'h0; else reg_result_11 <= result_11;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_12 <= 128'h0; else reg_result_12 <= result_12;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_13 <= 128'h0; else reg_result_13 <= result_13;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_14 <= 128'h0; else reg_result_14 <= result_14;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_15 <= 128'h0; else reg_result_15 <= result_15;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_16 <= 128'h0; else reg_result_16 <= result_16;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_17 <= 128'h0; else reg_result_17 <= result_17;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_18 <= 128'h0; else reg_result_18 <= result_18;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_19 <= 128'h0; else reg_result_19 <= result_19;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_20 <= 128'h0; else reg_result_20 <= result_20;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_21 <= 128'h0; else reg_result_21 <= result_21;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_22 <= 128'h0; else reg_result_22 <= result_22;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_23 <= 128'h0; else reg_result_23 <= result_23;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_24 <= 128'h0; else reg_result_24 <= result_24;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_25 <= 128'h0; else reg_result_25 <= result_25;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_26 <= 128'h0; else reg_result_26 <= result_26;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_27 <= 128'h0; else reg_result_27 <= result_27;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_28 <= 128'h0; else reg_result_28 <= result_28;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_29 <= 128'h0; else reg_result_29 <= result_29;
    always@(posedge clk or negedge reset_n) if(!reset_n) reg_result_30 <= 128'h0; else reg_result_30 <= result_30;
    always@(posedge clk or negedge reset_n) if(!reset_n) result_out    <= 128'h0; else result_out    <= reversed_result_31;
        
                                                    
endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package sm4_reg_pkg;

  // Param list
  parameter int NumRegsData = 4;
  parameter int NumRegsKey = 4;

  // Address widths within the block
  parameter int BlockAw = 6;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } sm4_enable_in;
    struct packed {
      logic        q;
      logic        qe;
    } encdec_sel_in;
    struct packed {
      logic        q;
      logic        qe;
    } enable_key_exp_in;
    struct packed {
      logic        q;
      logic        qe;
    } user_key_valid_in;
    struct packed {
      logic        q;
      logic        qe;
    } encdec_enable_in;
    struct packed {
      logic        q;
      logic        qe;
    } valid_in;
  } sm4_reg2hw_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } key_exp_ready_out;
    struct packed {
      logic        q;
    } valid_out;
  } sm4_reg2hw_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } sm4_reg2hw_key_mreg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } sm4_reg2hw_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } sm4_reg2hw_result_out_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } sm4_enable_in;
    struct packed {
      logic        d;
      logic        de;
    } encdec_sel_in;
    struct packed {
      logic        d;
      logic        de;
    } enable_key_exp_in;
    struct packed {
      logic        d;
      logic        de;
    } user_key_valid_in;
    struct packed {
      logic        d;
      logic        de;
    } encdec_enable_in;
    struct packed {
      logic        d;
      logic        de;
    } valid_in;
  } sm4_hw2reg_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } key_exp_ready_out;
    struct packed {
      logic        d;
      logic        de;
    } valid_out;
  } sm4_hw2reg_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } sm4_hw2reg_key_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } sm4_hw2reg_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } sm4_hw2reg_result_out_mreg_t;

  // Register -> HW type
  typedef struct packed {
    sm4_reg2hw_ctrl_signals_reg_t ctrl_signals; // [405:394]
    sm4_reg2hw_state_signals_reg_t state_signals; // [393:392]
    sm4_reg2hw_key_mreg_t [3:0] key; // [391:260]
    sm4_reg2hw_data_in_mreg_t [3:0] data_in; // [259:128]
    sm4_reg2hw_result_out_mreg_t [3:0] result_out; // [127:0]
  } sm4_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    sm4_hw2reg_ctrl_signals_reg_t ctrl_signals; // [411:400]
    sm4_hw2reg_state_signals_reg_t state_signals; // [399:396]
    sm4_hw2reg_key_mreg_t [3:0] key; // [395:264]
    sm4_hw2reg_data_in_mreg_t [3:0] data_in; // [263:132]
    sm4_hw2reg_result_out_mreg_t [3:0] result_out; // [131:0]
  } sm4_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] SM4_CTRL_SIGNALS_OFFSET = 6'h 0;
  parameter logic [BlockAw-1:0] SM4_STATE_SIGNALS_OFFSET = 6'h 4;
  parameter logic [BlockAw-1:0] SM4_KEY_0_OFFSET = 6'h 8;
  parameter logic [BlockAw-1:0] SM4_KEY_1_OFFSET = 6'h c;
  parameter logic [BlockAw-1:0] SM4_KEY_2_OFFSET = 6'h 10;
  parameter logic [BlockAw-1:0] SM4_KEY_3_OFFSET = 6'h 14;
  parameter logic [BlockAw-1:0] SM4_DATA_IN_0_OFFSET = 6'h 18;
  parameter logic [BlockAw-1:0] SM4_DATA_IN_1_OFFSET = 6'h 1c;
  parameter logic [BlockAw-1:0] SM4_DATA_IN_2_OFFSET = 6'h 20;
  parameter logic [BlockAw-1:0] SM4_DATA_IN_3_OFFSET = 6'h 24;
  parameter logic [BlockAw-1:0] SM4_RESULT_OUT_0_OFFSET = 6'h 28;
  parameter logic [BlockAw-1:0] SM4_RESULT_OUT_1_OFFSET = 6'h 2c;
  parameter logic [BlockAw-1:0] SM4_RESULT_OUT_2_OFFSET = 6'h 30;
  parameter logic [BlockAw-1:0] SM4_RESULT_OUT_3_OFFSET = 6'h 34;

  // Register index
  typedef enum int {
    SM4_CTRL_SIGNALS,
    SM4_STATE_SIGNALS,
    SM4_KEY_0,
    SM4_KEY_1,
    SM4_KEY_2,
    SM4_KEY_3,
    SM4_DATA_IN_0,
    SM4_DATA_IN_1,
    SM4_DATA_IN_2,
    SM4_DATA_IN_3,
    SM4_RESULT_OUT_0,
    SM4_RESULT_OUT_1,
    SM4_RESULT_OUT_2,
    SM4_RESULT_OUT_3
  } sm4_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] SM4_PERMIT [14] = '{
    4'b 0001, // index[ 0] SM4_CTRL_SIGNALS
    4'b 0001, // index[ 1] SM4_STATE_SIGNALS
    4'b 1111, // index[ 2] SM4_KEY_0
    4'b 1111, // index[ 3] SM4_KEY_1
    4'b 1111, // index[ 4] SM4_KEY_2
    4'b 1111, // index[ 5] SM4_KEY_3
    4'b 1111, // index[ 6] SM4_DATA_IN_0
    4'b 1111, // index[ 7] SM4_DATA_IN_1
    4'b 1111, // index[ 8] SM4_DATA_IN_2
    4'b 1111, // index[ 9] SM4_DATA_IN_3
    4'b 1111, // index[10] SM4_RESULT_OUT_0
    4'b 1111, // index[11] SM4_RESULT_OUT_1
    4'b 1111, // index[12] SM4_RESULT_OUT_2
    4'b 1111  // index[13] SM4_RESULT_OUT_3
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module sm4_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output sm4_reg_pkg::sm4_reg2hw_t reg2hw, // Write
  input  sm4_reg_pkg::sm4_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import sm4_reg_pkg::* ;

  localparam int AW = 6;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [13:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(14)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic ctrl_signals_we;
  logic ctrl_signals_sm4_enable_in_qs;
  logic ctrl_signals_sm4_enable_in_wd;
  logic ctrl_signals_encdec_sel_in_qs;
  logic ctrl_signals_encdec_sel_in_wd;
  logic ctrl_signals_enable_key_exp_in_qs;
  logic ctrl_signals_enable_key_exp_in_wd;
  logic ctrl_signals_user_key_valid_in_qs;
  logic ctrl_signals_user_key_valid_in_wd;
  logic ctrl_signals_encdec_enable_in_qs;
  logic ctrl_signals_encdec_enable_in_wd;
  logic ctrl_signals_valid_in_qs;
  logic ctrl_signals_valid_in_wd;
  logic state_signals_key_exp_ready_out_qs;
  logic state_signals_valid_out_qs;
  logic key_0_we;
  logic [31:0] key_0_qs;
  logic [31:0] key_0_wd;
  logic key_1_we;
  logic [31:0] key_1_qs;
  logic [31:0] key_1_wd;
  logic key_2_we;
  logic [31:0] key_2_qs;
  logic [31:0] key_2_wd;
  logic key_3_we;
  logic [31:0] key_3_qs;
  logic [31:0] key_3_wd;
  logic data_in_0_we;
  logic [31:0] data_in_0_qs;
  logic [31:0] data_in_0_wd;
  logic data_in_1_we;
  logic [31:0] data_in_1_qs;
  logic [31:0] data_in_1_wd;
  logic data_in_2_we;
  logic [31:0] data_in_2_qs;
  logic [31:0] data_in_2_wd;
  logic data_in_3_we;
  logic [31:0] data_in_3_qs;
  logic [31:0] data_in_3_wd;
  logic [31:0] result_out_0_qs;
  logic [31:0] result_out_1_qs;
  logic [31:0] result_out_2_qs;
  logic [31:0] result_out_3_qs;

  // Register instances
  // R[ctrl_signals]: V(False)
  logic ctrl_signals_qe;
  logic [5:0] ctrl_signals_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_ctrl_signals0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&ctrl_signals_flds_we),
    .q_o(ctrl_signals_qe)
  );
  //   F[sm4_enable_in]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_sm4_enable_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_sm4_enable_in_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.sm4_enable_in.de),
    .d      (hw2reg.ctrl_signals.sm4_enable_in.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[0]),
    .q      (reg2hw.ctrl_signals.sm4_enable_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_sm4_enable_in_qs)
  );
  assign reg2hw.ctrl_signals.sm4_enable_in.qe = ctrl_signals_qe;

  //   F[encdec_sel_in]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_encdec_sel_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_encdec_sel_in_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.encdec_sel_in.de),
    .d      (hw2reg.ctrl_signals.encdec_sel_in.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[1]),
    .q      (reg2hw.ctrl_signals.encdec_sel_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_encdec_sel_in_qs)
  );
  assign reg2hw.ctrl_signals.encdec_sel_in.qe = ctrl_signals_qe;

  //   F[enable_key_exp_in]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_enable_key_exp_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_enable_key_exp_in_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.enable_key_exp_in.de),
    .d      (hw2reg.ctrl_signals.enable_key_exp_in.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[2]),
    .q      (reg2hw.ctrl_signals.enable_key_exp_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_enable_key_exp_in_qs)
  );
  assign reg2hw.ctrl_signals.enable_key_exp_in.qe = ctrl_signals_qe;

  //   F[user_key_valid_in]: 3:3
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_user_key_valid_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_user_key_valid_in_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.user_key_valid_in.de),
    .d      (hw2reg.ctrl_signals.user_key_valid_in.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[3]),
    .q      (reg2hw.ctrl_signals.user_key_valid_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_user_key_valid_in_qs)
  );
  assign reg2hw.ctrl_signals.user_key_valid_in.qe = ctrl_signals_qe;

  //   F[encdec_enable_in]: 4:4
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_encdec_enable_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_encdec_enable_in_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.encdec_enable_in.de),
    .d      (hw2reg.ctrl_signals.encdec_enable_in.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[4]),
    .q      (reg2hw.ctrl_signals.encdec_enable_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_encdec_enable_in_qs)
  );
  assign reg2hw.ctrl_signals.encdec_enable_in.qe = ctrl_signals_qe;

  //   F[valid_in]: 5:5
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_valid_in (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_valid_in_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.valid_in.de),
    .d      (hw2reg.ctrl_signals.valid_in.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[5]),
    .q      (reg2hw.ctrl_signals.valid_in.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_valid_in_qs)
  );
  assign reg2hw.ctrl_signals.valid_in.qe = ctrl_signals_qe;


  // R[state_signals]: V(False)
  //   F[key_exp_ready_out]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_key_exp_ready_out (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.key_exp_ready_out.de),
    .d      (hw2reg.state_signals.key_exp_ready_out.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.key_exp_ready_out.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_key_exp_ready_out_qs)
  );

  //   F[valid_out]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_valid_out (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.valid_out.de),
    .d      (hw2reg.state_signals.valid_out.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.valid_out.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_valid_out_qs)
  );


  // Subregister 0 of Multireg key
  // R[key_0]: V(False)
  logic key_0_qe;
  logic [0:0] key_0_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_key0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&key_0_flds_we),
    .q_o(key_0_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_key_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (key_0_we),
    .wd     (key_0_wd),

    // from internal hardware
    .de     (hw2reg.key[0].de),
    .d      (hw2reg.key[0].d),

    // to internal hardware
    .qe     (key_0_flds_we[0]),
    .q      (reg2hw.key[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (key_0_qs)
  );
  assign reg2hw.key[0].qe = key_0_qe;


  // Subregister 1 of Multireg key
  // R[key_1]: V(False)
  logic key_1_qe;
  logic [0:0] key_1_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_key1_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&key_1_flds_we),
    .q_o(key_1_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_key_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (key_1_we),
    .wd     (key_1_wd),

    // from internal hardware
    .de     (hw2reg.key[1].de),
    .d      (hw2reg.key[1].d),

    // to internal hardware
    .qe     (key_1_flds_we[0]),
    .q      (reg2hw.key[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (key_1_qs)
  );
  assign reg2hw.key[1].qe = key_1_qe;


  // Subregister 2 of Multireg key
  // R[key_2]: V(False)
  logic key_2_qe;
  logic [0:0] key_2_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_key2_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&key_2_flds_we),
    .q_o(key_2_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_key_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (key_2_we),
    .wd     (key_2_wd),

    // from internal hardware
    .de     (hw2reg.key[2].de),
    .d      (hw2reg.key[2].d),

    // to internal hardware
    .qe     (key_2_flds_we[0]),
    .q      (reg2hw.key[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (key_2_qs)
  );
  assign reg2hw.key[2].qe = key_2_qe;


  // Subregister 3 of Multireg key
  // R[key_3]: V(False)
  logic key_3_qe;
  logic [0:0] key_3_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_key3_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&key_3_flds_we),
    .q_o(key_3_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_key_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (key_3_we),
    .wd     (key_3_wd),

    // from internal hardware
    .de     (hw2reg.key[3].de),
    .d      (hw2reg.key[3].d),

    // to internal hardware
    .qe     (key_3_flds_we[0]),
    .q      (reg2hw.key[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (key_3_qs)
  );
  assign reg2hw.key[3].qe = key_3_qe;


  // Subregister 0 of Multireg data_in
  // R[data_in_0]: V(False)
  logic data_in_0_qe;
  logic [0:0] data_in_0_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_0_flds_we),
    .q_o(data_in_0_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_0_we),
    .wd     (data_in_0_wd),

    // from internal hardware
    .de     (hw2reg.data_in[0].de),
    .d      (hw2reg.data_in[0].d),

    // to internal hardware
    .qe     (data_in_0_flds_we[0]),
    .q      (reg2hw.data_in[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_0_qs)
  );
  assign reg2hw.data_in[0].qe = data_in_0_qe;


  // Subregister 1 of Multireg data_in
  // R[data_in_1]: V(False)
  logic data_in_1_qe;
  logic [0:0] data_in_1_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in1_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_1_flds_we),
    .q_o(data_in_1_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_1_we),
    .wd     (data_in_1_wd),

    // from internal hardware
    .de     (hw2reg.data_in[1].de),
    .d      (hw2reg.data_in[1].d),

    // to internal hardware
    .qe     (data_in_1_flds_we[0]),
    .q      (reg2hw.data_in[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_1_qs)
  );
  assign reg2hw.data_in[1].qe = data_in_1_qe;


  // Subregister 2 of Multireg data_in
  // R[data_in_2]: V(False)
  logic data_in_2_qe;
  logic [0:0] data_in_2_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in2_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_2_flds_we),
    .q_o(data_in_2_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_2_we),
    .wd     (data_in_2_wd),

    // from internal hardware
    .de     (hw2reg.data_in[2].de),
    .d      (hw2reg.data_in[2].d),

    // to internal hardware
    .qe     (data_in_2_flds_we[0]),
    .q      (reg2hw.data_in[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_2_qs)
  );
  assign reg2hw.data_in[2].qe = data_in_2_qe;


  // Subregister 3 of Multireg data_in
  // R[data_in_3]: V(False)
  logic data_in_3_qe;
  logic [0:0] data_in_3_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in3_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_3_flds_we),
    .q_o(data_in_3_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_3_we),
    .wd     (data_in_3_wd),

    // from internal hardware
    .de     (hw2reg.data_in[3].de),
    .d      (hw2reg.data_in[3].d),

    // to internal hardware
    .qe     (data_in_3_flds_we[0]),
    .q      (reg2hw.data_in[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_3_qs)
  );
  assign reg2hw.data_in[3].qe = data_in_3_qe;


  // Subregister 0 of Multireg result_out
  // R[result_out_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[0].de),
    .d      (hw2reg.result_out[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_0_qs)
  );


  // Subregister 1 of Multireg result_out
  // R[result_out_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[1].de),
    .d      (hw2reg.result_out[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_1_qs)
  );


  // Subregister 2 of Multireg result_out
  // R[result_out_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[2].de),
    .d      (hw2reg.result_out[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_2_qs)
  );


  // Subregister 3 of Multireg result_out
  // R[result_out_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_result_out_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.result_out[3].de),
    .d      (hw2reg.result_out[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.result_out[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (result_out_3_qs)
  );



  logic [13:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == SM4_CTRL_SIGNALS_OFFSET);
    addr_hit[ 1] = (reg_addr == SM4_STATE_SIGNALS_OFFSET);
    addr_hit[ 2] = (reg_addr == SM4_KEY_0_OFFSET);
    addr_hit[ 3] = (reg_addr == SM4_KEY_1_OFFSET);
    addr_hit[ 4] = (reg_addr == SM4_KEY_2_OFFSET);
    addr_hit[ 5] = (reg_addr == SM4_KEY_3_OFFSET);
    addr_hit[ 6] = (reg_addr == SM4_DATA_IN_0_OFFSET);
    addr_hit[ 7] = (reg_addr == SM4_DATA_IN_1_OFFSET);
    addr_hit[ 8] = (reg_addr == SM4_DATA_IN_2_OFFSET);
    addr_hit[ 9] = (reg_addr == SM4_DATA_IN_3_OFFSET);
    addr_hit[10] = (reg_addr == SM4_RESULT_OUT_0_OFFSET);
    addr_hit[11] = (reg_addr == SM4_RESULT_OUT_1_OFFSET);
    addr_hit[12] = (reg_addr == SM4_RESULT_OUT_2_OFFSET);
    addr_hit[13] = (reg_addr == SM4_RESULT_OUT_3_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(SM4_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(SM4_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(SM4_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(SM4_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(SM4_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(SM4_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(SM4_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(SM4_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(SM4_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(SM4_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(SM4_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(SM4_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(SM4_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(SM4_PERMIT[13] & ~reg_be)))));
  end

  // Generate write-enables
  assign ctrl_signals_we = addr_hit[0] & reg_we & !reg_error;

  assign ctrl_signals_sm4_enable_in_wd = reg_wdata[0];

  assign ctrl_signals_encdec_sel_in_wd = reg_wdata[1];

  assign ctrl_signals_enable_key_exp_in_wd = reg_wdata[2];

  assign ctrl_signals_user_key_valid_in_wd = reg_wdata[3];

  assign ctrl_signals_encdec_enable_in_wd = reg_wdata[4];

  assign ctrl_signals_valid_in_wd = reg_wdata[5];
  assign key_0_we = addr_hit[2] & reg_we & !reg_error;

  assign key_0_wd = reg_wdata[31:0];
  assign key_1_we = addr_hit[3] & reg_we & !reg_error;

  assign key_1_wd = reg_wdata[31:0];
  assign key_2_we = addr_hit[4] & reg_we & !reg_error;

  assign key_2_wd = reg_wdata[31:0];
  assign key_3_we = addr_hit[5] & reg_we & !reg_error;

  assign key_3_wd = reg_wdata[31:0];
  assign data_in_0_we = addr_hit[6] & reg_we & !reg_error;

  assign data_in_0_wd = reg_wdata[31:0];
  assign data_in_1_we = addr_hit[7] & reg_we & !reg_error;

  assign data_in_1_wd = reg_wdata[31:0];
  assign data_in_2_we = addr_hit[8] & reg_we & !reg_error;

  assign data_in_2_wd = reg_wdata[31:0];
  assign data_in_3_we = addr_hit[9] & reg_we & !reg_error;

  assign data_in_3_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = ctrl_signals_we;
    reg_we_check[1] = 1'b0;
    reg_we_check[2] = key_0_we;
    reg_we_check[3] = key_1_we;
    reg_we_check[4] = key_2_we;
    reg_we_check[5] = key_3_we;
    reg_we_check[6] = data_in_0_we;
    reg_we_check[7] = data_in_1_we;
    reg_we_check[8] = data_in_2_we;
    reg_we_check[9] = data_in_3_we;
    reg_we_check[10] = 1'b0;
    reg_we_check[11] = 1'b0;
    reg_we_check[12] = 1'b0;
    reg_we_check[13] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = ctrl_signals_sm4_enable_in_qs;
        reg_rdata_next[1] = ctrl_signals_encdec_sel_in_qs;
        reg_rdata_next[2] = ctrl_signals_enable_key_exp_in_qs;
        reg_rdata_next[3] = ctrl_signals_user_key_valid_in_qs;
        reg_rdata_next[4] = ctrl_signals_encdec_enable_in_qs;
        reg_rdata_next[5] = ctrl_signals_valid_in_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = state_signals_key_exp_ready_out_qs;
        reg_rdata_next[1] = state_signals_valid_out_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = key_0_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = key_1_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = key_2_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = key_3_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = data_in_0_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = data_in_1_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = data_in_2_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = data_in_3_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = result_out_0_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = result_out_1_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = result_out_2_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = result_out_3_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


`include "prim_assert.sv"

module sm4
  import sm4_reg_pkg::*;
(
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  // Bus interface
  input  tlul_pkg::tl_h2d_t                         tl_i,
  output tlul_pkg::tl_d2h_t                         tl_o
);

  sm4_reg2hw_t               reg2hw;
  sm4_hw2reg_t               hw2reg;
  //wire                       ready_out;

sm4_reg_top  u_sm4_reg_top (
    .clk_i                             ( clk_i        ),
    .rst_ni                            ( rst_ni       ),
    .tl_i                              ( tl_i         ),
    .hw2reg                            ( hw2reg       ),
    .devmode_i                         ( 1'b1         ),

    .tl_o                              ( tl_o         ),
    .reg2hw                            ( reg2hw       ),
    .intg_err_o                        (   )
);

/*assign hw2reg.result_out[0].de={32(ready_out)};
assign hw2reg.result_out[1].de={32(ready_out)};
assign hw2reg.result_out[2].de={32(ready_out)};
assign hw2reg.result_out[3].de={32(ready_out)};
*/

assign hw2reg.ctrl_signals.sm4_enable_in.de = 1'd0;
assign hw2reg.ctrl_signals.encdec_enable_in.de = 1'd0;
assign hw2reg.ctrl_signals.encdec_sel_in.de = 1'd0;
assign hw2reg.ctrl_signals.valid_in.de = 1'd0;
assign hw2reg.data_in[0].de = 1'd0;
assign hw2reg.data_in[1].de = 1'd0;
assign hw2reg.data_in[2].de = 1'd0;
assign hw2reg.data_in[3].de = 1'd0;
assign hw2reg.ctrl_signals.enable_key_exp_in.de = 1'd0;
assign hw2reg.ctrl_signals.user_key_valid_in.de = 1'd0;
assign hw2reg.key[0].de = 1'd0;
assign hw2reg.key[1].de = 1'd0;
assign hw2reg.key[2].de = 1'd0;
assign hw2reg.key[3].de = 1'd0;


sm4_top  u_sm4_top (
    .clk                     ( clk_i        ),
    .reset_n                 ( rst_ni       ),
    .sm4_enable_in           ( reg2hw.ctrl_signals.sm4_enable_in.q),
    .encdec_enable_in        ( reg2hw.ctrl_signals.encdec_enable_in.q ),
    .encdec_sel_in           ( reg2hw.ctrl_signals.encdec_sel_in.q ),
    .valid_in                ( reg2hw.ctrl_signals.valid_in.q ),
    .data_in                 ( {reg2hw.data_in[3].q,reg2hw.data_in[2].q,reg2hw.data_in[1].q,reg2hw.data_in[0].q}),
    .enable_key_exp_in       ( reg2hw.ctrl_signals.enable_key_exp_in.q  ),
    .user_key_valid_in       ( reg2hw.ctrl_signals.user_key_valid_in.q ),
    .user_key_in             ( {reg2hw.key[3].q,reg2hw.key[2].q,reg2hw.key[1].q,reg2hw.key[0].q} ),

    //.ready_out               ( ready_out ),
    .result_out              ( {hw2reg.result_out[3].d,hw2reg.result_out[2].d,hw2reg.result_out[1].d,hw2reg.result_out[0].d} ),
    .valid_out               ( hw2reg.state_signals.valid_out.d),
    .key_exp_ready_out       ( hw2reg.state_signals.key_exp_ready_out.d),
    .ready_out_de            ( {hw2reg.result_out[3].de,hw2reg.result_out[2].de,hw2reg.result_out[1].de,hw2reg.result_out[0].de }),
    .valid_out_de            (hw2reg.state_signals.valid_out.de)
);
    
endmodule

// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/10 12:06:49
// Design Name: 
// Module Name: sm4_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module sm4_top(
    clk		            ,
    reset_n	            ,
    sm4_enable_in       ,
    encdec_enable_in    ,
    encdec_sel_in       ,
    valid_in            ,
    data_in             ,
    enable_key_exp_in   ,
    user_key_valid_in   ,
    user_key_in         ,
    key_exp_ready_out   ,
    result_out          ,
    valid_out           ,
    ready_out_de        ,
    valid_out_de
);
    
    input			 clk		        ;
    input			 reset_n	        ;
    input            sm4_enable_in      ;
    input            encdec_enable_in   ;
    input            encdec_sel_in      ;
    input            valid_in           ;
    input   [127: 0] data_in            ;
    input            enable_key_exp_in  ;
    input            user_key_valid_in  ;
    input   [127: 0] user_key_in        ;
    output  [3: 0] ready_out_de       ;
    output           valid_out_de       ;
    output  [127: 0] result_out         ;
    
    output           valid_out          ;
    output           key_exp_ready_out  ;
    wire             ready_out          ;
    wire    [31 : 0] rk_00              ;
    wire    [31 : 0] rk_01              ;
    wire    [31 : 0] rk_02              ;
    wire    [31 : 0] rk_03              ;
    wire    [31 : 0] rk_04              ;
    wire    [31 : 0] rk_05              ;
    wire    [31 : 0] rk_06              ;
    wire    [31 : 0] rk_07              ;
    wire    [31 : 0] rk_08              ;
    wire    [31 : 0] rk_09              ;
    wire    [31 : 0] rk_10              ;
    wire    [31 : 0] rk_11              ;
    wire    [31 : 0] rk_12              ;
    wire    [31 : 0] rk_13              ;
    wire    [31 : 0] rk_14              ;
    wire    [31 : 0] rk_15              ;
    wire    [31 : 0] rk_16              ;
    wire    [31 : 0] rk_17              ;
    wire    [31 : 0] rk_18              ;
    wire    [31 : 0] rk_19              ;
    wire    [31 : 0] rk_20              ;
    wire    [31 : 0] rk_21              ;
    wire    [31 : 0] rk_22              ;
    wire    [31 : 0] rk_23              ;
    wire    [31 : 0] rk_24              ;
    wire    [31 : 0] rk_25              ;
    wire    [31 : 0] rk_26              ;
    wire    [31 : 0] rk_27              ;
    wire    [31 : 0] rk_28              ;
    wire    [31 : 0] rk_29              ;
    wire    [31 : 0] rk_30              ;
    wire    [31 : 0] rk_31              ;
    
    ready_valid u_ready_valid(
      .clk              (clk              ),
      .ready_out        (ready_out        ),
      .encdec_enable_in (encdec_enable_in ),
      .valid_out        (valid_out        )
    );
  
    sm4_encdec u_encdec (
        .clk                    (clk                 ),
        .reset_n                (reset_n             ),
        .sm4_enable_in          (sm4_enable_in       ),
        .encdec_enable_in       (encdec_enable_in    ),
        .key_exp_ready_in       (key_exp_ready_out   ),
        .valid_in               (valid_in            ),
        .data_in                (data_in             ),
        .rk_00_in               (rk_00               ),
        .rk_01_in               (rk_01               ),
        .rk_02_in               (rk_02               ),
        .rk_03_in               (rk_03               ),
        .rk_04_in               (rk_04               ),
        .rk_05_in               (rk_05               ),
        .rk_06_in               (rk_06               ),
        .rk_07_in               (rk_07               ),
        .rk_08_in               (rk_08               ),
        .rk_09_in               (rk_09               ),
        .rk_10_in               (rk_10               ),
        .rk_11_in               (rk_11               ),
        .rk_12_in               (rk_12               ),
        .rk_13_in               (rk_13               ),
        .rk_14_in               (rk_14               ),
        .rk_15_in               (rk_15               ),
        .rk_16_in               (rk_16               ),
        .rk_17_in               (rk_17               ),
        .rk_18_in               (rk_18               ),
        .rk_19_in               (rk_19               ),
        .rk_20_in               (rk_20               ),
        .rk_21_in               (rk_21               ),
        .rk_22_in               (rk_22               ),
        .rk_23_in               (rk_23               ),
        .rk_24_in               (rk_24               ),
        .rk_25_in               (rk_25               ),
        .rk_26_in               (rk_26               ),
        .rk_27_in               (rk_27               ),
        .rk_28_in               (rk_28               ),
        .rk_29_in               (rk_29               ),
        .rk_30_in               (rk_30               ),
        .rk_31_in               (rk_31               ),
        .ready_out              (ready_out           ),
        .result_out             (result_out          )
    );
    
    assign ready_out_de = {4{ready_out}};
    assign valid_out_de=valid_out;

    key_expansion u_key
	(
        .clk					(clk					),
        .reset_n				(reset_n				),
        .sm4_enable_in		    (sm4_enable_in		    ),
        .encdec_sel_in		    (encdec_sel_in		    ),
        .enable_key_exp_in	    (enable_key_exp_in	    ),
        .user_key_in			(user_key_in			),
        .user_key_valid_in	    (user_key_valid_in	    ),
        .key_exp_finished_out   (key_exp_ready_out      ),
        .rk00_out			    (rk_00    			    ),
        .rk01_out			    (rk_01    			    ),
        .rk02_out			    (rk_02    			    ),
        .rk03_out			    (rk_03    			    ),
        .rk04_out			    (rk_04    			    ),
        .rk05_out			    (rk_05    			    ),
        .rk06_out			    (rk_06    			    ),
        .rk07_out			    (rk_07    			    ),
        .rk08_out			    (rk_08    			    ),
        .rk09_out			    (rk_09    			    ),
        .rk10_out			    (rk_10    			    ),
        .rk11_out			    (rk_11    			    ),
        .rk12_out			    (rk_12    			    ),
        .rk13_out			    (rk_13    			    ),
        .rk14_out			    (rk_14    			    ),
        .rk15_out			    (rk_15    			    ),
        .rk16_out			    (rk_16    			    ),
        .rk17_out			    (rk_17    			    ),
        .rk18_out			    (rk_18    			    ),
        .rk19_out			    (rk_19    			    ),
        .rk20_out			    (rk_20    			    ),
        .rk21_out			    (rk_21    			    ),
        .rk22_out			    (rk_22    			    ),
        .rk23_out			    (rk_23    			    ),
        .rk24_out			    (rk_24    			    ),
        .rk25_out			    (rk_25    			    ),
        .rk26_out			    (rk_26    			    ),
        .rk27_out			    (rk_27    			    ),
        .rk28_out			    (rk_28    			    ),
        .rk29_out			    (rk_29    			    ),
        .rk30_out			    (rk_30    			    ),
        .rk31_out			    (rk_31    			    )
    );
    
endmodule


// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/10 10:22:18
// Design Name: 
// Module Name: transform_for_encdec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module transform_for_encdec(
		data_in,
		result_out
	);
input	[31:0]	data_in;
output	[31:0]	result_out;			

wire	[7:0]	byte_0;
wire	[7:0]	byte_1;
wire	[7:0]	byte_2;
wire	[7:0]	byte_3;
wire	[7:0]	byte_0_replaced;
wire	[7:0]	byte_1_replaced;
wire	[7:0]	byte_2_replaced;
wire	[7:0]	byte_3_replaced;
wire	[31:0]	word_replaced;
wire	[31:0]	data_after_linear;
wire	[31:0]	data_after_linear_key;

assign	{ byte_0, byte_1, byte_2, byte_3 } = data_in;
assign	word_replaced = {byte_0_replaced, byte_1_replaced, byte_2_replaced,byte_3_replaced};

sbox_replace	u_0
	(
		.data_in(byte_0),
		.result_out(byte_0_replaced)														
	);
	
sbox_replace	u_1
	(
		.data_in(byte_1),
		.result_out(byte_1_replaced)														
	);
	
sbox_replace	u_2
	(
		.data_in(byte_2),
		.result_out(byte_2_replaced)														
	);
	
sbox_replace	u_3
	(
		.data_in(byte_3),
		.result_out(byte_3_replaced)														
	);	

assign	result_out = ( 	 (word_replaced ^ {word_replaced[29:0], word_replaced[31:30]}) 
                       ^ ({word_replaced[21:0], word_replaced[31:22]} ^ {word_replaced[13:0], word_replaced[31:14]})) 
				   ^ {word_replaced[7:0], word_replaced[31:8]};
													
endmodule		

// `timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Raymond Rui Chen, raymond.rui.chen@qq.com
// 
// Create Date: 2018/03/09 21:16:22
// Design Name: 
// Module Name: transform_for_key_exp
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module transform_for_key_exp
	(
		data_in,
		data_after_linear_key_out
	);
input	[31 : 0]	data_in;

output	[31 : 0]	data_after_linear_key_out; 	

wire	[7:0]	byte_0;
wire	[7:0]	byte_1;
wire	[7:0]	byte_2;
wire	[7:0]	byte_3;
wire	[7:0]	byte_0_replaced;
wire	[7:0]	byte_1_replaced;
wire	[7:0]	byte_2_replaced;
wire	[7:0]	byte_3_replaced;
wire	[31:0]	word_replaced;

assign	{	byte_0,
			byte_1,
			byte_2,
			byte_3}	=	data_in;

assign	word_replaced	=	{	byte_0_replaced,
								byte_1_replaced,
								byte_2_replaced,
								byte_3_replaced};

sbox_replace u_0
	(
		.data_in(byte_0),
		.result_out(byte_0_replaced)														
	);

sbox_replace	u_1
	(
		.data_in(byte_1),
		.result_out(byte_1_replaced)														
	);
	
sbox_replace	u_2
	(
		.data_in(byte_2),
		.result_out(byte_2_replaced)														
	);
	
sbox_replace	u_3
	(
		.data_in(byte_3),
		.result_out(byte_3_replaced)														
	);																																				

assign	data_after_linear_key_out	= (word_replaced ^ {word_replaced[18:0], word_replaced[31:19]}) 
					^ {word_replaced[8:0], word_replaced[31:9]};

endmodule											
																								


// -------------------------------------------------------------------------
//Berlekamp circuit for Reed-Solomon decoder
//Copyright (C) Tue Apr  2 17:07:10 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module rsdec_berl (lambda_out, omega_out, syndrome0, syndrome1, syndrome2, syndrome3, syndrome4, syndrome5, syndrome6, syndrome7, syndrome8, syndrome9, syndrome10, syndrome11, syndrome12, syndrome13, syndrome14, syndrome15, syndrome16, syndrome17, syndrome18, syndrome19, syndrome20, syndrome21, syndrome22, syndrome23, syndrome24, syndrome25, syndrome26, syndrome27, syndrome28, syndrome29, syndrome30, syndrome31, 
		D, DI, count, phase0, phase32, enable, clk, clrn);
	input clk, clrn, enable, phase0, phase32;
	input [7:0] syndrome0;
	input [7:0] syndrome1;
	input [7:0] syndrome2;
	input [7:0] syndrome3;
	input [7:0] syndrome4;
	input [7:0] syndrome5;
	input [7:0] syndrome6;
	input [7:0] syndrome7;
	input [7:0] syndrome8;
	input [7:0] syndrome9;
	input [7:0] syndrome10;
	input [7:0] syndrome11;
	input [7:0] syndrome12;
	input [7:0] syndrome13;
	input [7:0] syndrome14;
	input [7:0] syndrome15;
	input [7:0] syndrome16;
	input [7:0] syndrome17;
	input [7:0] syndrome18;
	input [7:0] syndrome19;
	input [7:0] syndrome20;
	input [7:0] syndrome21;
	input [7:0] syndrome22;
	input [7:0] syndrome23;
	input [7:0] syndrome24;
	input [7:0] syndrome25;
	input [7:0] syndrome26;
	input [7:0] syndrome27;
	input [7:0] syndrome28;
	input [7:0] syndrome29;
	input [7:0] syndrome30;
	input [7:0] syndrome31;
	input [7:0] DI;
	input [5:0] count;
	output [7:0] lambda_out;
	output [7:0] omega_out;
	reg [7:0] lambda_out;
	reg [7:0] omega_out;
	output [7:0] D;
	reg [7:0] D;

	integer j;
	reg init, delta;
	reg [4:0] L;
	reg [7:0] lambda[31:0];
	reg [7:0] omega[31:0];
	reg [7:0] A[30:0];
	reg [7:0] B[30:0];
	wire [7:0] tmp0;
	wire [7:0] tmp1;
	wire [7:0] tmp2;
	wire [7:0] tmp3;
	wire [7:0] tmp4;
	wire [7:0] tmp5;
	wire [7:0] tmp6;
	wire [7:0] tmp7;
	wire [7:0] tmp8;
	wire [7:0] tmp9;
	wire [7:0] tmp10;
	wire [7:0] tmp11;
	wire [7:0] tmp12;
	wire [7:0] tmp13;
	wire [7:0] tmp14;
	wire [7:0] tmp15;
	wire [7:0] tmp16;
	wire [7:0] tmp17;
	wire [7:0] tmp18;
	wire [7:0] tmp19;
	wire [7:0] tmp20;
	wire [7:0] tmp21;
	wire [7:0] tmp22;
	wire [7:0] tmp23;
	wire [7:0] tmp24;
	wire [7:0] tmp25;
	wire [7:0] tmp26;
	wire [7:0] tmp27;
	wire [7:0] tmp28;
	wire [7:0] tmp29;
	wire [7:0] tmp30;
	wire [7:0] tmp31;

	always @ (tmp1) lambda_out = tmp1;
	always @ (tmp3) omega_out = tmp3;

	always @ (L or D or count)
		// delta = (D != 0 && 2*L <= i);
		if (D != 0 && count >= {L, 1'b0}) delta = 1;
		else delta = 0;

	rsdec_berl_multiply x0 (tmp0, B[30], D, lambda[0], syndrome0, phase0);
	rsdec_berl_multiply x1 (tmp1, lambda[31], DI, lambda[1], syndrome1, phase0);
	rsdec_berl_multiply x2 (tmp2, A[30], D, lambda[2], syndrome2, phase0);
	rsdec_berl_multiply x3 (tmp3, omega[31], DI, lambda[3], syndrome3, phase0);
	multiply x4 (tmp4, lambda[4], syndrome4);
	multiply x5 (tmp5, lambda[5], syndrome5);
	multiply x6 (tmp6, lambda[6], syndrome6);
	multiply x7 (tmp7, lambda[7], syndrome7);
	multiply x8 (tmp8, lambda[8], syndrome8);
	multiply x9 (tmp9, lambda[9], syndrome9);
	multiply x10 (tmp10, lambda[10], syndrome10);
	multiply x11 (tmp11, lambda[11], syndrome11);
	multiply x12 (tmp12, lambda[12], syndrome12);
	multiply x13 (tmp13, lambda[13], syndrome13);
	multiply x14 (tmp14, lambda[14], syndrome14);
	multiply x15 (tmp15, lambda[15], syndrome15);
	multiply x16 (tmp16, lambda[16], syndrome16);
	multiply x17 (tmp17, lambda[17], syndrome17);
	multiply x18 (tmp18, lambda[18], syndrome18);
	multiply x19 (tmp19, lambda[19], syndrome19);
	multiply x20 (tmp20, lambda[20], syndrome20);
	multiply x21 (tmp21, lambda[21], syndrome21);
	multiply x22 (tmp22, lambda[22], syndrome22);
	multiply x23 (tmp23, lambda[23], syndrome23);
	multiply x24 (tmp24, lambda[24], syndrome24);
	multiply x25 (tmp25, lambda[25], syndrome25);
	multiply x26 (tmp26, lambda[26], syndrome26);
	multiply x27 (tmp27, lambda[27], syndrome27);
	multiply x28 (tmp28, lambda[28], syndrome28);
	multiply x29 (tmp29, lambda[29], syndrome29);
	multiply x30 (tmp30, lambda[30], syndrome30);
	multiply x31 (tmp31, lambda[31], syndrome31);

	always @ (posedge clk or negedge clrn)
	begin
		// for (j = t-1; j >=0; j--)
		//	if (j != 0) lambda[j] += D * B[j-1];
		if (~clrn)
		begin
			for (j = 0; j < 32; j = j + 1) lambda[j] <= 0;
			for (j = 0; j < 31; j = j + 1) B[j] <= 0;
			for (j = 0; j < 32; j = j + 1) omega[j] <= 0;
			for (j = 0; j < 31; j = j + 1) A[j] <= 0;
			L <= 0;
			D <= 0;
		end
		else if (~enable)
		begin
			lambda[0] <= 1;
			for (j = 1; j < 32; j = j +1) lambda[j] <= 0;
			B[0] <= 1;
			for (j = 1; j < 31; j = j +1) B[j] <= 0;
			omega[0] <= 1;
			for (j = 1; j < 32; j = j +1) omega[j] <= 0;
			for (j = 0; j < 31; j = j + 1) A[j] <= 0;
			L <= 0;
			D <= 0;
		end
		else
		begin
			if (~phase0)
			begin
				if (~phase32) lambda[0] <= lambda[31] ^ tmp0;
				else lambda[0] <= lambda[31];
				for (j = 1; j < 32; j = j + 1)
					lambda[j] <= lambda[j-1];
			end

		// for (j = t-1; j >=0; j--)
		//	if (delta) B[j] = lambda[j] *DI;
		//	else if (j != 0) B[j] = B[j-1];
		//	else B[j] = 0;
			if (~phase0)
			begin
				if (delta)	B[0] <= tmp1;
				else if (~phase32) B[0] <= B[30];
				else B[0] <= 0;
				for (j = 1; j < 31; j = j + 1)
					B[j] <= B[j-1];
			end

		// for (j = t-1; j >=0; j--)
		//	if (j != 0) omega[j] += D * A[j-1];
			if (~phase0)
			begin
				if (~phase32) omega[0] <= omega[31] ^ tmp2;
				else omega[0] <= omega[31];
				for (j = 1; j < 32; j = j + 1)
					omega[j] <= omega[j-1];
			end

		// for (j = t-1; j >=0; j--)
		//	if (delta) A[j] = omega[j] *DI;
		//	else if (j != 0) A[j] = A[j-1];
		//	else A[j] = 0;
			if (~phase0)
			begin
				if (delta)	A[0] <= tmp3;
				else if (~phase32) A[0] <= A[30];
				else A[0] <= 0;
				for (j = 1; j < 31; j = j + 1)
					A[j] <= A[j-1];
			end

		// if (delta) L = i - L + 1;
			if ((phase0 & delta) && (count != -1)) L <= count - L + 1;

		//for (D = j = 0; j < t; j = j + 1)
		//	D += lambda[j] * syndrome[t-j-1];
			if (phase0)
				D <= tmp0 ^ tmp1 ^ tmp2 ^ tmp3 ^ tmp4 ^ tmp5 ^ tmp6 ^ tmp7 ^ tmp8 ^ tmp9 ^ tmp10 ^ tmp11 ^ tmp12 ^ tmp13 ^ tmp14 ^ tmp15 ^ tmp16 ^ tmp17 ^ tmp18 ^ tmp19 ^ tmp20 ^ tmp21 ^ tmp22 ^ tmp23 ^ tmp24 ^ tmp25 ^ tmp26 ^ tmp27 ^ tmp28 ^ tmp29 ^ tmp30 ^ tmp31;

		end
	end

endmodule


module rsdec_berl_multiply (y, a, b, c, d, e);
	input [7:0] a, b, c, d;
	input e;
	output [7:0] y;
	wire [7:0] y;
	reg [7:0] p, q;

	always @ (a or c or e)
		if (e) p = c;
		else p = a;
	always @ (b or d or e)
		if (e) q = d;
		else q = b;

	multiply x0 (y, p, q);

endmodule

module multiply (y, a, b);
	input [7:0] a, b;
	output [7:0] y;
	reg [7:0] y;
	always @ (a or b)
	begin
		y[0] = (a[0] & b[0]) ^ (a[1] & b[7]) ^ (a[2] & b[6]) ^ (a[2] & b[7]) ^ (a[3] & b[5]) ^ (a[3] & b[6]) ^ (a[3] & b[7]) ^ (a[4] & b[4]) ^ (a[4] & b[5]) ^ (a[4] & b[6]) ^ (a[4] & b[7]) ^ (a[5] & b[3]) ^ (a[5] & b[4]) ^ (a[5] & b[5]) ^ (a[5] & b[6]) ^ (a[5] & b[7]) ^ (a[6] & b[2]) ^ (a[6] & b[3]) ^ (a[6] & b[4]) ^ (a[6] & b[5]) ^ (a[6] & b[6]) ^ (a[6] & b[7]) ^ (a[7] & b[1]) ^ (a[7] & b[2]) ^ (a[7] & b[3]) ^ (a[7] & b[4]) ^ (a[7] & b[5]) ^ (a[7] & b[6]);
		y[1] = (a[0] & b[1]) ^ (a[1] & b[0]) ^ (a[1] & b[7]) ^ (a[2] & b[6]) ^ (a[3] & b[5]) ^ (a[4] & b[4]) ^ (a[5] & b[3]) ^ (a[6] & b[2]) ^ (a[7] & b[1]) ^ (a[7] & b[7]);
		y[2] = (a[0] & b[2]) ^ (a[1] & b[1]) ^ (a[1] & b[7]) ^ (a[2] & b[0]) ^ (a[2] & b[6]) ^ (a[3] & b[5]) ^ (a[3] & b[7]) ^ (a[4] & b[4]) ^ (a[4] & b[6]) ^ (a[4] & b[7]) ^ (a[5] & b[3]) ^ (a[5] & b[5]) ^ (a[5] & b[6]) ^ (a[5] & b[7]) ^ (a[6] & b[2]) ^ (a[6] & b[4]) ^ (a[6] & b[5]) ^ (a[6] & b[6]) ^ (a[6] & b[7]) ^ (a[7] & b[1]) ^ (a[7] & b[3]) ^ (a[7] & b[4]) ^ (a[7] & b[5]) ^ (a[7] & b[6]);
		y[3] = (a[0] & b[3]) ^ (a[1] & b[2]) ^ (a[2] & b[1]) ^ (a[2] & b[7]) ^ (a[3] & b[0]) ^ (a[3] & b[6]) ^ (a[4] & b[5]) ^ (a[4] & b[7]) ^ (a[5] & b[4]) ^ (a[5] & b[6]) ^ (a[5] & b[7]) ^ (a[6] & b[3]) ^ (a[6] & b[5]) ^ (a[6] & b[6]) ^ (a[6] & b[7]) ^ (a[7] & b[2]) ^ (a[7] & b[4]) ^ (a[7] & b[5]) ^ (a[7] & b[6]) ^ (a[7] & b[7]);
		y[4] = (a[0] & b[4]) ^ (a[1] & b[3]) ^ (a[2] & b[2]) ^ (a[3] & b[1]) ^ (a[3] & b[7]) ^ (a[4] & b[0]) ^ (a[4] & b[6]) ^ (a[5] & b[5]) ^ (a[5] & b[7]) ^ (a[6] & b[4]) ^ (a[6] & b[6]) ^ (a[6] & b[7]) ^ (a[7] & b[3]) ^ (a[7] & b[5]) ^ (a[7] & b[6]) ^ (a[7] & b[7]);
		y[5] = (a[0] & b[5]) ^ (a[1] & b[4]) ^ (a[2] & b[3]) ^ (a[3] & b[2]) ^ (a[4] & b[1]) ^ (a[4] & b[7]) ^ (a[5] & b[0]) ^ (a[5] & b[6]) ^ (a[6] & b[5]) ^ (a[6] & b[7]) ^ (a[7] & b[4]) ^ (a[7] & b[6]) ^ (a[7] & b[7]);
		y[6] = (a[0] & b[6]) ^ (a[1] & b[5]) ^ (a[2] & b[4]) ^ (a[3] & b[3]) ^ (a[4] & b[2]) ^ (a[5] & b[1]) ^ (a[5] & b[7]) ^ (a[6] & b[0]) ^ (a[6] & b[6]) ^ (a[7] & b[5]) ^ (a[7] & b[7]);
		y[7] = (a[0] & b[7]) ^ (a[1] & b[6]) ^ (a[1] & b[7]) ^ (a[2] & b[5]) ^ (a[2] & b[6]) ^ (a[2] & b[7]) ^ (a[3] & b[4]) ^ (a[3] & b[5]) ^ (a[3] & b[6]) ^ (a[3] & b[7]) ^ (a[4] & b[3]) ^ (a[4] & b[4]) ^ (a[4] & b[5]) ^ (a[4] & b[6]) ^ (a[4] & b[7]) ^ (a[5] & b[2]) ^ (a[5] & b[3]) ^ (a[5] & b[4]) ^ (a[5] & b[5]) ^ (a[5] & b[6]) ^ (a[5] & b[7]) ^ (a[6] & b[1]) ^ (a[6] & b[2]) ^ (a[6] & b[3]) ^ (a[6] & b[4]) ^ (a[6] & b[5]) ^ (a[6] & b[6]) ^ (a[7] & b[0]) ^ (a[7] & b[1]) ^ (a[7] & b[2]) ^ (a[7] & b[3]) ^ (a[7] & b[4]) ^ (a[7] & b[5]);
	end
endmodule



// -------------------------------------------------------------------------
//Chien-Forney search circuit for Reed-Solomon decoder
//Copyright (C) Tue Apr  2 17:07:16 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module rsdec_chien_scale0 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0];
		y[1] = x[1];
		y[2] = x[2];
		y[3] = x[3];
		y[4] = x[4];
		y[5] = x[5];
		y[6] = x[6];
		y[7] = x[7];
	end
endmodule

module rsdec_chien_scale1 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[7];
		y[1] = x[0] ^ x[7];
		y[2] = x[1] ^ x[7];
		y[3] = x[2];
		y[4] = x[3];
		y[5] = x[4];
		y[6] = x[5];
		y[7] = x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale2 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[6] ^ x[7];
		y[1] = x[6];
		y[2] = x[0] ^ x[6];
		y[3] = x[1] ^ x[7];
		y[4] = x[2];
		y[5] = x[3];
		y[6] = x[4];
		y[7] = x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale3 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[5] ^ x[6] ^ x[7];
		y[1] = x[5];
		y[2] = x[5] ^ x[7];
		y[3] = x[0] ^ x[6];
		y[4] = x[1] ^ x[7];
		y[5] = x[2];
		y[6] = x[3];
		y[7] = x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale4 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[4];
		y[2] = x[4] ^ x[6] ^ x[7];
		y[3] = x[5] ^ x[7];
		y[4] = x[0] ^ x[6];
		y[5] = x[1] ^ x[7];
		y[6] = x[2];
		y[7] = x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale5 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[3];
		y[2] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[4] ^ x[6] ^ x[7];
		y[4] = x[5] ^ x[7];
		y[5] = x[0] ^ x[6];
		y[6] = x[1] ^ x[7];
		y[7] = x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale6 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[2];
		y[2] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[4] ^ x[6] ^ x[7];
		y[5] = x[5] ^ x[7];
		y[6] = x[0] ^ x[6];
		y[7] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_chien_scale7 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[1] = x[1] ^ x[7];
		y[2] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[4] ^ x[6] ^ x[7];
		y[6] = x[5] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
	end
endmodule

module rsdec_chien_scale8 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[1] = x[0] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[4] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
	end
endmodule

module rsdec_chien_scale9 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
		y[1] = x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6];
	end
endmodule

module rsdec_chien_scale10 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6];
		y[1] = x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_chien_scale11 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[7];
		y[1] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[6] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[4] ^ x[6];
	end
endmodule

module rsdec_chien_scale12 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[4] ^ x[6];
		y[1] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[0] ^ x[3] ^ x[5];
	end
endmodule

module rsdec_chien_scale13 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[5];
		y[1] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[4] ^ x[7];
	end
endmodule

module rsdec_chien_scale14 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[2] ^ x[4] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[6];
	end
endmodule

module rsdec_chien_scale15 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[6];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_chien_scale16 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[1] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale17 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[4] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[3] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_chien_scale18 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[5] ^ x[6];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[4] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_chien_scale19 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[2] ^ x[4] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[4] ^ x[6];
	end
endmodule

module rsdec_chien_scale20 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[4] ^ x[6];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[6] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_chien_scale21 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[7] = x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale22 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[5];
		y[3] = x[0] ^ x[1] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale23 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[2] = x[4] ^ x[7];
		y[3] = x[0] ^ x[5];
		y[4] = x[0] ^ x[1] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[7] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale24 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[2] = x[3] ^ x[6] ^ x[7];
		y[3] = x[4] ^ x[7];
		y[4] = x[0] ^ x[5];
		y[5] = x[0] ^ x[1] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien_scale25 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[2] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[3] ^ x[6] ^ x[7];
		y[4] = x[4] ^ x[7];
		y[5] = x[0] ^ x[5];
		y[6] = x[0] ^ x[1] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_chien_scale26 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[2] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[3] ^ x[6] ^ x[7];
		y[5] = x[4] ^ x[7];
		y[6] = x[0] ^ x[5];
		y[7] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
	end
endmodule

module rsdec_chien_scale27 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[1] = x[0] ^ x[1] ^ x[6];
		y[2] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[3] ^ x[6] ^ x[7];
		y[6] = x[4] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4];
	end
endmodule

module rsdec_chien_scale28 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4];
		y[1] = x[0] ^ x[5];
		y[2] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[3] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[3] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[7];
	end
endmodule

module rsdec_chien_scale29 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[7];
		y[1] = x[4] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[3] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[4] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[6];
	end
endmodule

module rsdec_chien_scale30 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[6];
		y[1] = x[3] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[4] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[5] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[6] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_chien_scale31 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[5] ^ x[7];
		y[1] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[5] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[6] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[0] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_chien (error, alpha, lambda, omega, even, D, search, load, shorten, clk, clrn);
	input clk, clrn, load, search, shorten;
	input [7:0] D;
	input [7:0] lambda;
	input [7:0] omega;
	output [7:0] even, error;
	output [7:0] alpha;
	reg [7:0] even, error;
	reg [7:0] alpha;

	wire [7:0] scale0;
	wire [7:0] scale1;
	wire [7:0] scale2;
	wire [7:0] scale3;
	wire [7:0] scale4;
	wire [7:0] scale5;
	wire [7:0] scale6;
	wire [7:0] scale7;
	wire [7:0] scale8;
	wire [7:0] scale9;
	wire [7:0] scale10;
	wire [7:0] scale11;
	wire [7:0] scale12;
	wire [7:0] scale13;
	wire [7:0] scale14;
	wire [7:0] scale15;
	wire [7:0] scale16;
	wire [7:0] scale17;
	wire [7:0] scale18;
	wire [7:0] scale19;
	wire [7:0] scale20;
	wire [7:0] scale21;
	wire [7:0] scale22;
	wire [7:0] scale23;
	wire [7:0] scale24;
	wire [7:0] scale25;
	wire [7:0] scale26;
	wire [7:0] scale27;
	wire [7:0] scale28;
	wire [7:0] scale29;
	wire [7:0] scale30;
	wire [7:0] scale31;
	wire [7:0] scale32;
	wire [7:0] scale33;
	wire [7:0] scale34;
	wire [7:0] scale35;
	wire [7:0] scale36;
	wire [7:0] scale37;
	wire [7:0] scale38;
	wire [7:0] scale39;
	wire [7:0] scale40;
	wire [7:0] scale41;
	wire [7:0] scale42;
	wire [7:0] scale43;
	wire [7:0] scale44;
	wire [7:0] scale45;
	wire [7:0] scale46;
	wire [7:0] scale47;
	wire [7:0] scale48;
	wire [7:0] scale49;
	wire [7:0] scale50;
	wire [7:0] scale51;
	wire [7:0] scale52;
	wire [7:0] scale53;
	wire [7:0] scale54;
	wire [7:0] scale55;
	wire [7:0] scale56;
	wire [7:0] scale57;
	wire [7:0] scale58;
	wire [7:0] scale59;
	wire [7:0] scale60;
	wire [7:0] scale61;
	wire [7:0] scale62;
	wire [7:0] scale63;
	reg [7:0] data0;
	reg [7:0] data1;
	reg [7:0] data2;
	reg [7:0] data3;
	reg [7:0] data4;
	reg [7:0] data5;
	reg [7:0] data6;
	reg [7:0] data7;
	reg [7:0] data8;
	reg [7:0] data9;
	reg [7:0] data10;
	reg [7:0] data11;
	reg [7:0] data12;
	reg [7:0] data13;
	reg [7:0] data14;
	reg [7:0] data15;
	reg [7:0] data16;
	reg [7:0] data17;
	reg [7:0] data18;
	reg [7:0] data19;
	reg [7:0] data20;
	reg [7:0] data21;
	reg [7:0] data22;
	reg [7:0] data23;
	reg [7:0] data24;
	reg [7:0] data25;
	reg [7:0] data26;
	reg [7:0] data27;
	reg [7:0] data28;
	reg [7:0] data29;
	reg [7:0] data30;
	reg [7:0] data31;
	reg [7:0] a0;
	reg [7:0] a1;
	reg [7:0] a2;
	reg [7:0] a3;
	reg [7:0] a4;
	reg [7:0] a5;
	reg [7:0] a6;
	reg [7:0] a7;
	reg [7:0] a8;
	reg [7:0] a9;
	reg [7:0] a10;
	reg [7:0] a11;
	reg [7:0] a12;
	reg [7:0] a13;
	reg [7:0] a14;
	reg [7:0] a15;
	reg [7:0] a16;
	reg [7:0] a17;
	reg [7:0] a18;
	reg [7:0] a19;
	reg [7:0] a20;
	reg [7:0] a21;
	reg [7:0] a22;
	reg [7:0] a23;
	reg [7:0] a24;
	reg [7:0] a25;
	reg [7:0] a26;
	reg [7:0] a27;
	reg [7:0] a28;
	reg [7:0] a29;
	reg [7:0] a30;
	reg [7:0] a31;
	reg [7:0] l0;
	reg [7:0] l1;
	reg [7:0] l2;
	reg [7:0] l3;
	reg [7:0] l4;
	reg [7:0] l5;
	reg [7:0] l6;
	reg [7:0] l7;
	reg [7:0] l8;
	reg [7:0] l9;
	reg [7:0] l10;
	reg [7:0] l11;
	reg [7:0] l12;
	reg [7:0] l13;
	reg [7:0] l14;
	reg [7:0] l15;
	reg [7:0] l16;
	reg [7:0] l17;
	reg [7:0] l18;
	reg [7:0] l19;
	reg [7:0] l20;
	reg [7:0] l21;
	reg [7:0] l22;
	reg [7:0] l23;
	reg [7:0] l24;
	reg [7:0] l25;
	reg [7:0] l26;
	reg [7:0] l27;
	reg [7:0] l28;
	reg [7:0] l29;
	reg [7:0] l30;
	reg [7:0] l31;
	reg [7:0] o0;
	reg [7:0] o1;
	reg [7:0] o2;
	reg [7:0] o3;
	reg [7:0] o4;
	reg [7:0] o5;
	reg [7:0] o6;
	reg [7:0] o7;
	reg [7:0] o8;
	reg [7:0] o9;
	reg [7:0] o10;
	reg [7:0] o11;
	reg [7:0] o12;
	reg [7:0] o13;
	reg [7:0] o14;
	reg [7:0] o15;
	reg [7:0] o16;
	reg [7:0] o17;
	reg [7:0] o18;
	reg [7:0] o19;
	reg [7:0] o20;
	reg [7:0] o21;
	reg [7:0] o22;
	reg [7:0] o23;
	reg [7:0] o24;
	reg [7:0] o25;
	reg [7:0] o26;
	reg [7:0] o27;
	reg [7:0] o28;
	reg [7:0] o29;
	reg [7:0] o30;
	reg [7:0] o31;
	reg [7:0] odd, numerator;
	wire [7:0] tmp;
	integer j;

	rsdec_chien_scale0 x0 (scale0, data0);
	rsdec_chien_scale1 x1 (scale1, data1);
	rsdec_chien_scale2 x2 (scale2, data2);
	rsdec_chien_scale3 x3 (scale3, data3);
	rsdec_chien_scale4 x4 (scale4, data4);
	rsdec_chien_scale5 x5 (scale5, data5);
	rsdec_chien_scale6 x6 (scale6, data6);
	rsdec_chien_scale7 x7 (scale7, data7);
	rsdec_chien_scale8 x8 (scale8, data8);
	rsdec_chien_scale9 x9 (scale9, data9);
	rsdec_chien_scale10 x10 (scale10, data10);
	rsdec_chien_scale11 x11 (scale11, data11);
	rsdec_chien_scale12 x12 (scale12, data12);
	rsdec_chien_scale13 x13 (scale13, data13);
	rsdec_chien_scale14 x14 (scale14, data14);
	rsdec_chien_scale15 x15 (scale15, data15);
	rsdec_chien_scale16 x16 (scale16, data16);
	rsdec_chien_scale17 x17 (scale17, data17);
	rsdec_chien_scale18 x18 (scale18, data18);
	rsdec_chien_scale19 x19 (scale19, data19);
	rsdec_chien_scale20 x20 (scale20, data20);
	rsdec_chien_scale21 x21 (scale21, data21);
	rsdec_chien_scale22 x22 (scale22, data22);
	rsdec_chien_scale23 x23 (scale23, data23);
	rsdec_chien_scale24 x24 (scale24, data24);
	rsdec_chien_scale25 x25 (scale25, data25);
	rsdec_chien_scale26 x26 (scale26, data26);
	rsdec_chien_scale27 x27 (scale27, data27);
	rsdec_chien_scale28 x28 (scale28, data28);
	rsdec_chien_scale29 x29 (scale29, data29);
	rsdec_chien_scale30 x30 (scale30, data30);
	rsdec_chien_scale31 x31 (scale31, data31);
	rsdec_chien_scale0 x32 (scale32, o0);
	rsdec_chien_scale1 x33 (scale33, o1);
	rsdec_chien_scale2 x34 (scale34, o2);
	rsdec_chien_scale3 x35 (scale35, o3);
	rsdec_chien_scale4 x36 (scale36, o4);
	rsdec_chien_scale5 x37 (scale37, o5);
	rsdec_chien_scale6 x38 (scale38, o6);
	rsdec_chien_scale7 x39 (scale39, o7);
	rsdec_chien_scale8 x40 (scale40, o8);
	rsdec_chien_scale9 x41 (scale41, o9);
	rsdec_chien_scale10 x42 (scale42, o10);
	rsdec_chien_scale11 x43 (scale43, o11);
	rsdec_chien_scale12 x44 (scale44, o12);
	rsdec_chien_scale13 x45 (scale45, o13);
	rsdec_chien_scale14 x46 (scale46, o14);
	rsdec_chien_scale15 x47 (scale47, o15);
	rsdec_chien_scale16 x48 (scale48, o16);
	rsdec_chien_scale17 x49 (scale49, o17);
	rsdec_chien_scale18 x50 (scale50, o18);
	rsdec_chien_scale19 x51 (scale51, o19);
	rsdec_chien_scale20 x52 (scale52, o20);
	rsdec_chien_scale21 x53 (scale53, o21);
	rsdec_chien_scale22 x54 (scale54, o22);
	rsdec_chien_scale23 x55 (scale55, o23);
	rsdec_chien_scale24 x56 (scale56, o24);
	rsdec_chien_scale25 x57 (scale57, o25);
	rsdec_chien_scale26 x58 (scale58, o26);
	rsdec_chien_scale27 x59 (scale59, o27);
	rsdec_chien_scale28 x60 (scale60, o28);
	rsdec_chien_scale29 x61 (scale61, o29);
	rsdec_chien_scale30 x62 (scale62, o30);
	rsdec_chien_scale31 x63 (scale63, o31);

	always @ (shorten or a0 or l0)
		if (shorten) data0 = a0;
		else data0 = l0;

	always @ (shorten or a1 or l1)
		if (shorten) data1 = a1;
		else data1 = l1;

	always @ (shorten or a2 or l2)
		if (shorten) data2 = a2;
		else data2 = l2;

	always @ (shorten or a3 or l3)
		if (shorten) data3 = a3;
		else data3 = l3;

	always @ (shorten or a4 or l4)
		if (shorten) data4 = a4;
		else data4 = l4;

	always @ (shorten or a5 or l5)
		if (shorten) data5 = a5;
		else data5 = l5;

	always @ (shorten or a6 or l6)
		if (shorten) data6 = a6;
		else data6 = l6;

	always @ (shorten or a7 or l7)
		if (shorten) data7 = a7;
		else data7 = l7;

	always @ (shorten or a8 or l8)
		if (shorten) data8 = a8;
		else data8 = l8;

	always @ (shorten or a9 or l9)
		if (shorten) data9 = a9;
		else data9 = l9;

	always @ (shorten or a10 or l10)
		if (shorten) data10 = a10;
		else data10 = l10;

	always @ (shorten or a11 or l11)
		if (shorten) data11 = a11;
		else data11 = l11;

	always @ (shorten or a12 or l12)
		if (shorten) data12 = a12;
		else data12 = l12;

	always @ (shorten or a13 or l13)
		if (shorten) data13 = a13;
		else data13 = l13;

	always @ (shorten or a14 or l14)
		if (shorten) data14 = a14;
		else data14 = l14;

	always @ (shorten or a15 or l15)
		if (shorten) data15 = a15;
		else data15 = l15;

	always @ (shorten or a16 or l16)
		if (shorten) data16 = a16;
		else data16 = l16;

	always @ (shorten or a17 or l17)
		if (shorten) data17 = a17;
		else data17 = l17;

	always @ (shorten or a18 or l18)
		if (shorten) data18 = a18;
		else data18 = l18;

	always @ (shorten or a19 or l19)
		if (shorten) data19 = a19;
		else data19 = l19;

	always @ (shorten or a20 or l20)
		if (shorten) data20 = a20;
		else data20 = l20;

	always @ (shorten or a21 or l21)
		if (shorten) data21 = a21;
		else data21 = l21;

	always @ (shorten or a22 or l22)
		if (shorten) data22 = a22;
		else data22 = l22;

	always @ (shorten or a23 or l23)
		if (shorten) data23 = a23;
		else data23 = l23;

	always @ (shorten or a24 or l24)
		if (shorten) data24 = a24;
		else data24 = l24;

	always @ (shorten or a25 or l25)
		if (shorten) data25 = a25;
		else data25 = l25;

	always @ (shorten or a26 or l26)
		if (shorten) data26 = a26;
		else data26 = l26;

	always @ (shorten or a27 or l27)
		if (shorten) data27 = a27;
		else data27 = l27;

	always @ (shorten or a28 or l28)
		if (shorten) data28 = a28;
		else data28 = l28;

	always @ (shorten or a29 or l29)
		if (shorten) data29 = a29;
		else data29 = l29;

	always @ (shorten or a30 or l30)
		if (shorten) data30 = a30;
		else data30 = l30;

	always @ (shorten or a31 or l31)
		if (shorten) data31 = a31;
		else data31 = l31;

	always @ (posedge clk or negedge clrn)
	begin
		if (~clrn)
		begin
			l0 <= 0;
			l1 <= 0;
			l2 <= 0;
			l3 <= 0;
			l4 <= 0;
			l5 <= 0;
			l6 <= 0;
			l7 <= 0;
			l8 <= 0;
			l9 <= 0;
			l10 <= 0;
			l11 <= 0;
			l12 <= 0;
			l13 <= 0;
			l14 <= 0;
			l15 <= 0;
			l16 <= 0;
			l17 <= 0;
			l18 <= 0;
			l19 <= 0;
			l20 <= 0;
			l21 <= 0;
			l22 <= 0;
			l23 <= 0;
			l24 <= 0;
			l25 <= 0;
			l26 <= 0;
			l27 <= 0;
			l28 <= 0;
			l29 <= 0;
			l30 <= 0;
			l31 <= 0;
			o0 <= 0;
			o1 <= 0;
			o2 <= 0;
			o3 <= 0;
			o4 <= 0;
			o5 <= 0;
			o6 <= 0;
			o7 <= 0;
			o8 <= 0;
			o9 <= 0;
			o10 <= 0;
			o11 <= 0;
			o12 <= 0;
			o13 <= 0;
			o14 <= 0;
			o15 <= 0;
			o16 <= 0;
			o17 <= 0;
			o18 <= 0;
			o19 <= 0;
			o20 <= 0;
			o21 <= 0;
			o22 <= 0;
			o23 <= 0;
			o24 <= 0;
			o25 <= 0;
			o26 <= 0;
			o27 <= 0;
			o28 <= 0;
			o29 <= 0;
			o30 <= 0;
			o31 <= 0;
			a0 <= 1;
			a1 <= 1;
			a2 <= 1;
			a3 <= 1;
			a4 <= 1;
			a5 <= 1;
			a6 <= 1;
			a7 <= 1;
			a8 <= 1;
			a9 <= 1;
			a10 <= 1;
			a11 <= 1;
			a12 <= 1;
			a13 <= 1;
			a14 <= 1;
			a15 <= 1;
			a16 <= 1;
			a17 <= 1;
			a18 <= 1;
			a19 <= 1;
			a20 <= 1;
			a21 <= 1;
			a22 <= 1;
			a23 <= 1;
			a24 <= 1;
			a25 <= 1;
			a26 <= 1;
			a27 <= 1;
			a28 <= 1;
			a29 <= 1;
			a30 <= 1;
			a31 <= 1;
		end
		else if (shorten)
		begin
			a0 <= scale0;
			a1 <= scale1;
			a2 <= scale2;
			a3 <= scale3;
			a4 <= scale4;
			a5 <= scale5;
			a6 <= scale6;
			a7 <= scale7;
			a8 <= scale8;
			a9 <= scale9;
			a10 <= scale10;
			a11 <= scale11;
			a12 <= scale12;
			a13 <= scale13;
			a14 <= scale14;
			a15 <= scale15;
			a16 <= scale16;
			a17 <= scale17;
			a18 <= scale18;
			a19 <= scale19;
			a20 <= scale20;
			a21 <= scale21;
			a22 <= scale22;
			a23 <= scale23;
			a24 <= scale24;
			a25 <= scale25;
			a26 <= scale26;
			a27 <= scale27;
			a28 <= scale28;
			a29 <= scale29;
			a30 <= scale30;
			a31 <= scale31;
		end
		else if (search)
		begin
			l0 <= scale0;
			l1 <= scale1;
			l2 <= scale2;
			l3 <= scale3;
			l4 <= scale4;
			l5 <= scale5;
			l6 <= scale6;
			l7 <= scale7;
			l8 <= scale8;
			l9 <= scale9;
			l10 <= scale10;
			l11 <= scale11;
			l12 <= scale12;
			l13 <= scale13;
			l14 <= scale14;
			l15 <= scale15;
			l16 <= scale16;
			l17 <= scale17;
			l18 <= scale18;
			l19 <= scale19;
			l20 <= scale20;
			l21 <= scale21;
			l22 <= scale22;
			l23 <= scale23;
			l24 <= scale24;
			l25 <= scale25;
			l26 <= scale26;
			l27 <= scale27;
			l28 <= scale28;
			l29 <= scale29;
			l30 <= scale30;
			l31 <= scale31;
			o0 <= scale32;
			o1 <= scale33;
			o2 <= scale34;
			o3 <= scale35;
			o4 <= scale36;
			o5 <= scale37;
			o6 <= scale38;
			o7 <= scale39;
			o8 <= scale40;
			o9 <= scale41;
			o10 <= scale42;
			o11 <= scale43;
			o12 <= scale44;
			o13 <= scale45;
			o14 <= scale46;
			o15 <= scale47;
			o16 <= scale48;
			o17 <= scale49;
			o18 <= scale50;
			o19 <= scale51;
			o20 <= scale52;
			o21 <= scale53;
			o22 <= scale54;
			o23 <= scale55;
			o24 <= scale56;
			o25 <= scale57;
			o26 <= scale58;
			o27 <= scale59;
			o28 <= scale60;
			o29 <= scale61;
			o30 <= scale62;
			o31 <= scale63;
		end
		else if (load)
		begin
			l0 <= lambda;
			l1 <= l0;
			l2 <= l1;
			l3 <= l2;
			l4 <= l3;
			l5 <= l4;
			l6 <= l5;
			l7 <= l6;
			l8 <= l7;
			l9 <= l8;
			l10 <= l9;
			l11 <= l10;
			l12 <= l11;
			l13 <= l12;
			l14 <= l13;
			l15 <= l14;
			l16 <= l15;
			l17 <= l16;
			l18 <= l17;
			l19 <= l18;
			l20 <= l19;
			l21 <= l20;
			l22 <= l21;
			l23 <= l22;
			l24 <= l23;
			l25 <= l24;
			l26 <= l25;
			l27 <= l26;
			l28 <= l27;
			l29 <= l28;
			l30 <= l29;
			l31 <= l30;
			o0 <= omega;
			o1 <= o0;
			o2 <= o1;
			o3 <= o2;
			o4 <= o3;
			o5 <= o4;
			o6 <= o5;
			o7 <= o6;
			o8 <= o7;
			o9 <= o8;
			o10 <= o9;
			o11 <= o10;
			o12 <= o11;
			o13 <= o12;
			o14 <= o13;
			o15 <= o14;
			o16 <= o15;
			o17 <= o16;
			o18 <= o17;
			o19 <= o18;
			o20 <= o19;
			o21 <= o20;
			o22 <= o21;
			o23 <= o22;
			o24 <= o23;
			o25 <= o24;
			o26 <= o25;
			o27 <= o26;
			o28 <= o27;
			o29 <= o28;
			o30 <= o29;
			o31 <= o30;
			a0 <= a31;
			a1 <= a0;
			a2 <= a1;
			a3 <= a2;
			a4 <= a3;
			a5 <= a4;
			a6 <= a5;
			a7 <= a6;
			a8 <= a7;
			a9 <= a8;
			a10 <= a9;
			a11 <= a10;
			a12 <= a11;
			a13 <= a12;
			a14 <= a13;
			a15 <= a14;
			a16 <= a15;
			a17 <= a16;
			a18 <= a17;
			a19 <= a18;
			a20 <= a19;
			a21 <= a20;
			a22 <= a21;
			a23 <= a22;
			a24 <= a23;
			a25 <= a24;
			a26 <= a25;
			a27 <= a26;
			a28 <= a27;
			a29 <= a28;
			a30 <= a29;
			a31 <= a30;
		end
	end

	always @ (l0 or l2 or l4 or l6 or l8 or l10 or l12 or l14 or l16 or l18 or l20 or l22 or l24 or l26 or l28 or l30)
		even = l0 ^ l2 ^ l4 ^ l6 ^ l8 ^ l10 ^ l12 ^ l14 ^ l16 ^ l18 ^ l20 ^ l22 ^ l24 ^ l26 ^ l28 ^ l30;

	always @ (l1 or l3 or l5 or l7 or l9 or l11 or l13 or l15 or l17 or l19 or l21 or l23 or l25 or l27 or l29 or l31)
		odd = l1 ^ l3 ^ l5 ^ l7 ^ l9 ^ l11 ^ l13 ^ l15 ^ l17 ^ l19 ^ l21 ^ l23 ^ l25 ^ l27 ^ l29 ^ l31;

	always @ (o0 or o1 or o2 or o3 or o4 or o5 or o6 or o7 or o8 or o9 or o10 or o11 or o12 or o13 or o14 or o15 or o16 or o17 or o18 or o19 or o20 or o21 or o22 or o23 or o24 or o25 or o26 or o27 or o28 or o29 or o30 or o31)
		numerator = o0 ^ o1 ^ o2 ^ o3 ^ o4 ^ o5 ^ o6 ^ o7 ^ o8 ^ o9 ^ o10 ^ o11 ^ o12 ^ o13 ^ o14 ^ o15 ^ o16 ^ o17 ^ o18 ^ o19 ^ o20 ^ o21 ^ o22 ^ o23 ^ o24 ^ o25 ^ o26 ^ o27 ^ o28 ^ o29 ^ o30 ^ o31;

	multiply m0 (tmp, numerator, D);

	always @ (even or odd or tmp)
		if (even == odd) error = tmp;
		else error = 0;

	always @ (a31) alpha = a31;

endmodule



// -------------------------------------------------------------------------
// a sample ROM, feeding data to encoder
//Copyright (C) Tue Apr  2 14:40:09 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module sigin(data, address);
	input [7:0] address;
	output [7:0] data;
	reg [7:0] data;
	
	// an arbitrary data source here
	always @ (address) data = address + 1;
endmodule



// -------------------------------------------------------------------------
//The inverse lookup table for Galois field
//Copyright (C) Tue Apr  2 17:07:28 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module inverse(y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	case (x) // synopsys full_case parallel_case
		1: y = 1; // 0 -> 255
		2: y = 195; // 1 -> 254
		4: y = 162; // 2 -> 253
		8: y = 81; // 3 -> 252
		16: y = 235; // 4 -> 251
		32: y = 182; // 5 -> 250
		64: y = 91; // 6 -> 249
		128: y = 238; // 7 -> 248
		135: y = 119; // 8 -> 247
		137: y = 248; // 9 -> 246
		149: y = 124; // 10 -> 245
		173: y = 62; // 11 -> 244
		221: y = 31; // 12 -> 243
		61: y = 204; // 13 -> 242
		122: y = 102; // 14 -> 241
		244: y = 51; // 15 -> 240
		111: y = 218; // 16 -> 239
		222: y = 109; // 17 -> 238
		59: y = 245; // 18 -> 237
		118: y = 185; // 19 -> 236
		236: y = 159; // 20 -> 235
		95: y = 140; // 21 -> 234
		190: y = 70; // 22 -> 233
		251: y = 35; // 23 -> 232
		113: y = 210; // 24 -> 231
		226: y = 105; // 25 -> 230
		67: y = 247; // 26 -> 229
		134: y = 184; // 27 -> 228
		139: y = 92; // 28 -> 227
		145: y = 46; // 29 -> 226
		165: y = 23; // 30 -> 225
		205: y = 200; // 31 -> 224
		29: y = 100; // 32 -> 223
		58: y = 50; // 33 -> 222
		116: y = 25; // 34 -> 221
		232: y = 207; // 35 -> 220
		87: y = 164; // 36 -> 219
		174: y = 82; // 37 -> 218
		219: y = 41; // 38 -> 217
		49: y = 215; // 39 -> 216
		98: y = 168; // 40 -> 215
		196: y = 84; // 41 -> 214
		15: y = 42; // 42 -> 213
		30: y = 21; // 43 -> 212
		60: y = 201; // 44 -> 211
		120: y = 167; // 45 -> 210
		240: y = 144; // 46 -> 209
		103: y = 72; // 47 -> 208
		206: y = 36; // 48 -> 207
		27: y = 18; // 49 -> 206
		54: y = 9; // 50 -> 205
		108: y = 199; // 51 -> 204
		216: y = 160; // 52 -> 203
		55: y = 80; // 53 -> 202
		110: y = 40; // 54 -> 201
		220: y = 20; // 55 -> 200
		63: y = 10; // 56 -> 199
		126: y = 5; // 57 -> 198
		252: y = 193; // 58 -> 197
		127: y = 163; // 59 -> 196
		254: y = 146; // 60 -> 195
		123: y = 73; // 61 -> 194
		246: y = 231; // 62 -> 193
		107: y = 176; // 63 -> 192
		214: y = 88; // 64 -> 191
		43: y = 44; // 65 -> 190
		86: y = 22; // 66 -> 189
		172: y = 11; // 67 -> 188
		223: y = 198; // 68 -> 187
		57: y = 99; // 69 -> 186
		114: y = 242; // 70 -> 185
		228: y = 121; // 71 -> 184
		79: y = 255; // 72 -> 183
		158: y = 188; // 73 -> 182
		187: y = 94; // 74 -> 181
		241: y = 47; // 75 -> 180
		101: y = 212; // 76 -> 179
		202: y = 106; // 77 -> 178
		19: y = 53; // 78 -> 177
		38: y = 217; // 79 -> 176
		76: y = 175; // 80 -> 175
		152: y = 148; // 81 -> 174
		183: y = 74; // 82 -> 173
		233: y = 37; // 83 -> 172
		85: y = 209; // 84 -> 171
		170: y = 171; // 85 -> 170
		211: y = 150; // 86 -> 169
		33: y = 75; // 87 -> 168
		66: y = 230; // 88 -> 167
		132: y = 115; // 89 -> 166
		143: y = 250; // 90 -> 165
		153: y = 125; // 91 -> 164
		181: y = 253; // 92 -> 163
		237: y = 189; // 93 -> 162
		93: y = 157; // 94 -> 161
		186: y = 141; // 95 -> 160
		243: y = 133; // 96 -> 159
		97: y = 129; // 97 -> 158
		194: y = 131; // 98 -> 157
		3: y = 130; // 99 -> 156
		6: y = 65; // 100 -> 155
		12: y = 227; // 101 -> 154
		24: y = 178; // 102 -> 153
		48: y = 89; // 103 -> 152
		96: y = 239; // 104 -> 151
		192: y = 180; // 105 -> 150
		7: y = 90; // 106 -> 149
		14: y = 45; // 107 -> 148
		28: y = 213; // 108 -> 147
		56: y = 169; // 109 -> 146
		112: y = 151; // 110 -> 145
		224: y = 136; // 111 -> 144
		71: y = 68; // 112 -> 143
		142: y = 34; // 113 -> 142
		155: y = 17; // 114 -> 141
		177: y = 203; // 115 -> 140
		229: y = 166; // 116 -> 139
		77: y = 83; // 117 -> 138
		154: y = 234; // 118 -> 137
		179: y = 117; // 119 -> 136
		225: y = 249; // 120 -> 135
		69: y = 191; // 121 -> 134
		138: y = 156; // 122 -> 133
		147: y = 78; // 123 -> 132
		161: y = 39; // 124 -> 131
		197: y = 208; // 125 -> 130
		13: y = 104; // 126 -> 129
		26: y = 52; // 127 -> 128
		52: y = 26; // 128 -> 127
		104: y = 13; // 129 -> 126
		208: y = 197; // 130 -> 125
		39: y = 161; // 131 -> 124
		78: y = 147; // 132 -> 123
		156: y = 138; // 133 -> 122
		191: y = 69; // 134 -> 121
		249: y = 225; // 135 -> 120
		117: y = 179; // 136 -> 119
		234: y = 154; // 137 -> 118
		83: y = 77; // 138 -> 117
		166: y = 229; // 139 -> 116
		203: y = 177; // 140 -> 115
		17: y = 155; // 141 -> 114
		34: y = 142; // 142 -> 113
		68: y = 71; // 143 -> 112
		136: y = 224; // 144 -> 111
		151: y = 112; // 145 -> 110
		169: y = 56; // 146 -> 109
		213: y = 28; // 147 -> 108
		45: y = 14; // 148 -> 107
		90: y = 7; // 149 -> 106
		180: y = 192; // 150 -> 105
		239: y = 96; // 151 -> 104
		89: y = 48; // 152 -> 103
		178: y = 24; // 153 -> 102
		227: y = 12; // 154 -> 101
		65: y = 6; // 155 -> 100
		130: y = 3; // 156 -> 99
		131: y = 194; // 157 -> 98
		129: y = 97; // 158 -> 97
		133: y = 243; // 159 -> 96
		141: y = 186; // 160 -> 95
		157: y = 93; // 161 -> 94
		189: y = 237; // 162 -> 93
		253: y = 181; // 163 -> 92
		125: y = 153; // 164 -> 91
		250: y = 143; // 165 -> 90
		115: y = 132; // 166 -> 89
		230: y = 66; // 167 -> 88
		75: y = 33; // 168 -> 87
		150: y = 211; // 169 -> 86
		171: y = 170; // 170 -> 85
		209: y = 85; // 171 -> 84
		37: y = 233; // 172 -> 83
		74: y = 183; // 173 -> 82
		148: y = 152; // 174 -> 81
		175: y = 76; // 175 -> 80
		217: y = 38; // 176 -> 79
		53: y = 19; // 177 -> 78
		106: y = 202; // 178 -> 77
		212: y = 101; // 179 -> 76
		47: y = 241; // 180 -> 75
		94: y = 187; // 181 -> 74
		188: y = 158; // 182 -> 73
		255: y = 79; // 183 -> 72
		121: y = 228; // 184 -> 71
		242: y = 114; // 185 -> 70
		99: y = 57; // 186 -> 69
		198: y = 223; // 187 -> 68
		11: y = 172; // 188 -> 67
		22: y = 86; // 189 -> 66
		44: y = 43; // 190 -> 65
		88: y = 214; // 191 -> 64
		176: y = 107; // 192 -> 63
		231: y = 246; // 193 -> 62
		73: y = 123; // 194 -> 61
		146: y = 254; // 195 -> 60
		163: y = 127; // 196 -> 59
		193: y = 252; // 197 -> 58
		5: y = 126; // 198 -> 57
		10: y = 63; // 199 -> 56
		20: y = 220; // 200 -> 55
		40: y = 110; // 201 -> 54
		80: y = 55; // 202 -> 53
		160: y = 216; // 203 -> 52
		199: y = 108; // 204 -> 51
		9: y = 54; // 205 -> 50
		18: y = 27; // 206 -> 49
		36: y = 206; // 207 -> 48
		72: y = 103; // 208 -> 47
		144: y = 240; // 209 -> 46
		167: y = 120; // 210 -> 45
		201: y = 60; // 211 -> 44
		21: y = 30; // 212 -> 43
		42: y = 15; // 213 -> 42
		84: y = 196; // 214 -> 41
		168: y = 98; // 215 -> 40
		215: y = 49; // 216 -> 39
		41: y = 219; // 217 -> 38
		82: y = 174; // 218 -> 37
		164: y = 87; // 219 -> 36
		207: y = 232; // 220 -> 35
		25: y = 116; // 221 -> 34
		50: y = 58; // 222 -> 33
		100: y = 29; // 223 -> 32
		200: y = 205; // 224 -> 31
		23: y = 165; // 225 -> 30
		46: y = 145; // 226 -> 29
		92: y = 139; // 227 -> 28
		184: y = 134; // 228 -> 27
		247: y = 67; // 229 -> 26
		105: y = 226; // 230 -> 25
		210: y = 113; // 231 -> 24
		35: y = 251; // 232 -> 23
		70: y = 190; // 233 -> 22
		140: y = 95; // 234 -> 21
		159: y = 236; // 235 -> 20
		185: y = 118; // 236 -> 19
		245: y = 59; // 237 -> 18
		109: y = 222; // 238 -> 17
		218: y = 111; // 239 -> 16
		51: y = 244; // 240 -> 15
		102: y = 122; // 241 -> 14
		204: y = 61; // 242 -> 13
		31: y = 221; // 243 -> 12
		62: y = 173; // 244 -> 11
		124: y = 149; // 245 -> 10
		248: y = 137; // 246 -> 9
		119: y = 135; // 247 -> 8
		238: y = 128; // 248 -> 7
		91: y = 64; // 249 -> 6
		182: y = 32; // 250 -> 5
		235: y = 16; // 251 -> 4
		81: y = 8; // 252 -> 3
		162: y = 4; // 253 -> 2
		195: y = 2; // 254 -> 1
		default: y = 0;
	endcase
endmodule


// -------------------------------------------------------------------------
//Syndrome generator circuit in Reed-Solomon Decoder
//Copyright (C) Tue Apr  2 17:07:53 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module rsdec_syn_m0 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[7];
		y[1] = x[0] ^ x[7];
		y[2] = x[1] ^ x[7];
		y[3] = x[2];
		y[4] = x[3];
		y[5] = x[4];
		y[6] = x[5];
		y[7] = x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m1 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[6] ^ x[7];
		y[1] = x[6];
		y[2] = x[0] ^ x[6];
		y[3] = x[1] ^ x[7];
		y[4] = x[2];
		y[5] = x[3];
		y[6] = x[4];
		y[7] = x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m2 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[5] ^ x[6] ^ x[7];
		y[1] = x[5];
		y[2] = x[5] ^ x[7];
		y[3] = x[0] ^ x[6];
		y[4] = x[1] ^ x[7];
		y[5] = x[2];
		y[6] = x[3];
		y[7] = x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m3 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[4];
		y[2] = x[4] ^ x[6] ^ x[7];
		y[3] = x[5] ^ x[7];
		y[4] = x[0] ^ x[6];
		y[5] = x[1] ^ x[7];
		y[6] = x[2];
		y[7] = x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m4 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[3];
		y[2] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[4] ^ x[6] ^ x[7];
		y[4] = x[5] ^ x[7];
		y[5] = x[0] ^ x[6];
		y[6] = x[1] ^ x[7];
		y[7] = x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m5 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[2];
		y[2] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[4] ^ x[6] ^ x[7];
		y[5] = x[5] ^ x[7];
		y[6] = x[0] ^ x[6];
		y[7] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_syn_m6 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[1] = x[1] ^ x[7];
		y[2] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[4] ^ x[6] ^ x[7];
		y[6] = x[5] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
	end
endmodule

module rsdec_syn_m7 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[1] = x[0] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[4] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
	end
endmodule

module rsdec_syn_m8 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
		y[1] = x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6];
	end
endmodule

module rsdec_syn_m9 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6];
		y[1] = x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_syn_m10 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[7];
		y[1] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[6] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[4] ^ x[6];
	end
endmodule

module rsdec_syn_m11 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[4] ^ x[6];
		y[1] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[0] ^ x[3] ^ x[5];
	end
endmodule

module rsdec_syn_m12 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[5];
		y[1] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[4] ^ x[7];
	end
endmodule

module rsdec_syn_m13 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[2] ^ x[4] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[6];
	end
endmodule

module rsdec_syn_m14 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[6];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_syn_m15 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[1] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m16 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[4] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[3] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_syn_m17 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[5] ^ x[6];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[4] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_syn_m18 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[2] ^ x[4] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[4] ^ x[6];
	end
endmodule

module rsdec_syn_m19 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[4] ^ x[6];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[6] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_syn_m20 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[7] = x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m21 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[5];
		y[3] = x[0] ^ x[1] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m22 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[2] = x[4] ^ x[7];
		y[3] = x[0] ^ x[5];
		y[4] = x[0] ^ x[1] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[7] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m23 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[2] = x[3] ^ x[6] ^ x[7];
		y[3] = x[4] ^ x[7];
		y[4] = x[0] ^ x[5];
		y[5] = x[0] ^ x[1] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m24 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[2] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[3] ^ x[6] ^ x[7];
		y[4] = x[4] ^ x[7];
		y[5] = x[0] ^ x[5];
		y[6] = x[0] ^ x[1] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_syn_m25 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[2] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[3] ^ x[6] ^ x[7];
		y[5] = x[4] ^ x[7];
		y[6] = x[0] ^ x[5];
		y[7] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
	end
endmodule

module rsdec_syn_m26 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[1] = x[0] ^ x[1] ^ x[6];
		y[2] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[3] ^ x[6] ^ x[7];
		y[6] = x[4] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4];
	end
endmodule

module rsdec_syn_m27 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4];
		y[1] = x[0] ^ x[5];
		y[2] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[3] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[3] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[7];
	end
endmodule

module rsdec_syn_m28 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[7];
		y[1] = x[4] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[3] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[4] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[6];
	end
endmodule

module rsdec_syn_m29 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[6];
		y[1] = x[3] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[4] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[5] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[6] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[5] ^ x[7];
	end
endmodule

module rsdec_syn_m30 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[5] ^ x[7];
		y[1] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[5] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[6] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[0] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rsdec_syn_m31 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[4] ^ x[6] ^ x[7];
		y[1] = x[1] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[4] ^ x[5];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[6] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[7] = x[3] ^ x[5] ^ x[6];
	end
endmodule

module rsdec_syn (y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, u, enable, shift, init, clk, clrn);
	input [7:0] u;
	input clk, clrn, shift, init, enable;
	output [7:0] y0;
	output [7:0] y1;
	output [7:0] y2;
	output [7:0] y3;
	output [7:0] y4;
	output [7:0] y5;
	output [7:0] y6;
	output [7:0] y7;
	output [7:0] y8;
	output [7:0] y9;
	output [7:0] y10;
	output [7:0] y11;
	output [7:0] y12;
	output [7:0] y13;
	output [7:0] y14;
	output [7:0] y15;
	output [7:0] y16;
	output [7:0] y17;
	output [7:0] y18;
	output [7:0] y19;
	output [7:0] y20;
	output [7:0] y21;
	output [7:0] y22;
	output [7:0] y23;
	output [7:0] y24;
	output [7:0] y25;
	output [7:0] y26;
	output [7:0] y27;
	output [7:0] y28;
	output [7:0] y29;
	output [7:0] y30;
	output [7:0] y31;
	reg [7:0] y0;
	reg [7:0] y1;
	reg [7:0] y2;
	reg [7:0] y3;
	reg [7:0] y4;
	reg [7:0] y5;
	reg [7:0] y6;
	reg [7:0] y7;
	reg [7:0] y8;
	reg [7:0] y9;
	reg [7:0] y10;
	reg [7:0] y11;
	reg [7:0] y12;
	reg [7:0] y13;
	reg [7:0] y14;
	reg [7:0] y15;
	reg [7:0] y16;
	reg [7:0] y17;
	reg [7:0] y18;
	reg [7:0] y19;
	reg [7:0] y20;
	reg [7:0] y21;
	reg [7:0] y22;
	reg [7:0] y23;
	reg [7:0] y24;
	reg [7:0] y25;
	reg [7:0] y26;
	reg [7:0] y27;
	reg [7:0] y28;
	reg [7:0] y29;
	reg [7:0] y30;
	reg [7:0] y31;

	wire [7:0] scale0;
	wire [7:0] scale1;
	wire [7:0] scale2;
	wire [7:0] scale3;
	wire [7:0] scale4;
	wire [7:0] scale5;
	wire [7:0] scale6;
	wire [7:0] scale7;
	wire [7:0] scale8;
	wire [7:0] scale9;
	wire [7:0] scale10;
	wire [7:0] scale11;
	wire [7:0] scale12;
	wire [7:0] scale13;
	wire [7:0] scale14;
	wire [7:0] scale15;
	wire [7:0] scale16;
	wire [7:0] scale17;
	wire [7:0] scale18;
	wire [7:0] scale19;
	wire [7:0] scale20;
	wire [7:0] scale21;
	wire [7:0] scale22;
	wire [7:0] scale23;
	wire [7:0] scale24;
	wire [7:0] scale25;
	wire [7:0] scale26;
	wire [7:0] scale27;
	wire [7:0] scale28;
	wire [7:0] scale29;
	wire [7:0] scale30;
	wire [7:0] scale31;

	rsdec_syn_m0 m0 (scale0, y0);
	rsdec_syn_m1 m1 (scale1, y1);
	rsdec_syn_m2 m2 (scale2, y2);
	rsdec_syn_m3 m3 (scale3, y3);
	rsdec_syn_m4 m4 (scale4, y4);
	rsdec_syn_m5 m5 (scale5, y5);
	rsdec_syn_m6 m6 (scale6, y6);
	rsdec_syn_m7 m7 (scale7, y7);
	rsdec_syn_m8 m8 (scale8, y8);
	rsdec_syn_m9 m9 (scale9, y9);
	rsdec_syn_m10 m10 (scale10, y10);
	rsdec_syn_m11 m11 (scale11, y11);
	rsdec_syn_m12 m12 (scale12, y12);
	rsdec_syn_m13 m13 (scale13, y13);
	rsdec_syn_m14 m14 (scale14, y14);
	rsdec_syn_m15 m15 (scale15, y15);
	rsdec_syn_m16 m16 (scale16, y16);
	rsdec_syn_m17 m17 (scale17, y17);
	rsdec_syn_m18 m18 (scale18, y18);
	rsdec_syn_m19 m19 (scale19, y19);
	rsdec_syn_m20 m20 (scale20, y20);
	rsdec_syn_m21 m21 (scale21, y21);
	rsdec_syn_m22 m22 (scale22, y22);
	rsdec_syn_m23 m23 (scale23, y23);
	rsdec_syn_m24 m24 (scale24, y24);
	rsdec_syn_m25 m25 (scale25, y25);
	rsdec_syn_m26 m26 (scale26, y26);
	rsdec_syn_m27 m27 (scale27, y27);
	rsdec_syn_m28 m28 (scale28, y28);
	rsdec_syn_m29 m29 (scale29, y29);
	rsdec_syn_m30 m30 (scale30, y30);
	rsdec_syn_m31 m31 (scale31, y31);

	always @ (posedge clk or negedge clrn)
	begin
		if (~clrn)
		begin
			y0 <= 0;
			y1 <= 0;
			y2 <= 0;
			y3 <= 0;
			y4 <= 0;
			y5 <= 0;
			y6 <= 0;
			y7 <= 0;
			y8 <= 0;
			y9 <= 0;
			y10 <= 0;
			y11 <= 0;
			y12 <= 0;
			y13 <= 0;
			y14 <= 0;
			y15 <= 0;
			y16 <= 0;
			y17 <= 0;
			y18 <= 0;
			y19 <= 0;
			y20 <= 0;
			y21 <= 0;
			y22 <= 0;
			y23 <= 0;
			y24 <= 0;
			y25 <= 0;
			y26 <= 0;
			y27 <= 0;
			y28 <= 0;
			y29 <= 0;
			y30 <= 0;
			y31 <= 0;
		end
		else if (init)
		begin
			y0 <= u;
			y1 <= u;
			y2 <= u;
			y3 <= u;
			y4 <= u;
			y5 <= u;
			y6 <= u;
			y7 <= u;
			y8 <= u;
			y9 <= u;
			y10 <= u;
			y11 <= u;
			y12 <= u;
			y13 <= u;
			y14 <= u;
			y15 <= u;
			y16 <= u;
			y17 <= u;
			y18 <= u;
			y19 <= u;
			y20 <= u;
			y21 <= u;
			y22 <= u;
			y23 <= u;
			y24 <= u;
			y25 <= u;
			y26 <= u;
			y27 <= u;
			y28 <= u;
			y29 <= u;
			y30 <= u;
			y31 <= u;
		end
		else if (enable)
		begin
			y0 <= scale0 ^ u;
			y1 <= scale1 ^ u;
			y2 <= scale2 ^ u;
			y3 <= scale3 ^ u;
			y4 <= scale4 ^ u;
			y5 <= scale5 ^ u;
			y6 <= scale6 ^ u;
			y7 <= scale7 ^ u;
			y8 <= scale8 ^ u;
			y9 <= scale9 ^ u;
			y10 <= scale10 ^ u;
			y11 <= scale11 ^ u;
			y12 <= scale12 ^ u;
			y13 <= scale13 ^ u;
			y14 <= scale14 ^ u;
			y15 <= scale15 ^ u;
			y16 <= scale16 ^ u;
			y17 <= scale17 ^ u;
			y18 <= scale18 ^ u;
			y19 <= scale19 ^ u;
			y20 <= scale20 ^ u;
			y21 <= scale21 ^ u;
			y22 <= scale22 ^ u;
			y23 <= scale23 ^ u;
			y24 <= scale24 ^ u;
			y25 <= scale25 ^ u;
			y26 <= scale26 ^ u;
			y27 <= scale27 ^ u;
			y28 <= scale28 ^ u;
			y29 <= scale29 ^ u;
			y30 <= scale30 ^ u;
			y31 <= scale31 ^ u;
		end
		else if (shift)
		begin
			y0 <= y1;
			y1 <= y2;
			y2 <= y3;
			y3 <= y4;
			y4 <= y5;
			y5 <= y6;
			y6 <= y7;
			y7 <= y8;
			y8 <= y9;
			y9 <= y10;
			y10 <= y11;
			y11 <= y12;
			y12 <= y13;
			y13 <= y14;
			y14 <= y15;
			y15 <= y16;
			y16 <= y17;
			y17 <= y18;
			y18 <= y19;
			y19 <= y20;
			y20 <= y21;
			y21 <= y22;
			y22 <= y23;
			y23 <= y24;
			y24 <= y25;
			y25 <= y26;
			y26 <= y27;
			y27 <= y28;
			y28 <= y29;
			y29 <= y30;
			y30 <= y31;
			y31 <= y0;
		end
	end

endmodule


module AP0BP1 (    
    input wire clk,        
    input wire rst_n,     
    input wire A,          
    input wire B,          
    output reg C           
);

// 用于保存A和B信号前一个状态的寄存器  
reg A_prev, B_prev;
// 初始化输出C  

  
// 上升沿检测逻辑  
always @(posedge clk or negedge rst_n) begin  
    if (!rst_n) begin  
        // 如果复位信号有效，将C复位到初始状态  
        C <= 0; // 或者 1，取决于你的复位逻辑  
    end else begin  
        // 检查A和B的上升沿  
        if (A && ~A_prev) begin  
            // 当A从0变为1时，将C置为低  
            C <= 0;  
        end else if (B && ~B_prev) begin  
            // 当B从0变为1时，将C置为高  
            C <= 1;  
        end  
    end  
end  
  
  
  
// 在时钟上升沿更新A和B的前一个状态  
always @(posedge clk or negedge rst_n) begin  
    if (!rst_n) begin  
        // 复位时，将A和B的前一个状态都设置为0  
        A_prev <= 0;  
        B_prev <= 0;  
    end else begin  
        // 在每个时钟上升沿，保存A和B的当前状态  
        A_prev <= A;  
        B_prev <= B;  
    end  
end  
  
endmodule




module LUT1 #(parameter INIT = 2'h0) (
    output O,
    input I0
);

    INVD0BWP40P140HVT u_inv (
        .I(I0),
        .ZN(O)
    );
    // assign O=I0;

endmodule

module LUT3 #(parameter INIT = 8'h00) (
    output O,
    input I0,
    input I1,
    input I2
);

    ND3D0BWP40P140HVT u_nand3 (
        .ZN(O),
        .A1(I0),
        .A2(I1),
        .A3(I2)
    );

endmodule

// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/30 10:46:11
// Design Name:
// Module Name: Comp
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Comp(
    input clk,
    input rst,
    input [31:0] num1,
    input [31:0] num2,
    input comp_en,
    output reg done,
    output reg [1:0] result
);

//can add a mode signle to change comp mode
reg [31:0] num1_reg;
reg [31:0] num2_reg;

always @(posedge clk or negedge rst) begin
    if(!rst) begin
        done <= 0;
        result <= 2'd0;
        num1_reg <= 32'd0;
        num2_reg <= 32'd0;
    end else begin
        if(comp_en) begin
            num1_reg <= num1;
            num2_reg <= num2;
            if(num1 > num2) begin
                done <= 1;
                result <= 2'b11;
            end else if(num1 == num2) begin
                done <= 1;
                result <= 2'b01;
            end else begin
                done <= 1;
                result <= 2'b00;
            end
        end else begin
            done <= 0;
            result <= 2'b00;
            num1_reg <= 32'd0;
            num2_reg <= 32'd0;
        end
    end
end

endmodule





// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/29 16:58:55
// Design Name:
// Module Name: Counter
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module Counter(
    input cnt_in,                //counter clk
    input clk,
    input rst,
    input cnt_ctrl,             //cnt_ctrl=1, counter start; cnt_ctrl=0,counter stop
    input clear,                //clear = 1,cnt_out reset to 0; else cnt_out retain
    output done,                //cnt_ctrl transmit form 1 to 0, than done=1
    output reg [31:0] cnt_out
);

    reg done_reg;
    // reg cnt_flag;
    reg cnt_ctrl_delayed;

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            done_reg <= 1'b0;
            cnt_ctrl_delayed <= 1'b1; 
        end else begin
            if (cnt_ctrl_delayed && !cnt_ctrl) begin
                done_reg <= 1'b1;
            end else begin
                done_reg <= 1'b0;
            end
            cnt_ctrl_delayed <= cnt_ctrl;
        end
    end


    assign done = done_reg;

    always @(posedge cnt_in or negedge rst) begin
        if (!rst) begin
            cnt_out <= 32'd0;
        end else if (clear) begin
            cnt_out <= 32'd0;
        end else if (cnt_ctrl) begin
            cnt_out <= cnt_out + 1'd1;
        end else begin
            cnt_out <= cnt_out ;
        end
    end

endmodule



// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/29 14:50:53
// Design Name:
// Module Name: PUF128
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

//`define WIDTH  256
`include "header.sv"

module PUF128(
    input clk,
    input rst,
    input enable,             //PUF start
    input mode,              // 0: rng mode; 1: puf mode;
    input [127:0] challenge,
    output request,          //request a new challenge for rng mode
    input ready_challenge,   //new challenge ready
    output response_done,             //response generated
    output [`WIDTH - 1:0] response,
    output response_done_2bit,
    output [1:0] response2bit
);

parameter VOTE_NUM = 10;
// parameter CHALLENGE_NUM = 1000;

reg timer_enable;          //timer start to work
reg request_reg;
reg [8:0] shift_cnt;       // shift for 128 cycle
reg [5:0] vote_cnt;        //num of one response collect
reg [127:0] challenge_reg;
// wire response_done_2bit;   //PUF generate one bit response
// wire [1:0] response2bit;
reg [`WIDTH - 1:0] response_one;  //one 128bit response
reg one_resp_ready;        //one 128bit response ready to write to voter
reg vote_start;            //start to vote response
reg vote_clear;            //clear data in voter
//wire response_done;        //response after voting done
//reg [ `WIDTH - 1 :0] response_reg;  //final output response
reg [3:0] state;            // state reg for FSM

localparam                       IDLE =  0;            //wait for PUF start
localparam                       REQUEST  =  1;        //request new challenge for rng mode
localparam                       UPDATE = 2;           //challenge upated for rng mode
localparam                       RNG = 3;              //rng output gen
localparam                       SHIFT = 4;            //shift challenge (128)
localparam                       VOTE_STORE = 5;       //writ data to voter
localparam                       VOTE = 6;              //start vote
localparam                       ALL_DONE = 7;          //all tings done


PUF1bit puf_inst (
    .clk(clk),
    .rst(rst),
    .timer_enable(timer_enable),
    .challenge(challenge_reg),
    .response_done(response_done_2bit),
    .response(response2bit)
);

//vote
Voter #(.Threshold(5)) u_voter(
  .clk(clk),
  .rst(rst),
  .ready(one_resp_ready),
  .vote(vote_start),
  .clear(vote_clear),
  .done(response_done),
  .data_in(response_one),
  .data_out(response)
);

assign request = request_reg;
//assign response = response_reg;

always @(posedge clk or negedge rst) begin
    if (!rst) begin
        state <= IDLE;
        timer_enable <= 1'd0;
        request_reg <= 1'd0;
        shift_cnt <= 9'd0;
        vote_start <= 1'd0;
        vote_clear <= 1'd0;
        one_resp_ready <= 1'd0;
        vote_cnt <= 6'd0;
        response_one <= `WIDTH'd0;
        challenge_reg <= 128'd0;
    end else begin
        case(state)
            IDLE: begin
                if (enable) begin
                    if (!mode) begin              // jump to rng mode, request new challenge
                        state <= REQUEST;
                        timer_enable <= 1'd0;
                        request_reg <= 1'd0;
                        shift_cnt <= 9'd0;
                        vote_start <= 1'd0;
                        vote_clear <= 1'd0;
                        one_resp_ready <= 1'd0;
                        vote_cnt <= 6'd0;
                        response_one <= `WIDTH'd0;
                        challenge_reg <= 128'd0;
                    end else if (mode & (challenge != 0)) begin              // jump to puf mode, use challenge from primary input
                        state <= SHIFT;
                        timer_enable <= 1'd0;
                        request_reg <= 1'd0;
                        shift_cnt <= 9'd0;
                        vote_start <= 1'd0;
                        vote_clear <= 1'd0;
                        one_resp_ready <= 1'd0;
                        vote_cnt <= 6'd0;
                        response_one <= `WIDTH'd0;
                        challenge_reg <= challenge;
                    end
                end
            end
            REQUEST: begin
                if (enable & !mode) begin
                    state <= UPDATE;
                    timer_enable <= 1'd0;
                    request_reg <= 1'd1;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd1;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    challenge_reg <= 128'd0;
                end else begin
                    state <= ALL_DONE;
                    timer_enable <= 1'd0;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    challenge_reg <= 128'd0;
                end
            end
            UPDATE: begin
                if (ready_challenge) begin
                    state <= RNG;
                    timer_enable <= 1'd0;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    challenge_reg <= challenge;
                end
            end
            RNG: begin
                if (!response_done_2bit) begin
                    timer_enable <= 1'd1;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    state <= RNG;
                end else if (response_done_2bit) begin
                    timer_enable <= 1'd0;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    state <= REQUEST;
                end
            end
            SHIFT: begin
                if (shift_cnt < 9'd128) begin
                    if (!response_done_2bit) begin
                        timer_enable <= 1'd1;
                        challenge_reg <= challenge_reg;
                        request_reg <= 1'd0;
                        shift_cnt <= shift_cnt;
                        vote_start <= 1'd0;
                        vote_clear <= 1'd0;
                        one_resp_ready <= 1'd0;
                        vote_cnt <= vote_cnt;
                        response_one <= response_one;
                        state <= SHIFT;
                    end else if (response_done_2bit & timer_enable) begin
                        timer_enable <= 1'd0;
                        challenge_reg <= {challenge_reg[126:0], challenge_reg[127]};
                        request_reg <= 1'd0;
                        shift_cnt <= shift_cnt + 1'd1;
                        vote_start <= 1'd0;
                        vote_clear <= 1'd0;
                        one_resp_ready <= 1'd0;
                        vote_cnt <= vote_cnt;
                        response_one <= {response_one[`WIDTH-3:0],response2bit};
                        state <= SHIFT;
                    end else begin
                        timer_enable <= timer_enable;
                        challenge_reg <= challenge_reg;
                        request_reg <= 1'd0;
                        shift_cnt <= shift_cnt;
                        vote_start <= 1'd0;
                        vote_clear <= 1'd0;
                        one_resp_ready <= 1'd0;
                        vote_cnt <= vote_cnt;
                        response_one <= response_one;
                        state <= SHIFT;
                    end
                end else begin
                    timer_enable <= 1'd0;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd1;
                    vote_cnt <= vote_cnt;
                    response_one <= response_one;
                    state <= VOTE_STORE;
                end
            end
            VOTE_STORE: begin
                if (vote_cnt < VOTE_NUM -1 ) begin
                    timer_enable <= 1'd0;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= vote_cnt + 1'd1;
                    response_one <= `WIDTH'd0;
                    state <= SHIFT;
                end else if (vote_cnt >= VOTE_NUM -1 ) begin
                    timer_enable <= 1'd0;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd1;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    state <= VOTE;
                end
            end
            VOTE: begin
                if (response_done) begin
                    timer_enable <= 1'd0;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    state <= ALL_DONE;
                end else begin
                    timer_enable <= 1'd0;
                    challenge_reg <= challenge_reg;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd1;
                    vote_clear <= 1'd0;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    state <= VOTE;
                end
            end
            ALL_DONE: begin
                if (enable) begin
                    state <= ALL_DONE;
                    timer_enable <= 1'd0;
                    request_reg <= 1'd0;
                    shift_cnt <= 9'd0;
                    vote_start <= 1'd0;
                    vote_clear <= 1'd1;
                    one_resp_ready <= 1'd0;
                    vote_cnt <= 6'd0;
                    response_one <= `WIDTH'd0;
                    challenge_reg <= 128'd0;
                end else begin
                    state <= IDLE;
                end
            end

            default: state <= IDLE;
        endcase
    end
end

endmodule



// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/30 17:03:05
// Design Name:
// Module Name: PUF1bit
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
`include "header.sv"

module PUF1bit(
    input clk,
    input rst,
    input timer_enable,             //PUF start
    input [127:0] challenge,
    output response_done,             //response generated, can be sent form UART
    output [1:0] response
);

`ifdef SYNTHESIS_ZDR
// `define TEST
// `ifdef TEST
parameter NUM_LUTS = 5;
parameter  NUM_OSCILLATORS = 128;

wire [127:0]  mux_in_a;      //RO output to MUX
wire [127:0]  mux_in_b;
wire [127:0] dec_out_a;     //RO selected to work
wire [127:0] dec_out_b;
wire [6:0] dec_in_a;        //RO selected code(need to decode)
wire [6:0] dec_in_b;
wire [31:0] cnt_out_a;       // counter output
wire [31:0] cnt_out_b;
wire cnt_ctrl;              //timer output to control the counter
// (* keep="true" *) wire [639:0] ca;            //RO lines
// (* keep="true" *) wire [639:0] cb;
wire [127:0] ena;           //RO enable signle
wire [127:0] enb;
wire cnt_done, cnt_done_a, cnt_done_b;  //counter ready to read data
(* keep="true" *) wire mux_out_a, mux_out_b;

(* keep="true" *) wire [127:0] ro_a;
(* keep="true" *) wire [127:0] ro_b;

//wire [639:0] ca_test;            //RO lines
//wire [639:0] cb_test;

 genvar i;
  generate
    for (i=0; i < NUM_OSCILLATORS; i=i+1) begin: puf_a
    (* keep="true" *)  wire [NUM_LUTS-1:0] ca; 

      LUT3 #(.INIT(8'h7F)) LUTa_init (
        .O(ca[0]),
        .I0(ena[i]),
        .I1(rst),
        .I2(ca[NUM_LUTS-1])
      );

    //   assign #2 ca[0] = !(ena[i] & rst & ca[NUM_LUTS-1]);

      genvar j;
      for (j=1; j < NUM_LUTS; j=j+1) begin: LUT_chain
        LUT1 #(.INIT(2'h1)) LUT (
          .O(ca[j]),
          .I0(ca[j-1])
        );
      end

      LUT1 #(.INIT(2'h1)) LUTa_last (
        .O(ro_a[i]),
        .I0(ca[NUM_LUTS-3]) 
      );

      assign mux_in_a[i] = ro_a[i];
      assign ena[i] = dec_out_a[i];
    end
  endgenerate

genvar m;
  generate
    for (m=0; m < NUM_OSCILLATORS; m=m+1) begin: puf_b
    (* keep="true" *)  wire [NUM_LUTS-1:0] cb; 

      LUT3 #(.INIT(8'h7F)) LUTa_init (
        .O(cb[0]),
        .I0(enb[m]),
        .I1(rst),
        .I2(cb[NUM_LUTS-1])
      );
    //   assign #2 cb[0] = !(enb[m] & rst & cb[NUM_LUTS-1]);

      genvar n;
      for (n=1; n < NUM_LUTS; n=n+1) begin: LUT_chain
        LUT1 #(.INIT(2'h1)) LUT (
          .O(cb[n]),
          .I0(cb[n-1])
        );
      end

      LUT1 #(.INIT(2'h1)) LUTa_last (
        .O(ro_b[m]),
        .I0(cb[NUM_LUTS-3]) 
      );

      assign mux_in_b[m] = ro_b[m];
      assign enb[m] = dec_out_b[m];
    end
  endgenerate

// genvar i;
// generate
//   for (i=0; i < 128; i=i+1)
//   begin: puf_a
//      LUT3  #(.INIT(8'h7f)) LUTa0 (
//       .O(ca[0+5*i]),
//       .I0(ena[i]),
//       .I1(rst),
//       .I2(ca[4+5*i])
//      );
//      LUT1 #(.INIT(2'h1)) LUTa1(
//       .O(ca[1+5*i]),
//       .I0(ca[0+5*i])
//     );

//     LUT1 #(.INIT(2'h1)) LUTa2(
//         .O(ca[2+5*i]),
//         .I0(ca[1+5*i])
//     );

//     LUT1 #(.INIT(2'h1)) LUTa3(
//         .O(ca[3+5*i]),
//         .I0(ca[2+5*i])
//     );

//     LUT1 #(.INIT(2'h1)) LUTa4(
//         .O(ca[4+5*i]),
//         .I0(ca[3+5*i])
//     );

//     LUT1 #(.INIT(2'h1)) LUTa5(
//         .O(ro_a[i]),
//         .I0(ca[i*5+2])
//     );
//     assign mux_in_a[i] = ro_a[i];
//     assign ena[i] = dec_out_a[i];

//   end
// endgenerate

// genvar j;
// generate
//   for (j=0; j < 128; j=j+1)
//   begin: puf_b
//      LUT3  #(.INIT(8'h7f)) LUTb0 (
//       .O(cb[0+5*j]),
//       .I0(enb[j]),
//       .I1(rst),
//       .I2(cb[4+5*j])
//      );
//      LUT1 #(.INIT(2'h1)) LUTb1(
//       .O(cb[1+5*j]),
//       .I0(cb[0+5*j])
//     );

//     LUT1 #(.INIT(2'h1)) LUTb2(
//         .O(cb[2+5*j]),
//         .I0(cb[1+5*j])
//     );

//     LUT1 #(.INIT(2'h1)) LUTb3(
//         .O(cb[3+5*j]),
//         .I0(cb[2+5*j])
//     );

//     LUT1 #(.INIT(2'h1)) LUTb4(
//         .O(cb[4+5*j]),
//         .I0(cb[3+5*j])
//     );

//     LUT1 #(.INIT(2'h1)) LUTb5(
//         .O(ro_b[j]),
//         .I0(cb[j*5+2])
//     );
//    assign mux_in_b[j] = ro_b[j];
//    assign enb[j] = dec_out_b[j];

//   end
// endgenerate

//zdr: can be improved
assign dec_in_b = challenge[6:0];
assign dec_in_a = challenge[13:7];

PUFDec128 DecA(
    .i_Sel(dec_in_a),
    .o_Q(dec_out_a)
);

PUFDec128 DecB(
    .i_Sel(dec_in_b),
    .o_Q(dec_out_b)
);

PUFMux128 MuxA(
    .i_D(mux_in_a),
    .i_Sel(dec_in_a),
    .o_Q(mux_out_a)
);

PUFMux128 MuxB(
    .i_D(mux_in_b),
    .i_Sel(dec_in_b),
    .o_Q(mux_out_b)
);

Timer #(.target(5'd15)) u_timer(
    .rst(rst),
    .clk(clk),
    .enable(timer_enable),
    .ctrl(cnt_ctrl)
);

Counter CounterA(
    .cnt_in(mux_out_a),
    .clk(clk),
    .rst(rst),
    .cnt_out(cnt_out_a),
    .cnt_ctrl(cnt_ctrl),
    .done(cnt_done_a),
    .clear(cnt_clear)
);

Counter CounterB(
    .cnt_in(mux_out_b),
    .clk(clk),
    .rst(rst),
    .cnt_out(cnt_out_b),
    .cnt_ctrl(cnt_ctrl),
    .done(cnt_done_b),
    .clear(cnt_clear)
);

assign cnt_done = cnt_done_a && cnt_done_b;

Comp u_comp(
    .clk(clk),
    .rst(rst),
    .num1(cnt_out_a),
    .num2(cnt_out_b),
    .comp_en(cnt_done),
    .done(response_done),
    .result(response)
);

Timer #(.target(2)) u_cnt_clear(
    .rst(rst),
    .clk(clk),
    .enable(response_done),
    .ctrl(cnt_clear)
);

`else

localparam M = 15; // 定义LFSR运行周期的数量，根据需要修改
reg [127:0] lfsr; // 128位线性反馈移位寄存器
reg [3:0] done_counter; // 完成后的倒计时计数器
reg [7:0] run_counter; // LFSR运行计数器

reg [1:0] response_reg;
reg response_done_reg;

assign response = response_reg;
assign response_done = response_done_reg;

always @(posedge clk or negedge rst) begin
    if (!rst) begin
        lfsr <= 0;
        response_reg <= 0;
        response_done_reg <= 0;
        done_counter <= 0;
        run_counter <= 0;
    end else if (timer_enable) begin
        if (run_counter == 0) begin
            lfsr <= challenge;
            run_counter <= run_counter + 1;
        end  else if (run_counter < M) begin
            lfsr <= {lfsr[0]^lfsr[22]^lfsr[36]^lfsr[49]^lfsr[88],lfsr[37]^lfsr[85]^lfsr[96]^lfsr[108]^lfsr[122],lfsr[127:2]};
            run_counter <= run_counter + 1;
        end else  if (run_counter == M) begin
            response_reg <= lfsr[127:126]; // 取LFSR的高两位作为response
            response_done_reg <= 1; // 标记响应完成
            run_counter <= run_counter + 1; // 防止重复进入此条件分支
        end
    end else if (response_done_reg) begin
        if (done_counter < 2) begin
            done_counter <= done_counter + 1;
        end else begin
            response_done_reg <= 0; // 2个周期后将response_done置低
            done_counter <= 0; // 重置计数器
        end
    end else begin
        // 当timer_enable为低且response_done为低时，复位计数器
        run_counter <= 0;
        done_counter <= 0;
    end
end


`endif

endmodule



`include "header.sv"

module PUF_core (
    input clk,
    input rst_n,
    input enable,
    input mode,   // 0: rng mode; 1: puf mode
    input ready_challenge,  //new challenge ready
    input [127:0] challenge, // a 128bit challenge
    output response_done,
    output response_valid,
    output [`WIDTH - 1:0] response,
    output response_valid_re,
    output [`WIDTH/32 -1:0]response_re,
    output response_done_2bit_re,
    output response_done_2bit,
    output [1:0] response2bit,
    output [3:0] rng4bit,
    output rng4bit_done,
    output rng_mode,
    input es_rng_req
);

wire request;
wire [127:0] challenge_rng, challenge_puf;
wire ready_challenge_rng, ready_challenge_puf;
wire response_done_2bit_puf;
wire [1:0] response2bit_puf;

reg [3:0] rng4bit_reg;
reg rng4bit_done_reg;

assign challenge_puf = mode ? challenge : challenge_rng;
assign ready_challenge_puf = mode ? ready_challenge : ready_challenge_rng;

assign response_done_2bit = mode ? 0 : response_done_2bit_puf;
assign response2bit = mode ? 0 : response2bit_puf;

assign response_valid_re = 1;
assign response_re = {8{response_done}};
assign response_done_2bit_re = 1;
PUF128 #(.VOTE_NUM(10)) puf_128 (
    .clk(clk),
    .rst(rst_n),
    .enable(enable),
    .mode(mode),
    .challenge(challenge_puf),
    .ready_challenge(ready_challenge_puf),
    .response_done(response_done),
    .response(response),
    .request(request),
    .response_done_2bit(response_done_2bit_puf),
    .response2bit(response2bit_puf)
);

rng_puf #(.Challenge_repeat(1)) u_rng(
  .clk(clk),                // Clock input
  .request(request),        // Request input
  .rst(rst_n),                // Reset input
  .ready_challenge(ready_challenge_rng),  // Ready output
  .challenge(challenge_rng)     // Challenge output
);

AP0BP1 u_AP0BP1(
  .clk   (clk   ),
  .rst_n (rst_n ),
  .A     (ready_challenge),
  .B     (response_done),
  .C     (response_valid)
);

assign rng_mode = mode;

// Internal signals
reg [1:0] counter; // 2-bit counter to count the number of times response2bit_puf is received
reg response_done_2bit_puf_d; // Delayed version of response_done_2bit_puf for edge detection

// Edge detection for response_done_2bit_puf
wire response_done_2bit_puf_rising;
assign response_done_2bit_puf_rising = response_done_2bit_puf & ~response_done_2bit_puf_d;

assign rng4bit = es_rng_req ? rng4bit_reg : 0;
assign rng4bit_done = rng4bit_done_reg & es_rng_req;

// Sequential logic for updating rng4bit_reg and rng4bit_reg_done
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        // Reset state
        rng4bit_reg <= 4'b0000;
        rng4bit_done_reg <= 1'b0;
        counter <= 2'b00;
        response_done_2bit_puf_d <= 1'b0;
    end else begin
        // Default state
        rng4bit_done_reg <= 1'b0; // Clear rng4bit_done_reg flag every cycle
        response_done_2bit_puf_d <= response_done_2bit_puf; // Update the delayed version

        // Check if there is a rising edge on response_done_2bit_puf
        if (response_done_2bit_puf_rising) begin
            // Fill rng4bit_reg on successive rising edges
            if (counter < 2'b10) begin
                // Shift the response into rng4bit_reg
                rng4bit_reg <= {rng4bit_reg[1:0], response2bit_puf};
                // Increment the counter
                counter <= counter + 1;
            end
            // Check if rng4bit_reg is filled
            if (counter == 2'b01) begin // Counter was 0 before, now it's 1, so rng4bit_reg is full
                rng4bit_done_reg <= 1'b1; // Set rng4bit_done_reg high for one cycle
                counter <= 2'b00; // Reset the counter
                rng4bit_reg <= rng4bit_reg ^ challenge_rng[127:124];
            end
        end
    end
end

endmodule



// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/29 15:38:12
// Design Name:
// Module Name: PUFDec128
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module PUFDec128(
    input [6:0] i_Sel,
    output reg [127:0] o_Q
);

generate
    genvar i;
    for(i=0; i<128; i=i+1) begin
        always @ (i_Sel) begin
            if(i == i_Sel) begin
                o_Q[i] = 1'b1;
            end else begin
                o_Q[i] = 1'b0;
            end
        end
    end
endgenerate

endmodule




module PUFMux128 (
input [127:0] i_D,
input [6:0] i_Sel,
output reg o_Q
);

always @(*) begin
	case(i_Sel)
		7'b0000000: o_Q = i_D[0];
		7'b0000001: o_Q = i_D[1];
		7'b0000010: o_Q = i_D[2];
		7'b0000011: o_Q = i_D[3];
		7'b0000100: o_Q = i_D[4];
		7'b0000101: o_Q = i_D[5];
		7'b0000110: o_Q = i_D[6];
		7'b0000111: o_Q = i_D[7];
		7'b0001000: o_Q = i_D[8];
		7'b0001001: o_Q = i_D[9];
		7'b0001010: o_Q = i_D[10];
		7'b0001011: o_Q = i_D[11];
		7'b0001100: o_Q = i_D[12];
		7'b0001101: o_Q = i_D[13];
		7'b0001110: o_Q = i_D[14];
		7'b0001111: o_Q = i_D[15];
		7'b0010000: o_Q = i_D[16];
		7'b0010001: o_Q = i_D[17];
		7'b0010010: o_Q = i_D[18];
		7'b0010011: o_Q = i_D[19];
		7'b0010100: o_Q = i_D[20];
		7'b0010101: o_Q = i_D[21];
		7'b0010110: o_Q = i_D[22];
		7'b0010111: o_Q = i_D[23];
		7'b0011000: o_Q = i_D[24];
		7'b0011001: o_Q = i_D[25];
		7'b0011010: o_Q = i_D[26];
		7'b0011011: o_Q = i_D[27];
		7'b0011100: o_Q = i_D[28];
		7'b0011101: o_Q = i_D[29];
		7'b0011110: o_Q = i_D[30];
		7'b0011111: o_Q = i_D[31];
		7'b0100000: o_Q = i_D[32];
		7'b0100001: o_Q = i_D[33];
		7'b0100010: o_Q = i_D[34];
		7'b0100011: o_Q = i_D[35];
		7'b0100100: o_Q = i_D[36];
		7'b0100101: o_Q = i_D[37];
		7'b0100110: o_Q = i_D[38];
		7'b0100111: o_Q = i_D[39];
		7'b0101000: o_Q = i_D[40];
		7'b0101001: o_Q = i_D[41];
		7'b0101010: o_Q = i_D[42];
		7'b0101011: o_Q = i_D[43];
		7'b0101100: o_Q = i_D[44];
		7'b0101101: o_Q = i_D[45];
		7'b0101110: o_Q = i_D[46];
		7'b0101111: o_Q = i_D[47];
		7'b0110000: o_Q = i_D[48];
		7'b0110001: o_Q = i_D[49];
		7'b0110010: o_Q = i_D[50];
		7'b0110011: o_Q = i_D[51];
		7'b0110100: o_Q = i_D[52];
		7'b0110101: o_Q = i_D[53];
		7'b0110110: o_Q = i_D[54];
		7'b0110111: o_Q = i_D[55];
		7'b0111000: o_Q = i_D[56];
		7'b0111001: o_Q = i_D[57];
		7'b0111010: o_Q = i_D[58];
		7'b0111011: o_Q = i_D[59];
		7'b0111100: o_Q = i_D[60];
		7'b0111101: o_Q = i_D[61];
		7'b0111110: o_Q = i_D[62];
		7'b0111111: o_Q = i_D[63];
		7'b1000000: o_Q = i_D[64];
		7'b1000001: o_Q = i_D[65];
		7'b1000010: o_Q = i_D[66];
		7'b1000011: o_Q = i_D[67];
		7'b1000100: o_Q = i_D[68];
		7'b1000101: o_Q = i_D[69];
		7'b1000110: o_Q = i_D[70];
		7'b1000111: o_Q = i_D[71];
		7'b1001000: o_Q = i_D[72];
		7'b1001001: o_Q = i_D[73];
		7'b1001010: o_Q = i_D[74];
		7'b1001011: o_Q = i_D[75];
		7'b1001100: o_Q = i_D[76];
		7'b1001101: o_Q = i_D[77];
		7'b1001110: o_Q = i_D[78];
		7'b1001111: o_Q = i_D[79];
		7'b1010000: o_Q = i_D[80];
		7'b1010001: o_Q = i_D[81];
		7'b1010010: o_Q = i_D[82];
		7'b1010011: o_Q = i_D[83];
		7'b1010100: o_Q = i_D[84];
		7'b1010101: o_Q = i_D[85];
		7'b1010110: o_Q = i_D[86];
		7'b1010111: o_Q = i_D[87];
		7'b1011000: o_Q = i_D[88];
		7'b1011001: o_Q = i_D[89];
		7'b1011010: o_Q = i_D[90];
		7'b1011011: o_Q = i_D[91];
		7'b1011100: o_Q = i_D[92];
		7'b1011101: o_Q = i_D[93];
		7'b1011110: o_Q = i_D[94];
		7'b1011111: o_Q = i_D[95];
		7'b1100000: o_Q = i_D[96];
		7'b1100001: o_Q = i_D[97];
		7'b1100010: o_Q = i_D[98];
		7'b1100011: o_Q = i_D[99];
		7'b1100100: o_Q = i_D[100];
		7'b1100101: o_Q = i_D[101];
		7'b1100110: o_Q = i_D[102];
		7'b1100111: o_Q = i_D[103];
		7'b1101000: o_Q = i_D[104];
		7'b1101001: o_Q = i_D[105];
		7'b1101010: o_Q = i_D[106];
		7'b1101011: o_Q = i_D[107];
		7'b1101100: o_Q = i_D[108];
		7'b1101101: o_Q = i_D[109];
		7'b1101110: o_Q = i_D[110];
		7'b1101111: o_Q = i_D[111];
		7'b1110000: o_Q = i_D[112];
		7'b1110001: o_Q = i_D[113];
		7'b1110010: o_Q = i_D[114];
		7'b1110011: o_Q = i_D[115];
		7'b1110100: o_Q = i_D[116];
		7'b1110101: o_Q = i_D[117];
		7'b1110110: o_Q = i_D[118];
		7'b1110111: o_Q = i_D[119];
		7'b1111000: o_Q = i_D[120];
		7'b1111001: o_Q = i_D[121];
		7'b1111010: o_Q = i_D[122];
		7'b1111011: o_Q = i_D[123];
		7'b1111100: o_Q = i_D[124];
		7'b1111101: o_Q = i_D[125];
		7'b1111110: o_Q = i_D[126];
		default: o_Q = i_D[127];
	endcase
end

endmodule



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package puf_reg_pkg;

  // Param list
  parameter int NumRegs_challenge = 4;
  parameter int NumRegs_response = 8;

  // Address widths within the block
  parameter int BlockAw = 6;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } enable_puf;
    struct packed {
      logic        q;
      logic        qe;
    } mode_puf;
    struct packed {
      logic        q;
      logic        qe;
    } ready_cha;
  } puf_reg2hw_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } response_valid_bit;
    struct packed {
      logic        q;
    } response_done_2bit;
  } puf_reg2hw_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } puf_reg2hw_challenge_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } puf_reg2hw_response_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } enable_puf;
    struct packed {
      logic        d;
      logic        de;
    } mode_puf;
    struct packed {
      logic        d;
      logic        de;
    } ready_cha;
  } puf_hw2reg_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } response_valid_bit;
    struct packed {
      logic        d;
      logic        de;
    } response_done_2bit;
  } puf_hw2reg_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } puf_hw2reg_challenge_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } puf_hw2reg_response_mreg_t;

  // Register -> HW type
  typedef struct packed {
    puf_reg2hw_ctrl_signals_reg_t ctrl_signals; // [395:390]
    puf_reg2hw_state_signals_reg_t state_signals; // [389:388]
    puf_reg2hw_challenge_mreg_t [3:0] challenge; // [387:256]
    puf_reg2hw_response_mreg_t [7:0] response; // [255:0]
  } puf_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    puf_hw2reg_ctrl_signals_reg_t ctrl_signals; // [405:400]
    puf_hw2reg_state_signals_reg_t state_signals; // [399:396]
    puf_hw2reg_challenge_mreg_t [3:0] challenge; // [395:264]
    puf_hw2reg_response_mreg_t [7:0] response; // [263:0]
  } puf_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] PUF_CTRL_SIGNALS_OFFSET = 6'h 0;
  parameter logic [BlockAw-1:0] PUF_STATE_SIGNALS_OFFSET = 6'h 4;
  parameter logic [BlockAw-1:0] PUF_CHALLENGE_0_OFFSET = 6'h 8;
  parameter logic [BlockAw-1:0] PUF_CHALLENGE_1_OFFSET = 6'h c;
  parameter logic [BlockAw-1:0] PUF_CHALLENGE_2_OFFSET = 6'h 10;
  parameter logic [BlockAw-1:0] PUF_CHALLENGE_3_OFFSET = 6'h 14;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_0_OFFSET = 6'h 18;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_1_OFFSET = 6'h 1c;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_2_OFFSET = 6'h 20;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_3_OFFSET = 6'h 24;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_4_OFFSET = 6'h 28;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_5_OFFSET = 6'h 2c;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_6_OFFSET = 6'h 30;
  parameter logic [BlockAw-1:0] PUF_RESPONSE_7_OFFSET = 6'h 34;

  // Register index
  typedef enum int {
    PUF_CTRL_SIGNALS,
    PUF_STATE_SIGNALS,
    PUF_CHALLENGE_0,
    PUF_CHALLENGE_1,
    PUF_CHALLENGE_2,
    PUF_CHALLENGE_3,
    PUF_RESPONSE_0,
    PUF_RESPONSE_1,
    PUF_RESPONSE_2,
    PUF_RESPONSE_3,
    PUF_RESPONSE_4,
    PUF_RESPONSE_5,
    PUF_RESPONSE_6,
    PUF_RESPONSE_7
  } puf_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] PUF_PERMIT [14] = '{
    4'b 0001, // index[ 0] PUF_CTRL_SIGNALS
    4'b 0001, // index[ 1] PUF_STATE_SIGNALS
    4'b 1111, // index[ 2] PUF_CHALLENGE_0
    4'b 1111, // index[ 3] PUF_CHALLENGE_1
    4'b 1111, // index[ 4] PUF_CHALLENGE_2
    4'b 1111, // index[ 5] PUF_CHALLENGE_3
    4'b 1111, // index[ 6] PUF_RESPONSE_0
    4'b 1111, // index[ 7] PUF_RESPONSE_1
    4'b 1111, // index[ 8] PUF_RESPONSE_2
    4'b 1111, // index[ 9] PUF_RESPONSE_3
    4'b 1111, // index[10] PUF_RESPONSE_4
    4'b 1111, // index[11] PUF_RESPONSE_5
    4'b 1111, // index[12] PUF_RESPONSE_6
    4'b 1111  // index[13] PUF_RESPONSE_7
  };

endpackage



// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module puf_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output puf_reg_pkg::puf_reg2hw_t reg2hw, // Write
  input  puf_reg_pkg::puf_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import puf_reg_pkg::* ;

  localparam int AW = 6;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [13:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(14)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic ctrl_signals_we;
  logic ctrl_signals_enable_puf_qs;
  logic ctrl_signals_enable_puf_wd;
  logic ctrl_signals_mode_puf_qs;
  logic ctrl_signals_mode_puf_wd;
  logic ctrl_signals_ready_cha_qs;
  logic ctrl_signals_ready_cha_wd;
  logic state_signals_response_valid_bit_qs;
  logic state_signals_response_done_2bit_qs;
  logic challenge_0_we;
  logic [31:0] challenge_0_qs;
  logic [31:0] challenge_0_wd;
  logic challenge_1_we;
  logic [31:0] challenge_1_qs;
  logic [31:0] challenge_1_wd;
  logic challenge_2_we;
  logic [31:0] challenge_2_qs;
  logic [31:0] challenge_2_wd;
  logic challenge_3_we;
  logic [31:0] challenge_3_qs;
  logic [31:0] challenge_3_wd;
  logic [31:0] response_0_qs;
  logic [31:0] response_1_qs;
  logic [31:0] response_2_qs;
  logic [31:0] response_3_qs;
  logic [31:0] response_4_qs;
  logic [31:0] response_5_qs;
  logic [31:0] response_6_qs;
  logic [31:0] response_7_qs;

  // Register instances
  // R[ctrl_signals]: V(False)
  logic ctrl_signals_qe;
  logic [2:0] ctrl_signals_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_ctrl_signals0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&ctrl_signals_flds_we),
    .q_o(ctrl_signals_qe)
  );
  //   F[enable_puf]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_enable_puf (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_enable_puf_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.enable_puf.de),
    .d      (hw2reg.ctrl_signals.enable_puf.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[0]),
    .q      (reg2hw.ctrl_signals.enable_puf.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_enable_puf_qs)
  );
  assign reg2hw.ctrl_signals.enable_puf.qe = ctrl_signals_qe;

  //   F[mode_puf]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_mode_puf (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_mode_puf_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.mode_puf.de),
    .d      (hw2reg.ctrl_signals.mode_puf.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[1]),
    .q      (reg2hw.ctrl_signals.mode_puf.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_mode_puf_qs)
  );
  assign reg2hw.ctrl_signals.mode_puf.qe = ctrl_signals_qe;

  //   F[ready_cha]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_ready_cha (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_ready_cha_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.ready_cha.de),
    .d      (hw2reg.ctrl_signals.ready_cha.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[2]),
    .q      (reg2hw.ctrl_signals.ready_cha.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_ready_cha_qs)
  );
  assign reg2hw.ctrl_signals.ready_cha.qe = ctrl_signals_qe;


  // R[state_signals]: V(False)
  //   F[response_valid_bit]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_response_valid_bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.response_valid_bit.de),
    .d      (hw2reg.state_signals.response_valid_bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.response_valid_bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_response_valid_bit_qs)
  );

  //   F[response_done_2bit]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_response_done_2bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.response_done_2bit.de),
    .d      (hw2reg.state_signals.response_done_2bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.response_done_2bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_response_done_2bit_qs)
  );


  // Subregister 0 of Multireg challenge
  // R[challenge_0]: V(False)
  logic challenge_0_qe;
  logic [0:0] challenge_0_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_challenge0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&challenge_0_flds_we),
    .q_o(challenge_0_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_challenge_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (challenge_0_we),
    .wd     (challenge_0_wd),

    // from internal hardware
    .de     (hw2reg.challenge[0].de),
    .d      (hw2reg.challenge[0].d),

    // to internal hardware
    .qe     (challenge_0_flds_we[0]),
    .q      (reg2hw.challenge[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (challenge_0_qs)
  );
  assign reg2hw.challenge[0].qe = challenge_0_qe;


  // Subregister 1 of Multireg challenge
  // R[challenge_1]: V(False)
  logic challenge_1_qe;
  logic [0:0] challenge_1_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_challenge1_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&challenge_1_flds_we),
    .q_o(challenge_1_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_challenge_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (challenge_1_we),
    .wd     (challenge_1_wd),

    // from internal hardware
    .de     (hw2reg.challenge[1].de),
    .d      (hw2reg.challenge[1].d),

    // to internal hardware
    .qe     (challenge_1_flds_we[0]),
    .q      (reg2hw.challenge[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (challenge_1_qs)
  );
  assign reg2hw.challenge[1].qe = challenge_1_qe;


  // Subregister 2 of Multireg challenge
  // R[challenge_2]: V(False)
  logic challenge_2_qe;
  logic [0:0] challenge_2_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_challenge2_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&challenge_2_flds_we),
    .q_o(challenge_2_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_challenge_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (challenge_2_we),
    .wd     (challenge_2_wd),

    // from internal hardware
    .de     (hw2reg.challenge[2].de),
    .d      (hw2reg.challenge[2].d),

    // to internal hardware
    .qe     (challenge_2_flds_we[0]),
    .q      (reg2hw.challenge[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (challenge_2_qs)
  );
  assign reg2hw.challenge[2].qe = challenge_2_qe;


  // Subregister 3 of Multireg challenge
  // R[challenge_3]: V(False)
  logic challenge_3_qe;
  logic [0:0] challenge_3_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_challenge3_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&challenge_3_flds_we),
    .q_o(challenge_3_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_challenge_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (challenge_3_we),
    .wd     (challenge_3_wd),

    // from internal hardware
    .de     (hw2reg.challenge[3].de),
    .d      (hw2reg.challenge[3].d),

    // to internal hardware
    .qe     (challenge_3_flds_we[0]),
    .q      (reg2hw.challenge[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (challenge_3_qs)
  );
  assign reg2hw.challenge[3].qe = challenge_3_qe;


  // Subregister 0 of Multireg response
  // R[response_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[0].de),
    .d      (hw2reg.response[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_0_qs)
  );


  // Subregister 1 of Multireg response
  // R[response_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[1].de),
    .d      (hw2reg.response[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_1_qs)
  );


  // Subregister 2 of Multireg response
  // R[response_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[2].de),
    .d      (hw2reg.response[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_2_qs)
  );


  // Subregister 3 of Multireg response
  // R[response_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[3].de),
    .d      (hw2reg.response[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_3_qs)
  );


  // Subregister 4 of Multireg response
  // R[response_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[4].de),
    .d      (hw2reg.response[4].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_4_qs)
  );


  // Subregister 5 of Multireg response
  // R[response_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[5].de),
    .d      (hw2reg.response[5].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_5_qs)
  );


  // Subregister 6 of Multireg response
  // R[response_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[6].de),
    .d      (hw2reg.response[6].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_6_qs)
  );


  // Subregister 7 of Multireg response
  // R[response_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_response_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.response[7].de),
    .d      (hw2reg.response[7].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.response[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (response_7_qs)
  );



  logic [13:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == PUF_CTRL_SIGNALS_OFFSET);
    addr_hit[ 1] = (reg_addr == PUF_STATE_SIGNALS_OFFSET);
    addr_hit[ 2] = (reg_addr == PUF_CHALLENGE_0_OFFSET);
    addr_hit[ 3] = (reg_addr == PUF_CHALLENGE_1_OFFSET);
    addr_hit[ 4] = (reg_addr == PUF_CHALLENGE_2_OFFSET);
    addr_hit[ 5] = (reg_addr == PUF_CHALLENGE_3_OFFSET);
    addr_hit[ 6] = (reg_addr == PUF_RESPONSE_0_OFFSET);
    addr_hit[ 7] = (reg_addr == PUF_RESPONSE_1_OFFSET);
    addr_hit[ 8] = (reg_addr == PUF_RESPONSE_2_OFFSET);
    addr_hit[ 9] = (reg_addr == PUF_RESPONSE_3_OFFSET);
    addr_hit[10] = (reg_addr == PUF_RESPONSE_4_OFFSET);
    addr_hit[11] = (reg_addr == PUF_RESPONSE_5_OFFSET);
    addr_hit[12] = (reg_addr == PUF_RESPONSE_6_OFFSET);
    addr_hit[13] = (reg_addr == PUF_RESPONSE_7_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(PUF_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(PUF_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(PUF_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(PUF_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(PUF_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(PUF_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(PUF_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(PUF_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(PUF_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(PUF_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(PUF_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(PUF_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(PUF_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(PUF_PERMIT[13] & ~reg_be)))));
  end

  // Generate write-enables
  assign ctrl_signals_we = addr_hit[0] & reg_we & !reg_error;

  assign ctrl_signals_enable_puf_wd = reg_wdata[0];

  assign ctrl_signals_mode_puf_wd = reg_wdata[1];

  assign ctrl_signals_ready_cha_wd = reg_wdata[2];
  assign challenge_0_we = addr_hit[2] & reg_we & !reg_error;

  assign challenge_0_wd = reg_wdata[31:0];
  assign challenge_1_we = addr_hit[3] & reg_we & !reg_error;

  assign challenge_1_wd = reg_wdata[31:0];
  assign challenge_2_we = addr_hit[4] & reg_we & !reg_error;

  assign challenge_2_wd = reg_wdata[31:0];
  assign challenge_3_we = addr_hit[5] & reg_we & !reg_error;

  assign challenge_3_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = ctrl_signals_we;
    reg_we_check[1] = 1'b0;
    reg_we_check[2] = challenge_0_we;
    reg_we_check[3] = challenge_1_we;
    reg_we_check[4] = challenge_2_we;
    reg_we_check[5] = challenge_3_we;
    reg_we_check[6] = 1'b0;
    reg_we_check[7] = 1'b0;
    reg_we_check[8] = 1'b0;
    reg_we_check[9] = 1'b0;
    reg_we_check[10] = 1'b0;
    reg_we_check[11] = 1'b0;
    reg_we_check[12] = 1'b0;
    reg_we_check[13] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = ctrl_signals_enable_puf_qs;
        reg_rdata_next[1] = ctrl_signals_mode_puf_qs;
        reg_rdata_next[2] = ctrl_signals_ready_cha_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = state_signals_response_valid_bit_qs;
        reg_rdata_next[1] = state_signals_response_done_2bit_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = challenge_0_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = challenge_1_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = challenge_2_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = challenge_3_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = response_0_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = response_1_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = response_2_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = response_3_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = response_4_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = response_5_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = response_6_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = response_7_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule



`include "prim_assert.sv"

module puf
  import puf_reg_pkg::*;
(
  input  logic                                      clk_i,
  input  logic                                      rst_ni,

  output [3:0] rng4bit,
  output rng4bit_done,
  output rng_mode,
  input es_rng_req,

  // Bus interface
  input  tlul_pkg::tl_h2d_t                         tl_i,
  output tlul_pkg::tl_d2h_t                         tl_o
);

  puf_reg2hw_t               reg2hw;
  puf_hw2reg_t               hw2reg;
  //wire                       ready_out;

puf_reg_top  u_puf_reg_top (
    .clk_i                             ( clk_i  ),
    .rst_ni                            ( rst_ni ),
    .tl_i                              ( tl_i   ),
    .hw2reg                            ( hw2reg ),
    .devmode_i                         ( 1'b1   ),

    .tl_o                              ( tl_o   ),
    .reg2hw                            ( reg2hw ),
    .intg_err_o                        ( )
);

assign hw2reg.ctrl_signals.mode_puf.de = 1'd0;
assign hw2reg.ctrl_signals.enable_puf.de = 1'd0;
assign hw2reg.ctrl_signals.ready_cha.de = 1'd0;
assign hw2reg.challenge[0].de = 1'd0;
assign hw2reg.challenge[1].de = 1'd0;
assign hw2reg.challenge[2].de = 1'd0;
assign hw2reg.challenge[3].de = 1'd0;


PUF_core  u_PUF_core (
    .clk                     ( clk_i  ),
    .rst_n                   ( rst_ni ),
    .enable                  ( reg2hw.ctrl_signals.enable_puf.q ),
    .mode                    ( reg2hw.ctrl_signals.mode_puf.q ),
    .ready_challenge         ( reg2hw.ctrl_signals.ready_cha.q ),
    .challenge               ( {reg2hw.challenge[3].q,reg2hw.challenge[2].q,reg2hw.challenge[1].q,reg2hw.challenge[0].q} ),

    .response_done           (  ),//暂时无用
    .response_valid          ( hw2reg.state_signals.response_valid_bit.d ),
    .response                ( {hw2reg.response[7].d,hw2reg.response[6].d,hw2reg.response[5].d,hw2reg.response[4].d,hw2reg.response[3].d,hw2reg.response[2].d,hw2reg.response[1].d,hw2reg.response[0].d} ),
    .response_valid_re       ( hw2reg.state_signals.response_valid_bit.de ),
    .response_re             ( {hw2reg.response[7].de,hw2reg.response[6].de,hw2reg.response[5].de,hw2reg.response[4].de,hw2reg.response[3].de,hw2reg.response[2].de,hw2reg.response[1].de,hw2reg.response[0].de} ),
    .response_done_2bit_re   ( hw2reg.state_signals.response_done_2bit.de ),
    .response_done_2bit      ( hw2reg.state_signals.response_done_2bit.d ),
    .response2bit            (  ),//暂时无用
    .rng4bit                 ( rng4bit ),
    .rng4bit_done            ( rng4bit_done ),
    .rng_mode                ( rng_mode ),
    .es_rng_req              ( es_rng_req )
);

endmodule



// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/29 15:45:14
// Design Name:
// Module Name: rng
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module rng_puf(
    input clk,
    input request,
    input rst,
    output ready_challenge,
    output [127:0] challenge
);

parameter Challenge_repeat = 2;
//parameter initial_seed = 128'hC5141C0383F09022C512E99C9A2A50A4;
parameter initial_seed = 128'hC9F99D6C9F99D6C9F99D6C9F99D6C9F;

reg [127:0] seed;
reg ready_challenge_reg;

assign challenge = seed;

assign ready_challenge = ready_challenge_reg;

reg sig_delay;
reg out;

always @(posedge clk or negedge rst) begin
    if (!rst) begin
        out <= 0;
        sig_delay <= 0;
    end
    else begin
        sig_delay <= request;
        if (sig_delay == 0 && request == 1) begin
            out <= 1;
        end
        else begin
            out <= 0;
        end
    end
end

reg [5:0] request_cnt;

always @(posedge clk or negedge rst) begin
    if (!rst) begin
        seed <= initial_seed;
        ready_challenge_reg <= 1'd0;
        request_cnt <= 6'd0;
    end else if(out & request_cnt == Challenge_repeat-1) begin
        //seed[0] <= ~(seed[127] ^ seed[125] ^ seed[100] ^ seed[98]);
        //seed <= {seed[126:0],seed[0]};
        seed <= {seed[0]^seed[63]^seed[96]^seed[127],seed[127:1]};
        ready_challenge_reg <= 1'd1;
        request_cnt <= 6'd0;
    end else if (out) begin
        seed <= seed;
        ready_challenge_reg <= 1'd1;
        request_cnt <= request_cnt + 1'd1;
    end
    else begin
        seed <= seed;
        ready_challenge_reg <= 1'd0;
        request_cnt <= request_cnt;
     end
end

endmodule



// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/29 16:58:55
// Design Name:
// Module Name: Timer
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Timer(
    input clk,
    input rst,
    input enable,
    output reg ctrl
);

parameter [5:0] target = 5'd15;
reg [31:0] count;

//reg sig_delay;
//reg out;

//always @(posedge clk or negedge rst) begin
//    if (!rst) begin
//        out <= 0;
//        sig_delay <= 0;
//    end
//    else begin
//        sig_delay <= enable;
//        if (sig_delay == 0 && enable == 1) begin
//            out <= 1;
//        end
//        else begin
//            out <= 0;
//        end
//    end
//end

always @(posedge clk or negedge rst) begin
    if (!rst) begin
        count <= 31'd0;
        ctrl <= 0;
    end else if (enable) begin
        if (count < target) begin
            count <= count + 1;
            ctrl <= 1;
        end else begin
            ctrl <= 0;
            count <= count;
        end
    end else if (!enable) begin
        ctrl <= 0;
        count <= 31'd0;
    end
end

endmodule



// `timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2023/03/30 11:13:19
// Design Name:
// Module Name: Vote
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

`include "header.sv"

module Voter(
  input wire clk,
  input wire rst,
  input wire ready,
  input wire vote,
  input wire clear,
  output wire done,
  input wire [`WIDTH-1:0] data_in,
  output reg [`WIDTH-1:0] data_out
);

parameter  Threshold = 5; // ��ֵ

//reg [127:0] data_out_reg;
reg [5:0] sum [0:`WIDTH-1];
reg [`WIDTH-1:0] done_reg;

genvar i;
generate
  for (i = 0; i < `WIDTH; i = i + 1) begin : adder
    always@(posedge clk or negedge rst) begin
        if(!rst) begin
            sum[i] <= 0;
            data_out[i] <= 0;
            done_reg[i] <= 1'd0;
        end else if (ready) begin
            sum[i] <= data_in[i] + sum[i];
            data_out[i] <= 0;
            done_reg[i] <= 1'd0;
        end else if (vote) begin
            if ( sum[i] >= Threshold ) begin
                data_out[i] <= 1;
                done_reg[i] <= 1'd1;
            end else begin
                data_out[i] <= 0;
                done_reg[i] <= 1'd1;
            end
        end else if (clear) begin
            sum[i] <= 0;
            data_out[i] <= 0;
            done_reg[i] <= 1'd0;
        end else begin
            sum[i] <= sum[i];
            data_out[i] <= data_out[i];
            done_reg[i] <= done_reg[i];
        end
      end
    end
assign done = & done_reg;

endgenerate

//assign data_out = data_out_reg;

endmodule



// -------------------------------------------------------------------------
//Reed-Solomon decoder
//Copyright (C) Wed May 22 10:06:57 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module rsdec(x, error, with_error, enable, valid, k, clk, clrn);
	input enable, clk, clrn;
	input [7:0] k, x;
	output [7:0] error;
	wire [7:0] error;
	output with_error, valid;
	reg with_error, valid;

	wire [7:0] s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31;
	wire [7:0] lambda, omega, alpha;
	reg [5:0] count;
	reg [32:0] phase;
	wire [7:0] D0, D1, DI;
	reg [7:0] D, D2;
	reg [7:0] u, length0, length1, length2, length3;
	reg syn_enable, syn_init, syn_shift, berl_enable;
	reg chien_search, chien_load, shorten;

	always @ (chien_search or shorten)
		valid = chien_search & ~shorten;

	rsdec_syn x0 (s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, 
		u, syn_enable, syn_shift&phase[0], syn_init, clk, clrn);
	rsdec_berl x1 (lambda, omega,
		s0, s31, s30, s29, s28, s27, s26, s25, s24, s23, s22, s21, s20, s19, s18, s17, s16, s15, s14, s13, s12, s11, s10, s9, s8, s7, s6, s5, s4, s3, s2, s1, 
		D0, D2, count, phase[0], phase[32], berl_enable, clk, clrn);
	rsdec_chien x2 (error, alpha, lambda, omega,
		D1, DI, chien_search, chien_load, shorten, clk, clrn);
	inverse x3 (DI, D);

	always @ (posedge clk or negedge clrn)
	begin
		if (~clrn)
		begin
			syn_enable <= 0;
			syn_shift <= 0;
			berl_enable <= 0;
			chien_search <= 1;
			chien_load <= 0;
			length0 <= 0;
			length2 <= 255 - k;
			count <= -1;
			phase <= 1;
			u <= 0;
			shorten <= 1;
			syn_init <= 0;
		end
		else
		begin
			if (enable & ~syn_enable & ~syn_shift)
			begin
				syn_enable <= 1;
				syn_init <= 1;
			end
			if (syn_enable)
			begin
				length0 <= length1;
				syn_init <= 0;
				if (length1 == k)
				begin
					syn_enable <= 0;
					syn_shift <= 1;
					berl_enable <= 1;
				end
			end
			if (berl_enable & with_error)
			begin
				if (phase[0])
				begin
					count <= count + 1;
					if (count == 31)
					begin
						syn_shift <= 0;
						length0 <= 0;
						chien_load <= 1;
						length2 <= length0;
					end
				end
				phase <= {phase[31:0], phase[32]};
			end
			if (berl_enable & ~with_error)
				if (&count)
				begin
					syn_shift <= 0;
					length0 <= 0;
					berl_enable <= 0;
				end
				else
					phase <= {phase[31:0], phase[32]};
			if (chien_load & phase[32])
			begin
				berl_enable <= 0;
				chien_load <= 0;
				chien_search <= 1;
				count <= -1;
				phase <= 1;
			end
			if (chien_search)
			begin
				length2 <= length3;
				if (length3 == 0)
					chien_search <= 0;
			end
		if (enable) u <= x;
		if (shorten == 1 && length2 == 0)
			shorten <= 0;
		end

	end

	always @ (chien_search or D0 or D1)
		if (chien_search) D = D1;
		else D = D0;

	always @ (DI or alpha or chien_load)
		if (chien_load) D2 = alpha;
		else D2 = DI;

	always @ (length0) length1 = length0 + 1;
	always @ (length2) length3 = length2 - 1;
	always @ (syn_shift or s0 or s1 or s2 or s3 or s4 or s5 or s6 or s7 or s8 or s9 or s10 or s11 or s12 or s13 or s14 or s15 or s16 or s17 or s18 or s19 or s20 or s21 or s22 or s23 or s24 or s25 or s26 or s27 or s28 or s29 or s30 or s31)
		if (syn_shift && (s0 | s1 | s2 | s3 | s4 | s5 | s6 | s7 | s8 | s9 | s10 | s11 | s12 | s13 | s14 | s15 | s16 | s17 | s18 | s19 | s20 | s21 | s22 | s23 | s24 | s25 | s26 | s27 | s28 | s29 | s30 | s31)!= 0)
			with_error = 1;
		else with_error = 0;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package rs_decode_reg_pkg;

  // Param list
  parameter int NumRegs_encoded_data_in = 50;
  parameter int NumRegs_error_pos_out = 50;

  // Address widths within the block
  parameter int BlockAw = 9;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } decode_en;
    struct packed {
      logic        q;
      logic        qe;
    } clrn;
  } rs_decode_reg2hw_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } output_valid_bit;
    struct packed {
      logic        q;
    } ready_bit;
    struct packed {
      logic        q;
    } with_error_bit;
  } rs_decode_reg2hw_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } rs_decode_reg2hw_encoded_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } rs_decode_reg2hw_error_pos_out_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } decode_en;
    struct packed {
      logic        d;
      logic        de;
    } clrn;
  } rs_decode_hw2reg_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } output_valid_bit;
    struct packed {
      logic        d;
      logic        de;
    } ready_bit;
    struct packed {
      logic        d;
      logic        de;
    } with_error_bit;
  } rs_decode_hw2reg_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } rs_decode_hw2reg_encoded_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } rs_decode_hw2reg_error_pos_out_mreg_t;

  // Register -> HW type
  typedef struct packed {
    rs_decode_reg2hw_ctrl_signals_reg_t ctrl_signals; // [3256:3253]
    rs_decode_reg2hw_state_signals_reg_t state_signals; // [3252:3250]
    rs_decode_reg2hw_encoded_data_in_mreg_t [49:0] encoded_data_in; // [3249:1600]
    rs_decode_reg2hw_error_pos_out_mreg_t [49:0] error_pos_out; // [1599:0]
  } rs_decode_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    rs_decode_hw2reg_ctrl_signals_reg_t ctrl_signals; // [3309:3306]
    rs_decode_hw2reg_state_signals_reg_t state_signals; // [3305:3300]
    rs_decode_hw2reg_encoded_data_in_mreg_t [49:0] encoded_data_in; // [3299:1650]
    rs_decode_hw2reg_error_pos_out_mreg_t [49:0] error_pos_out; // [1649:0]
  } rs_decode_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] RS_DECODE_CTRL_SIGNALS_OFFSET = 9'h 0;
  parameter logic [BlockAw-1:0] RS_DECODE_STATE_SIGNALS_OFFSET = 9'h 4;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_0_OFFSET = 9'h 8;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_1_OFFSET = 9'h c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_2_OFFSET = 9'h 10;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_3_OFFSET = 9'h 14;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_4_OFFSET = 9'h 18;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_5_OFFSET = 9'h 1c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_6_OFFSET = 9'h 20;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_7_OFFSET = 9'h 24;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_8_OFFSET = 9'h 28;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_9_OFFSET = 9'h 2c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_10_OFFSET = 9'h 30;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_11_OFFSET = 9'h 34;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_12_OFFSET = 9'h 38;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_13_OFFSET = 9'h 3c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_14_OFFSET = 9'h 40;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_15_OFFSET = 9'h 44;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_16_OFFSET = 9'h 48;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_17_OFFSET = 9'h 4c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_18_OFFSET = 9'h 50;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_19_OFFSET = 9'h 54;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_20_OFFSET = 9'h 58;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_21_OFFSET = 9'h 5c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_22_OFFSET = 9'h 60;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_23_OFFSET = 9'h 64;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_24_OFFSET = 9'h 68;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_25_OFFSET = 9'h 6c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_26_OFFSET = 9'h 70;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_27_OFFSET = 9'h 74;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_28_OFFSET = 9'h 78;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_29_OFFSET = 9'h 7c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_30_OFFSET = 9'h 80;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_31_OFFSET = 9'h 84;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_32_OFFSET = 9'h 88;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_33_OFFSET = 9'h 8c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_34_OFFSET = 9'h 90;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_35_OFFSET = 9'h 94;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_36_OFFSET = 9'h 98;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_37_OFFSET = 9'h 9c;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_38_OFFSET = 9'h a0;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_39_OFFSET = 9'h a4;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_40_OFFSET = 9'h a8;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_41_OFFSET = 9'h ac;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_42_OFFSET = 9'h b0;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_43_OFFSET = 9'h b4;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_44_OFFSET = 9'h b8;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_45_OFFSET = 9'h bc;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_46_OFFSET = 9'h c0;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_47_OFFSET = 9'h c4;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_48_OFFSET = 9'h c8;
  parameter logic [BlockAw-1:0] RS_DECODE_ENCODED_DATA_IN_49_OFFSET = 9'h cc;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_0_OFFSET = 9'h d0;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_1_OFFSET = 9'h d4;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_2_OFFSET = 9'h d8;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_3_OFFSET = 9'h dc;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_4_OFFSET = 9'h e0;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_5_OFFSET = 9'h e4;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_6_OFFSET = 9'h e8;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_7_OFFSET = 9'h ec;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_8_OFFSET = 9'h f0;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_9_OFFSET = 9'h f4;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_10_OFFSET = 9'h f8;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_11_OFFSET = 9'h fc;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_12_OFFSET = 9'h 100;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_13_OFFSET = 9'h 104;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_14_OFFSET = 9'h 108;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_15_OFFSET = 9'h 10c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_16_OFFSET = 9'h 110;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_17_OFFSET = 9'h 114;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_18_OFFSET = 9'h 118;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_19_OFFSET = 9'h 11c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_20_OFFSET = 9'h 120;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_21_OFFSET = 9'h 124;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_22_OFFSET = 9'h 128;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_23_OFFSET = 9'h 12c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_24_OFFSET = 9'h 130;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_25_OFFSET = 9'h 134;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_26_OFFSET = 9'h 138;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_27_OFFSET = 9'h 13c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_28_OFFSET = 9'h 140;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_29_OFFSET = 9'h 144;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_30_OFFSET = 9'h 148;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_31_OFFSET = 9'h 14c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_32_OFFSET = 9'h 150;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_33_OFFSET = 9'h 154;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_34_OFFSET = 9'h 158;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_35_OFFSET = 9'h 15c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_36_OFFSET = 9'h 160;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_37_OFFSET = 9'h 164;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_38_OFFSET = 9'h 168;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_39_OFFSET = 9'h 16c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_40_OFFSET = 9'h 170;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_41_OFFSET = 9'h 174;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_42_OFFSET = 9'h 178;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_43_OFFSET = 9'h 17c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_44_OFFSET = 9'h 180;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_45_OFFSET = 9'h 184;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_46_OFFSET = 9'h 188;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_47_OFFSET = 9'h 18c;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_48_OFFSET = 9'h 190;
  parameter logic [BlockAw-1:0] RS_DECODE_ERROR_POS_OUT_49_OFFSET = 9'h 194;

  // Register index
  typedef enum int {
    RS_DECODE_CTRL_SIGNALS,
    RS_DECODE_STATE_SIGNALS,
    RS_DECODE_ENCODED_DATA_IN_0,
    RS_DECODE_ENCODED_DATA_IN_1,
    RS_DECODE_ENCODED_DATA_IN_2,
    RS_DECODE_ENCODED_DATA_IN_3,
    RS_DECODE_ENCODED_DATA_IN_4,
    RS_DECODE_ENCODED_DATA_IN_5,
    RS_DECODE_ENCODED_DATA_IN_6,
    RS_DECODE_ENCODED_DATA_IN_7,
    RS_DECODE_ENCODED_DATA_IN_8,
    RS_DECODE_ENCODED_DATA_IN_9,
    RS_DECODE_ENCODED_DATA_IN_10,
    RS_DECODE_ENCODED_DATA_IN_11,
    RS_DECODE_ENCODED_DATA_IN_12,
    RS_DECODE_ENCODED_DATA_IN_13,
    RS_DECODE_ENCODED_DATA_IN_14,
    RS_DECODE_ENCODED_DATA_IN_15,
    RS_DECODE_ENCODED_DATA_IN_16,
    RS_DECODE_ENCODED_DATA_IN_17,
    RS_DECODE_ENCODED_DATA_IN_18,
    RS_DECODE_ENCODED_DATA_IN_19,
    RS_DECODE_ENCODED_DATA_IN_20,
    RS_DECODE_ENCODED_DATA_IN_21,
    RS_DECODE_ENCODED_DATA_IN_22,
    RS_DECODE_ENCODED_DATA_IN_23,
    RS_DECODE_ENCODED_DATA_IN_24,
    RS_DECODE_ENCODED_DATA_IN_25,
    RS_DECODE_ENCODED_DATA_IN_26,
    RS_DECODE_ENCODED_DATA_IN_27,
    RS_DECODE_ENCODED_DATA_IN_28,
    RS_DECODE_ENCODED_DATA_IN_29,
    RS_DECODE_ENCODED_DATA_IN_30,
    RS_DECODE_ENCODED_DATA_IN_31,
    RS_DECODE_ENCODED_DATA_IN_32,
    RS_DECODE_ENCODED_DATA_IN_33,
    RS_DECODE_ENCODED_DATA_IN_34,
    RS_DECODE_ENCODED_DATA_IN_35,
    RS_DECODE_ENCODED_DATA_IN_36,
    RS_DECODE_ENCODED_DATA_IN_37,
    RS_DECODE_ENCODED_DATA_IN_38,
    RS_DECODE_ENCODED_DATA_IN_39,
    RS_DECODE_ENCODED_DATA_IN_40,
    RS_DECODE_ENCODED_DATA_IN_41,
    RS_DECODE_ENCODED_DATA_IN_42,
    RS_DECODE_ENCODED_DATA_IN_43,
    RS_DECODE_ENCODED_DATA_IN_44,
    RS_DECODE_ENCODED_DATA_IN_45,
    RS_DECODE_ENCODED_DATA_IN_46,
    RS_DECODE_ENCODED_DATA_IN_47,
    RS_DECODE_ENCODED_DATA_IN_48,
    RS_DECODE_ENCODED_DATA_IN_49,
    RS_DECODE_ERROR_POS_OUT_0,
    RS_DECODE_ERROR_POS_OUT_1,
    RS_DECODE_ERROR_POS_OUT_2,
    RS_DECODE_ERROR_POS_OUT_3,
    RS_DECODE_ERROR_POS_OUT_4,
    RS_DECODE_ERROR_POS_OUT_5,
    RS_DECODE_ERROR_POS_OUT_6,
    RS_DECODE_ERROR_POS_OUT_7,
    RS_DECODE_ERROR_POS_OUT_8,
    RS_DECODE_ERROR_POS_OUT_9,
    RS_DECODE_ERROR_POS_OUT_10,
    RS_DECODE_ERROR_POS_OUT_11,
    RS_DECODE_ERROR_POS_OUT_12,
    RS_DECODE_ERROR_POS_OUT_13,
    RS_DECODE_ERROR_POS_OUT_14,
    RS_DECODE_ERROR_POS_OUT_15,
    RS_DECODE_ERROR_POS_OUT_16,
    RS_DECODE_ERROR_POS_OUT_17,
    RS_DECODE_ERROR_POS_OUT_18,
    RS_DECODE_ERROR_POS_OUT_19,
    RS_DECODE_ERROR_POS_OUT_20,
    RS_DECODE_ERROR_POS_OUT_21,
    RS_DECODE_ERROR_POS_OUT_22,
    RS_DECODE_ERROR_POS_OUT_23,
    RS_DECODE_ERROR_POS_OUT_24,
    RS_DECODE_ERROR_POS_OUT_25,
    RS_DECODE_ERROR_POS_OUT_26,
    RS_DECODE_ERROR_POS_OUT_27,
    RS_DECODE_ERROR_POS_OUT_28,
    RS_DECODE_ERROR_POS_OUT_29,
    RS_DECODE_ERROR_POS_OUT_30,
    RS_DECODE_ERROR_POS_OUT_31,
    RS_DECODE_ERROR_POS_OUT_32,
    RS_DECODE_ERROR_POS_OUT_33,
    RS_DECODE_ERROR_POS_OUT_34,
    RS_DECODE_ERROR_POS_OUT_35,
    RS_DECODE_ERROR_POS_OUT_36,
    RS_DECODE_ERROR_POS_OUT_37,
    RS_DECODE_ERROR_POS_OUT_38,
    RS_DECODE_ERROR_POS_OUT_39,
    RS_DECODE_ERROR_POS_OUT_40,
    RS_DECODE_ERROR_POS_OUT_41,
    RS_DECODE_ERROR_POS_OUT_42,
    RS_DECODE_ERROR_POS_OUT_43,
    RS_DECODE_ERROR_POS_OUT_44,
    RS_DECODE_ERROR_POS_OUT_45,
    RS_DECODE_ERROR_POS_OUT_46,
    RS_DECODE_ERROR_POS_OUT_47,
    RS_DECODE_ERROR_POS_OUT_48,
    RS_DECODE_ERROR_POS_OUT_49
  } rs_decode_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] RS_DECODE_PERMIT [102] = '{
    4'b 0001, // index[  0] RS_DECODE_CTRL_SIGNALS
    4'b 0001, // index[  1] RS_DECODE_STATE_SIGNALS
    4'b 1111, // index[  2] RS_DECODE_ENCODED_DATA_IN_0
    4'b 1111, // index[  3] RS_DECODE_ENCODED_DATA_IN_1
    4'b 1111, // index[  4] RS_DECODE_ENCODED_DATA_IN_2
    4'b 1111, // index[  5] RS_DECODE_ENCODED_DATA_IN_3
    4'b 1111, // index[  6] RS_DECODE_ENCODED_DATA_IN_4
    4'b 1111, // index[  7] RS_DECODE_ENCODED_DATA_IN_5
    4'b 1111, // index[  8] RS_DECODE_ENCODED_DATA_IN_6
    4'b 1111, // index[  9] RS_DECODE_ENCODED_DATA_IN_7
    4'b 1111, // index[ 10] RS_DECODE_ENCODED_DATA_IN_8
    4'b 1111, // index[ 11] RS_DECODE_ENCODED_DATA_IN_9
    4'b 1111, // index[ 12] RS_DECODE_ENCODED_DATA_IN_10
    4'b 1111, // index[ 13] RS_DECODE_ENCODED_DATA_IN_11
    4'b 1111, // index[ 14] RS_DECODE_ENCODED_DATA_IN_12
    4'b 1111, // index[ 15] RS_DECODE_ENCODED_DATA_IN_13
    4'b 1111, // index[ 16] RS_DECODE_ENCODED_DATA_IN_14
    4'b 1111, // index[ 17] RS_DECODE_ENCODED_DATA_IN_15
    4'b 1111, // index[ 18] RS_DECODE_ENCODED_DATA_IN_16
    4'b 1111, // index[ 19] RS_DECODE_ENCODED_DATA_IN_17
    4'b 1111, // index[ 20] RS_DECODE_ENCODED_DATA_IN_18
    4'b 1111, // index[ 21] RS_DECODE_ENCODED_DATA_IN_19
    4'b 1111, // index[ 22] RS_DECODE_ENCODED_DATA_IN_20
    4'b 1111, // index[ 23] RS_DECODE_ENCODED_DATA_IN_21
    4'b 1111, // index[ 24] RS_DECODE_ENCODED_DATA_IN_22
    4'b 1111, // index[ 25] RS_DECODE_ENCODED_DATA_IN_23
    4'b 1111, // index[ 26] RS_DECODE_ENCODED_DATA_IN_24
    4'b 1111, // index[ 27] RS_DECODE_ENCODED_DATA_IN_25
    4'b 1111, // index[ 28] RS_DECODE_ENCODED_DATA_IN_26
    4'b 1111, // index[ 29] RS_DECODE_ENCODED_DATA_IN_27
    4'b 1111, // index[ 30] RS_DECODE_ENCODED_DATA_IN_28
    4'b 1111, // index[ 31] RS_DECODE_ENCODED_DATA_IN_29
    4'b 1111, // index[ 32] RS_DECODE_ENCODED_DATA_IN_30
    4'b 1111, // index[ 33] RS_DECODE_ENCODED_DATA_IN_31
    4'b 1111, // index[ 34] RS_DECODE_ENCODED_DATA_IN_32
    4'b 1111, // index[ 35] RS_DECODE_ENCODED_DATA_IN_33
    4'b 1111, // index[ 36] RS_DECODE_ENCODED_DATA_IN_34
    4'b 1111, // index[ 37] RS_DECODE_ENCODED_DATA_IN_35
    4'b 1111, // index[ 38] RS_DECODE_ENCODED_DATA_IN_36
    4'b 1111, // index[ 39] RS_DECODE_ENCODED_DATA_IN_37
    4'b 1111, // index[ 40] RS_DECODE_ENCODED_DATA_IN_38
    4'b 1111, // index[ 41] RS_DECODE_ENCODED_DATA_IN_39
    4'b 1111, // index[ 42] RS_DECODE_ENCODED_DATA_IN_40
    4'b 1111, // index[ 43] RS_DECODE_ENCODED_DATA_IN_41
    4'b 1111, // index[ 44] RS_DECODE_ENCODED_DATA_IN_42
    4'b 1111, // index[ 45] RS_DECODE_ENCODED_DATA_IN_43
    4'b 1111, // index[ 46] RS_DECODE_ENCODED_DATA_IN_44
    4'b 1111, // index[ 47] RS_DECODE_ENCODED_DATA_IN_45
    4'b 1111, // index[ 48] RS_DECODE_ENCODED_DATA_IN_46
    4'b 1111, // index[ 49] RS_DECODE_ENCODED_DATA_IN_47
    4'b 1111, // index[ 50] RS_DECODE_ENCODED_DATA_IN_48
    4'b 1111, // index[ 51] RS_DECODE_ENCODED_DATA_IN_49
    4'b 1111, // index[ 52] RS_DECODE_ERROR_POS_OUT_0
    4'b 1111, // index[ 53] RS_DECODE_ERROR_POS_OUT_1
    4'b 1111, // index[ 54] RS_DECODE_ERROR_POS_OUT_2
    4'b 1111, // index[ 55] RS_DECODE_ERROR_POS_OUT_3
    4'b 1111, // index[ 56] RS_DECODE_ERROR_POS_OUT_4
    4'b 1111, // index[ 57] RS_DECODE_ERROR_POS_OUT_5
    4'b 1111, // index[ 58] RS_DECODE_ERROR_POS_OUT_6
    4'b 1111, // index[ 59] RS_DECODE_ERROR_POS_OUT_7
    4'b 1111, // index[ 60] RS_DECODE_ERROR_POS_OUT_8
    4'b 1111, // index[ 61] RS_DECODE_ERROR_POS_OUT_9
    4'b 1111, // index[ 62] RS_DECODE_ERROR_POS_OUT_10
    4'b 1111, // index[ 63] RS_DECODE_ERROR_POS_OUT_11
    4'b 1111, // index[ 64] RS_DECODE_ERROR_POS_OUT_12
    4'b 1111, // index[ 65] RS_DECODE_ERROR_POS_OUT_13
    4'b 1111, // index[ 66] RS_DECODE_ERROR_POS_OUT_14
    4'b 1111, // index[ 67] RS_DECODE_ERROR_POS_OUT_15
    4'b 1111, // index[ 68] RS_DECODE_ERROR_POS_OUT_16
    4'b 1111, // index[ 69] RS_DECODE_ERROR_POS_OUT_17
    4'b 1111, // index[ 70] RS_DECODE_ERROR_POS_OUT_18
    4'b 1111, // index[ 71] RS_DECODE_ERROR_POS_OUT_19
    4'b 1111, // index[ 72] RS_DECODE_ERROR_POS_OUT_20
    4'b 1111, // index[ 73] RS_DECODE_ERROR_POS_OUT_21
    4'b 1111, // index[ 74] RS_DECODE_ERROR_POS_OUT_22
    4'b 1111, // index[ 75] RS_DECODE_ERROR_POS_OUT_23
    4'b 1111, // index[ 76] RS_DECODE_ERROR_POS_OUT_24
    4'b 1111, // index[ 77] RS_DECODE_ERROR_POS_OUT_25
    4'b 1111, // index[ 78] RS_DECODE_ERROR_POS_OUT_26
    4'b 1111, // index[ 79] RS_DECODE_ERROR_POS_OUT_27
    4'b 1111, // index[ 80] RS_DECODE_ERROR_POS_OUT_28
    4'b 1111, // index[ 81] RS_DECODE_ERROR_POS_OUT_29
    4'b 1111, // index[ 82] RS_DECODE_ERROR_POS_OUT_30
    4'b 1111, // index[ 83] RS_DECODE_ERROR_POS_OUT_31
    4'b 1111, // index[ 84] RS_DECODE_ERROR_POS_OUT_32
    4'b 1111, // index[ 85] RS_DECODE_ERROR_POS_OUT_33
    4'b 1111, // index[ 86] RS_DECODE_ERROR_POS_OUT_34
    4'b 1111, // index[ 87] RS_DECODE_ERROR_POS_OUT_35
    4'b 1111, // index[ 88] RS_DECODE_ERROR_POS_OUT_36
    4'b 1111, // index[ 89] RS_DECODE_ERROR_POS_OUT_37
    4'b 1111, // index[ 90] RS_DECODE_ERROR_POS_OUT_38
    4'b 1111, // index[ 91] RS_DECODE_ERROR_POS_OUT_39
    4'b 1111, // index[ 92] RS_DECODE_ERROR_POS_OUT_40
    4'b 1111, // index[ 93] RS_DECODE_ERROR_POS_OUT_41
    4'b 1111, // index[ 94] RS_DECODE_ERROR_POS_OUT_42
    4'b 1111, // index[ 95] RS_DECODE_ERROR_POS_OUT_43
    4'b 1111, // index[ 96] RS_DECODE_ERROR_POS_OUT_44
    4'b 1111, // index[ 97] RS_DECODE_ERROR_POS_OUT_45
    4'b 1111, // index[ 98] RS_DECODE_ERROR_POS_OUT_46
    4'b 1111, // index[ 99] RS_DECODE_ERROR_POS_OUT_47
    4'b 1111, // index[100] RS_DECODE_ERROR_POS_OUT_48
    4'b 1111  // index[101] RS_DECODE_ERROR_POS_OUT_49
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module rs_decode_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output rs_decode_reg_pkg::rs_decode_reg2hw_t reg2hw, // Write
  input  rs_decode_reg_pkg::rs_decode_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import rs_decode_reg_pkg::* ;

  localparam int AW = 9;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [101:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(102)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic ctrl_signals_we;
  logic ctrl_signals_decode_en_qs;
  logic ctrl_signals_decode_en_wd;
  logic ctrl_signals_clrn_qs;
  logic ctrl_signals_clrn_wd;
  logic state_signals_output_valid_bit_qs;
  logic state_signals_ready_bit_qs;
  logic state_signals_with_error_bit_qs;
  logic encoded_data_in_0_we;
  logic [31:0] encoded_data_in_0_qs;
  logic [31:0] encoded_data_in_0_wd;
  logic encoded_data_in_1_we;
  logic [31:0] encoded_data_in_1_qs;
  logic [31:0] encoded_data_in_1_wd;
  logic encoded_data_in_2_we;
  logic [31:0] encoded_data_in_2_qs;
  logic [31:0] encoded_data_in_2_wd;
  logic encoded_data_in_3_we;
  logic [31:0] encoded_data_in_3_qs;
  logic [31:0] encoded_data_in_3_wd;
  logic encoded_data_in_4_we;
  logic [31:0] encoded_data_in_4_qs;
  logic [31:0] encoded_data_in_4_wd;
  logic encoded_data_in_5_we;
  logic [31:0] encoded_data_in_5_qs;
  logic [31:0] encoded_data_in_5_wd;
  logic encoded_data_in_6_we;
  logic [31:0] encoded_data_in_6_qs;
  logic [31:0] encoded_data_in_6_wd;
  logic encoded_data_in_7_we;
  logic [31:0] encoded_data_in_7_qs;
  logic [31:0] encoded_data_in_7_wd;
  logic encoded_data_in_8_we;
  logic [31:0] encoded_data_in_8_qs;
  logic [31:0] encoded_data_in_8_wd;
  logic encoded_data_in_9_we;
  logic [31:0] encoded_data_in_9_qs;
  logic [31:0] encoded_data_in_9_wd;
  logic encoded_data_in_10_we;
  logic [31:0] encoded_data_in_10_qs;
  logic [31:0] encoded_data_in_10_wd;
  logic encoded_data_in_11_we;
  logic [31:0] encoded_data_in_11_qs;
  logic [31:0] encoded_data_in_11_wd;
  logic encoded_data_in_12_we;
  logic [31:0] encoded_data_in_12_qs;
  logic [31:0] encoded_data_in_12_wd;
  logic encoded_data_in_13_we;
  logic [31:0] encoded_data_in_13_qs;
  logic [31:0] encoded_data_in_13_wd;
  logic encoded_data_in_14_we;
  logic [31:0] encoded_data_in_14_qs;
  logic [31:0] encoded_data_in_14_wd;
  logic encoded_data_in_15_we;
  logic [31:0] encoded_data_in_15_qs;
  logic [31:0] encoded_data_in_15_wd;
  logic encoded_data_in_16_we;
  logic [31:0] encoded_data_in_16_qs;
  logic [31:0] encoded_data_in_16_wd;
  logic encoded_data_in_17_we;
  logic [31:0] encoded_data_in_17_qs;
  logic [31:0] encoded_data_in_17_wd;
  logic encoded_data_in_18_we;
  logic [31:0] encoded_data_in_18_qs;
  logic [31:0] encoded_data_in_18_wd;
  logic encoded_data_in_19_we;
  logic [31:0] encoded_data_in_19_qs;
  logic [31:0] encoded_data_in_19_wd;
  logic encoded_data_in_20_we;
  logic [31:0] encoded_data_in_20_qs;
  logic [31:0] encoded_data_in_20_wd;
  logic encoded_data_in_21_we;
  logic [31:0] encoded_data_in_21_qs;
  logic [31:0] encoded_data_in_21_wd;
  logic encoded_data_in_22_we;
  logic [31:0] encoded_data_in_22_qs;
  logic [31:0] encoded_data_in_22_wd;
  logic encoded_data_in_23_we;
  logic [31:0] encoded_data_in_23_qs;
  logic [31:0] encoded_data_in_23_wd;
  logic encoded_data_in_24_we;
  logic [31:0] encoded_data_in_24_qs;
  logic [31:0] encoded_data_in_24_wd;
  logic encoded_data_in_25_we;
  logic [31:0] encoded_data_in_25_qs;
  logic [31:0] encoded_data_in_25_wd;
  logic encoded_data_in_26_we;
  logic [31:0] encoded_data_in_26_qs;
  logic [31:0] encoded_data_in_26_wd;
  logic encoded_data_in_27_we;
  logic [31:0] encoded_data_in_27_qs;
  logic [31:0] encoded_data_in_27_wd;
  logic encoded_data_in_28_we;
  logic [31:0] encoded_data_in_28_qs;
  logic [31:0] encoded_data_in_28_wd;
  logic encoded_data_in_29_we;
  logic [31:0] encoded_data_in_29_qs;
  logic [31:0] encoded_data_in_29_wd;
  logic encoded_data_in_30_we;
  logic [31:0] encoded_data_in_30_qs;
  logic [31:0] encoded_data_in_30_wd;
  logic encoded_data_in_31_we;
  logic [31:0] encoded_data_in_31_qs;
  logic [31:0] encoded_data_in_31_wd;
  logic encoded_data_in_32_we;
  logic [31:0] encoded_data_in_32_qs;
  logic [31:0] encoded_data_in_32_wd;
  logic encoded_data_in_33_we;
  logic [31:0] encoded_data_in_33_qs;
  logic [31:0] encoded_data_in_33_wd;
  logic encoded_data_in_34_we;
  logic [31:0] encoded_data_in_34_qs;
  logic [31:0] encoded_data_in_34_wd;
  logic encoded_data_in_35_we;
  logic [31:0] encoded_data_in_35_qs;
  logic [31:0] encoded_data_in_35_wd;
  logic encoded_data_in_36_we;
  logic [31:0] encoded_data_in_36_qs;
  logic [31:0] encoded_data_in_36_wd;
  logic encoded_data_in_37_we;
  logic [31:0] encoded_data_in_37_qs;
  logic [31:0] encoded_data_in_37_wd;
  logic encoded_data_in_38_we;
  logic [31:0] encoded_data_in_38_qs;
  logic [31:0] encoded_data_in_38_wd;
  logic encoded_data_in_39_we;
  logic [31:0] encoded_data_in_39_qs;
  logic [31:0] encoded_data_in_39_wd;
  logic encoded_data_in_40_we;
  logic [31:0] encoded_data_in_40_qs;
  logic [31:0] encoded_data_in_40_wd;
  logic encoded_data_in_41_we;
  logic [31:0] encoded_data_in_41_qs;
  logic [31:0] encoded_data_in_41_wd;
  logic encoded_data_in_42_we;
  logic [31:0] encoded_data_in_42_qs;
  logic [31:0] encoded_data_in_42_wd;
  logic encoded_data_in_43_we;
  logic [31:0] encoded_data_in_43_qs;
  logic [31:0] encoded_data_in_43_wd;
  logic encoded_data_in_44_we;
  logic [31:0] encoded_data_in_44_qs;
  logic [31:0] encoded_data_in_44_wd;
  logic encoded_data_in_45_we;
  logic [31:0] encoded_data_in_45_qs;
  logic [31:0] encoded_data_in_45_wd;
  logic encoded_data_in_46_we;
  logic [31:0] encoded_data_in_46_qs;
  logic [31:0] encoded_data_in_46_wd;
  logic encoded_data_in_47_we;
  logic [31:0] encoded_data_in_47_qs;
  logic [31:0] encoded_data_in_47_wd;
  logic encoded_data_in_48_we;
  logic [31:0] encoded_data_in_48_qs;
  logic [31:0] encoded_data_in_48_wd;
  logic encoded_data_in_49_we;
  logic [31:0] encoded_data_in_49_qs;
  logic [31:0] encoded_data_in_49_wd;
  logic [31:0] error_pos_out_0_qs;
  logic [31:0] error_pos_out_1_qs;
  logic [31:0] error_pos_out_2_qs;
  logic [31:0] error_pos_out_3_qs;
  logic [31:0] error_pos_out_4_qs;
  logic [31:0] error_pos_out_5_qs;
  logic [31:0] error_pos_out_6_qs;
  logic [31:0] error_pos_out_7_qs;
  logic [31:0] error_pos_out_8_qs;
  logic [31:0] error_pos_out_9_qs;
  logic [31:0] error_pos_out_10_qs;
  logic [31:0] error_pos_out_11_qs;
  logic [31:0] error_pos_out_12_qs;
  logic [31:0] error_pos_out_13_qs;
  logic [31:0] error_pos_out_14_qs;
  logic [31:0] error_pos_out_15_qs;
  logic [31:0] error_pos_out_16_qs;
  logic [31:0] error_pos_out_17_qs;
  logic [31:0] error_pos_out_18_qs;
  logic [31:0] error_pos_out_19_qs;
  logic [31:0] error_pos_out_20_qs;
  logic [31:0] error_pos_out_21_qs;
  logic [31:0] error_pos_out_22_qs;
  logic [31:0] error_pos_out_23_qs;
  logic [31:0] error_pos_out_24_qs;
  logic [31:0] error_pos_out_25_qs;
  logic [31:0] error_pos_out_26_qs;
  logic [31:0] error_pos_out_27_qs;
  logic [31:0] error_pos_out_28_qs;
  logic [31:0] error_pos_out_29_qs;
  logic [31:0] error_pos_out_30_qs;
  logic [31:0] error_pos_out_31_qs;
  logic [31:0] error_pos_out_32_qs;
  logic [31:0] error_pos_out_33_qs;
  logic [31:0] error_pos_out_34_qs;
  logic [31:0] error_pos_out_35_qs;
  logic [31:0] error_pos_out_36_qs;
  logic [31:0] error_pos_out_37_qs;
  logic [31:0] error_pos_out_38_qs;
  logic [31:0] error_pos_out_39_qs;
  logic [31:0] error_pos_out_40_qs;
  logic [31:0] error_pos_out_41_qs;
  logic [31:0] error_pos_out_42_qs;
  logic [31:0] error_pos_out_43_qs;
  logic [31:0] error_pos_out_44_qs;
  logic [31:0] error_pos_out_45_qs;
  logic [31:0] error_pos_out_46_qs;
  logic [31:0] error_pos_out_47_qs;
  logic [31:0] error_pos_out_48_qs;
  logic [31:0] error_pos_out_49_qs;

  // Register instances
  // R[ctrl_signals]: V(False)
  logic ctrl_signals_qe;
  logic [1:0] ctrl_signals_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_ctrl_signals0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&ctrl_signals_flds_we),
    .q_o(ctrl_signals_qe)
  );
  //   F[decode_en]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_decode_en (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_decode_en_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.decode_en.de),
    .d      (hw2reg.ctrl_signals.decode_en.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[0]),
    .q      (reg2hw.ctrl_signals.decode_en.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_decode_en_qs)
  );
  assign reg2hw.ctrl_signals.decode_en.qe = ctrl_signals_qe;

  //   F[clrn]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h1)
  ) u_ctrl_signals_clrn (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_clrn_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.clrn.de),
    .d      (hw2reg.ctrl_signals.clrn.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[1]),
    .q      (reg2hw.ctrl_signals.clrn.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_clrn_qs)
  );
  assign reg2hw.ctrl_signals.clrn.qe = ctrl_signals_qe;


  // R[state_signals]: V(False)
  //   F[output_valid_bit]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_output_valid_bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.output_valid_bit.de),
    .d      (hw2reg.state_signals.output_valid_bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.output_valid_bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_output_valid_bit_qs)
  );

  //   F[ready_bit]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_ready_bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.ready_bit.de),
    .d      (hw2reg.state_signals.ready_bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.ready_bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_ready_bit_qs)
  );

  //   F[with_error_bit]: 2:2
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_with_error_bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.with_error_bit.de),
    .d      (hw2reg.state_signals.with_error_bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.with_error_bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_with_error_bit_qs)
  );


  // Subregister 0 of Multireg encoded_data_in
  // R[encoded_data_in_0]: V(False)
  logic encoded_data_in_0_qe;
  logic [0:0] encoded_data_in_0_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_0_flds_we),
    .q_o(encoded_data_in_0_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_0_we),
    .wd     (encoded_data_in_0_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[0].de),
    .d      (hw2reg.encoded_data_in[0].d),

    // to internal hardware
    .qe     (encoded_data_in_0_flds_we[0]),
    .q      (reg2hw.encoded_data_in[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_0_qs)
  );
  assign reg2hw.encoded_data_in[0].qe = encoded_data_in_0_qe;


  // Subregister 1 of Multireg encoded_data_in
  // R[encoded_data_in_1]: V(False)
  logic encoded_data_in_1_qe;
  logic [0:0] encoded_data_in_1_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in1_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_1_flds_we),
    .q_o(encoded_data_in_1_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_1_we),
    .wd     (encoded_data_in_1_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[1].de),
    .d      (hw2reg.encoded_data_in[1].d),

    // to internal hardware
    .qe     (encoded_data_in_1_flds_we[0]),
    .q      (reg2hw.encoded_data_in[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_1_qs)
  );
  assign reg2hw.encoded_data_in[1].qe = encoded_data_in_1_qe;


  // Subregister 2 of Multireg encoded_data_in
  // R[encoded_data_in_2]: V(False)
  logic encoded_data_in_2_qe;
  logic [0:0] encoded_data_in_2_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in2_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_2_flds_we),
    .q_o(encoded_data_in_2_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_2_we),
    .wd     (encoded_data_in_2_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[2].de),
    .d      (hw2reg.encoded_data_in[2].d),

    // to internal hardware
    .qe     (encoded_data_in_2_flds_we[0]),
    .q      (reg2hw.encoded_data_in[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_2_qs)
  );
  assign reg2hw.encoded_data_in[2].qe = encoded_data_in_2_qe;


  // Subregister 3 of Multireg encoded_data_in
  // R[encoded_data_in_3]: V(False)
  logic encoded_data_in_3_qe;
  logic [0:0] encoded_data_in_3_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in3_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_3_flds_we),
    .q_o(encoded_data_in_3_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_3_we),
    .wd     (encoded_data_in_3_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[3].de),
    .d      (hw2reg.encoded_data_in[3].d),

    // to internal hardware
    .qe     (encoded_data_in_3_flds_we[0]),
    .q      (reg2hw.encoded_data_in[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_3_qs)
  );
  assign reg2hw.encoded_data_in[3].qe = encoded_data_in_3_qe;


  // Subregister 4 of Multireg encoded_data_in
  // R[encoded_data_in_4]: V(False)
  logic encoded_data_in_4_qe;
  logic [0:0] encoded_data_in_4_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in4_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_4_flds_we),
    .q_o(encoded_data_in_4_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_4_we),
    .wd     (encoded_data_in_4_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[4].de),
    .d      (hw2reg.encoded_data_in[4].d),

    // to internal hardware
    .qe     (encoded_data_in_4_flds_we[0]),
    .q      (reg2hw.encoded_data_in[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_4_qs)
  );
  assign reg2hw.encoded_data_in[4].qe = encoded_data_in_4_qe;


  // Subregister 5 of Multireg encoded_data_in
  // R[encoded_data_in_5]: V(False)
  logic encoded_data_in_5_qe;
  logic [0:0] encoded_data_in_5_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in5_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_5_flds_we),
    .q_o(encoded_data_in_5_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_5_we),
    .wd     (encoded_data_in_5_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[5].de),
    .d      (hw2reg.encoded_data_in[5].d),

    // to internal hardware
    .qe     (encoded_data_in_5_flds_we[0]),
    .q      (reg2hw.encoded_data_in[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_5_qs)
  );
  assign reg2hw.encoded_data_in[5].qe = encoded_data_in_5_qe;


  // Subregister 6 of Multireg encoded_data_in
  // R[encoded_data_in_6]: V(False)
  logic encoded_data_in_6_qe;
  logic [0:0] encoded_data_in_6_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in6_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_6_flds_we),
    .q_o(encoded_data_in_6_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_6_we),
    .wd     (encoded_data_in_6_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[6].de),
    .d      (hw2reg.encoded_data_in[6].d),

    // to internal hardware
    .qe     (encoded_data_in_6_flds_we[0]),
    .q      (reg2hw.encoded_data_in[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_6_qs)
  );
  assign reg2hw.encoded_data_in[6].qe = encoded_data_in_6_qe;


  // Subregister 7 of Multireg encoded_data_in
  // R[encoded_data_in_7]: V(False)
  logic encoded_data_in_7_qe;
  logic [0:0] encoded_data_in_7_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in7_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_7_flds_we),
    .q_o(encoded_data_in_7_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_7_we),
    .wd     (encoded_data_in_7_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[7].de),
    .d      (hw2reg.encoded_data_in[7].d),

    // to internal hardware
    .qe     (encoded_data_in_7_flds_we[0]),
    .q      (reg2hw.encoded_data_in[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_7_qs)
  );
  assign reg2hw.encoded_data_in[7].qe = encoded_data_in_7_qe;


  // Subregister 8 of Multireg encoded_data_in
  // R[encoded_data_in_8]: V(False)
  logic encoded_data_in_8_qe;
  logic [0:0] encoded_data_in_8_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in8_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_8_flds_we),
    .q_o(encoded_data_in_8_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_8 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_8_we),
    .wd     (encoded_data_in_8_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[8].de),
    .d      (hw2reg.encoded_data_in[8].d),

    // to internal hardware
    .qe     (encoded_data_in_8_flds_we[0]),
    .q      (reg2hw.encoded_data_in[8].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_8_qs)
  );
  assign reg2hw.encoded_data_in[8].qe = encoded_data_in_8_qe;


  // Subregister 9 of Multireg encoded_data_in
  // R[encoded_data_in_9]: V(False)
  logic encoded_data_in_9_qe;
  logic [0:0] encoded_data_in_9_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in9_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_9_flds_we),
    .q_o(encoded_data_in_9_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_9 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_9_we),
    .wd     (encoded_data_in_9_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[9].de),
    .d      (hw2reg.encoded_data_in[9].d),

    // to internal hardware
    .qe     (encoded_data_in_9_flds_we[0]),
    .q      (reg2hw.encoded_data_in[9].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_9_qs)
  );
  assign reg2hw.encoded_data_in[9].qe = encoded_data_in_9_qe;


  // Subregister 10 of Multireg encoded_data_in
  // R[encoded_data_in_10]: V(False)
  logic encoded_data_in_10_qe;
  logic [0:0] encoded_data_in_10_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in10_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_10_flds_we),
    .q_o(encoded_data_in_10_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_10 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_10_we),
    .wd     (encoded_data_in_10_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[10].de),
    .d      (hw2reg.encoded_data_in[10].d),

    // to internal hardware
    .qe     (encoded_data_in_10_flds_we[0]),
    .q      (reg2hw.encoded_data_in[10].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_10_qs)
  );
  assign reg2hw.encoded_data_in[10].qe = encoded_data_in_10_qe;


  // Subregister 11 of Multireg encoded_data_in
  // R[encoded_data_in_11]: V(False)
  logic encoded_data_in_11_qe;
  logic [0:0] encoded_data_in_11_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in11_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_11_flds_we),
    .q_o(encoded_data_in_11_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_11 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_11_we),
    .wd     (encoded_data_in_11_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[11].de),
    .d      (hw2reg.encoded_data_in[11].d),

    // to internal hardware
    .qe     (encoded_data_in_11_flds_we[0]),
    .q      (reg2hw.encoded_data_in[11].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_11_qs)
  );
  assign reg2hw.encoded_data_in[11].qe = encoded_data_in_11_qe;


  // Subregister 12 of Multireg encoded_data_in
  // R[encoded_data_in_12]: V(False)
  logic encoded_data_in_12_qe;
  logic [0:0] encoded_data_in_12_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in12_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_12_flds_we),
    .q_o(encoded_data_in_12_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_12 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_12_we),
    .wd     (encoded_data_in_12_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[12].de),
    .d      (hw2reg.encoded_data_in[12].d),

    // to internal hardware
    .qe     (encoded_data_in_12_flds_we[0]),
    .q      (reg2hw.encoded_data_in[12].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_12_qs)
  );
  assign reg2hw.encoded_data_in[12].qe = encoded_data_in_12_qe;


  // Subregister 13 of Multireg encoded_data_in
  // R[encoded_data_in_13]: V(False)
  logic encoded_data_in_13_qe;
  logic [0:0] encoded_data_in_13_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in13_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_13_flds_we),
    .q_o(encoded_data_in_13_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_13 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_13_we),
    .wd     (encoded_data_in_13_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[13].de),
    .d      (hw2reg.encoded_data_in[13].d),

    // to internal hardware
    .qe     (encoded_data_in_13_flds_we[0]),
    .q      (reg2hw.encoded_data_in[13].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_13_qs)
  );
  assign reg2hw.encoded_data_in[13].qe = encoded_data_in_13_qe;


  // Subregister 14 of Multireg encoded_data_in
  // R[encoded_data_in_14]: V(False)
  logic encoded_data_in_14_qe;
  logic [0:0] encoded_data_in_14_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in14_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_14_flds_we),
    .q_o(encoded_data_in_14_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_14 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_14_we),
    .wd     (encoded_data_in_14_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[14].de),
    .d      (hw2reg.encoded_data_in[14].d),

    // to internal hardware
    .qe     (encoded_data_in_14_flds_we[0]),
    .q      (reg2hw.encoded_data_in[14].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_14_qs)
  );
  assign reg2hw.encoded_data_in[14].qe = encoded_data_in_14_qe;


  // Subregister 15 of Multireg encoded_data_in
  // R[encoded_data_in_15]: V(False)
  logic encoded_data_in_15_qe;
  logic [0:0] encoded_data_in_15_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in15_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_15_flds_we),
    .q_o(encoded_data_in_15_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_15 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_15_we),
    .wd     (encoded_data_in_15_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[15].de),
    .d      (hw2reg.encoded_data_in[15].d),

    // to internal hardware
    .qe     (encoded_data_in_15_flds_we[0]),
    .q      (reg2hw.encoded_data_in[15].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_15_qs)
  );
  assign reg2hw.encoded_data_in[15].qe = encoded_data_in_15_qe;


  // Subregister 16 of Multireg encoded_data_in
  // R[encoded_data_in_16]: V(False)
  logic encoded_data_in_16_qe;
  logic [0:0] encoded_data_in_16_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in16_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_16_flds_we),
    .q_o(encoded_data_in_16_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_16 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_16_we),
    .wd     (encoded_data_in_16_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[16].de),
    .d      (hw2reg.encoded_data_in[16].d),

    // to internal hardware
    .qe     (encoded_data_in_16_flds_we[0]),
    .q      (reg2hw.encoded_data_in[16].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_16_qs)
  );
  assign reg2hw.encoded_data_in[16].qe = encoded_data_in_16_qe;


  // Subregister 17 of Multireg encoded_data_in
  // R[encoded_data_in_17]: V(False)
  logic encoded_data_in_17_qe;
  logic [0:0] encoded_data_in_17_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in17_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_17_flds_we),
    .q_o(encoded_data_in_17_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_17 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_17_we),
    .wd     (encoded_data_in_17_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[17].de),
    .d      (hw2reg.encoded_data_in[17].d),

    // to internal hardware
    .qe     (encoded_data_in_17_flds_we[0]),
    .q      (reg2hw.encoded_data_in[17].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_17_qs)
  );
  assign reg2hw.encoded_data_in[17].qe = encoded_data_in_17_qe;


  // Subregister 18 of Multireg encoded_data_in
  // R[encoded_data_in_18]: V(False)
  logic encoded_data_in_18_qe;
  logic [0:0] encoded_data_in_18_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in18_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_18_flds_we),
    .q_o(encoded_data_in_18_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_18 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_18_we),
    .wd     (encoded_data_in_18_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[18].de),
    .d      (hw2reg.encoded_data_in[18].d),

    // to internal hardware
    .qe     (encoded_data_in_18_flds_we[0]),
    .q      (reg2hw.encoded_data_in[18].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_18_qs)
  );
  assign reg2hw.encoded_data_in[18].qe = encoded_data_in_18_qe;


  // Subregister 19 of Multireg encoded_data_in
  // R[encoded_data_in_19]: V(False)
  logic encoded_data_in_19_qe;
  logic [0:0] encoded_data_in_19_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in19_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_19_flds_we),
    .q_o(encoded_data_in_19_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_19 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_19_we),
    .wd     (encoded_data_in_19_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[19].de),
    .d      (hw2reg.encoded_data_in[19].d),

    // to internal hardware
    .qe     (encoded_data_in_19_flds_we[0]),
    .q      (reg2hw.encoded_data_in[19].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_19_qs)
  );
  assign reg2hw.encoded_data_in[19].qe = encoded_data_in_19_qe;


  // Subregister 20 of Multireg encoded_data_in
  // R[encoded_data_in_20]: V(False)
  logic encoded_data_in_20_qe;
  logic [0:0] encoded_data_in_20_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in20_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_20_flds_we),
    .q_o(encoded_data_in_20_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_20 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_20_we),
    .wd     (encoded_data_in_20_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[20].de),
    .d      (hw2reg.encoded_data_in[20].d),

    // to internal hardware
    .qe     (encoded_data_in_20_flds_we[0]),
    .q      (reg2hw.encoded_data_in[20].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_20_qs)
  );
  assign reg2hw.encoded_data_in[20].qe = encoded_data_in_20_qe;


  // Subregister 21 of Multireg encoded_data_in
  // R[encoded_data_in_21]: V(False)
  logic encoded_data_in_21_qe;
  logic [0:0] encoded_data_in_21_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in21_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_21_flds_we),
    .q_o(encoded_data_in_21_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_21 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_21_we),
    .wd     (encoded_data_in_21_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[21].de),
    .d      (hw2reg.encoded_data_in[21].d),

    // to internal hardware
    .qe     (encoded_data_in_21_flds_we[0]),
    .q      (reg2hw.encoded_data_in[21].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_21_qs)
  );
  assign reg2hw.encoded_data_in[21].qe = encoded_data_in_21_qe;


  // Subregister 22 of Multireg encoded_data_in
  // R[encoded_data_in_22]: V(False)
  logic encoded_data_in_22_qe;
  logic [0:0] encoded_data_in_22_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in22_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_22_flds_we),
    .q_o(encoded_data_in_22_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_22 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_22_we),
    .wd     (encoded_data_in_22_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[22].de),
    .d      (hw2reg.encoded_data_in[22].d),

    // to internal hardware
    .qe     (encoded_data_in_22_flds_we[0]),
    .q      (reg2hw.encoded_data_in[22].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_22_qs)
  );
  assign reg2hw.encoded_data_in[22].qe = encoded_data_in_22_qe;


  // Subregister 23 of Multireg encoded_data_in
  // R[encoded_data_in_23]: V(False)
  logic encoded_data_in_23_qe;
  logic [0:0] encoded_data_in_23_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in23_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_23_flds_we),
    .q_o(encoded_data_in_23_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_23 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_23_we),
    .wd     (encoded_data_in_23_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[23].de),
    .d      (hw2reg.encoded_data_in[23].d),

    // to internal hardware
    .qe     (encoded_data_in_23_flds_we[0]),
    .q      (reg2hw.encoded_data_in[23].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_23_qs)
  );
  assign reg2hw.encoded_data_in[23].qe = encoded_data_in_23_qe;


  // Subregister 24 of Multireg encoded_data_in
  // R[encoded_data_in_24]: V(False)
  logic encoded_data_in_24_qe;
  logic [0:0] encoded_data_in_24_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in24_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_24_flds_we),
    .q_o(encoded_data_in_24_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_24 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_24_we),
    .wd     (encoded_data_in_24_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[24].de),
    .d      (hw2reg.encoded_data_in[24].d),

    // to internal hardware
    .qe     (encoded_data_in_24_flds_we[0]),
    .q      (reg2hw.encoded_data_in[24].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_24_qs)
  );
  assign reg2hw.encoded_data_in[24].qe = encoded_data_in_24_qe;


  // Subregister 25 of Multireg encoded_data_in
  // R[encoded_data_in_25]: V(False)
  logic encoded_data_in_25_qe;
  logic [0:0] encoded_data_in_25_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in25_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_25_flds_we),
    .q_o(encoded_data_in_25_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_25 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_25_we),
    .wd     (encoded_data_in_25_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[25].de),
    .d      (hw2reg.encoded_data_in[25].d),

    // to internal hardware
    .qe     (encoded_data_in_25_flds_we[0]),
    .q      (reg2hw.encoded_data_in[25].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_25_qs)
  );
  assign reg2hw.encoded_data_in[25].qe = encoded_data_in_25_qe;


  // Subregister 26 of Multireg encoded_data_in
  // R[encoded_data_in_26]: V(False)
  logic encoded_data_in_26_qe;
  logic [0:0] encoded_data_in_26_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in26_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_26_flds_we),
    .q_o(encoded_data_in_26_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_26 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_26_we),
    .wd     (encoded_data_in_26_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[26].de),
    .d      (hw2reg.encoded_data_in[26].d),

    // to internal hardware
    .qe     (encoded_data_in_26_flds_we[0]),
    .q      (reg2hw.encoded_data_in[26].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_26_qs)
  );
  assign reg2hw.encoded_data_in[26].qe = encoded_data_in_26_qe;


  // Subregister 27 of Multireg encoded_data_in
  // R[encoded_data_in_27]: V(False)
  logic encoded_data_in_27_qe;
  logic [0:0] encoded_data_in_27_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in27_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_27_flds_we),
    .q_o(encoded_data_in_27_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_27 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_27_we),
    .wd     (encoded_data_in_27_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[27].de),
    .d      (hw2reg.encoded_data_in[27].d),

    // to internal hardware
    .qe     (encoded_data_in_27_flds_we[0]),
    .q      (reg2hw.encoded_data_in[27].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_27_qs)
  );
  assign reg2hw.encoded_data_in[27].qe = encoded_data_in_27_qe;


  // Subregister 28 of Multireg encoded_data_in
  // R[encoded_data_in_28]: V(False)
  logic encoded_data_in_28_qe;
  logic [0:0] encoded_data_in_28_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in28_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_28_flds_we),
    .q_o(encoded_data_in_28_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_28 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_28_we),
    .wd     (encoded_data_in_28_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[28].de),
    .d      (hw2reg.encoded_data_in[28].d),

    // to internal hardware
    .qe     (encoded_data_in_28_flds_we[0]),
    .q      (reg2hw.encoded_data_in[28].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_28_qs)
  );
  assign reg2hw.encoded_data_in[28].qe = encoded_data_in_28_qe;


  // Subregister 29 of Multireg encoded_data_in
  // R[encoded_data_in_29]: V(False)
  logic encoded_data_in_29_qe;
  logic [0:0] encoded_data_in_29_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in29_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_29_flds_we),
    .q_o(encoded_data_in_29_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_29 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_29_we),
    .wd     (encoded_data_in_29_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[29].de),
    .d      (hw2reg.encoded_data_in[29].d),

    // to internal hardware
    .qe     (encoded_data_in_29_flds_we[0]),
    .q      (reg2hw.encoded_data_in[29].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_29_qs)
  );
  assign reg2hw.encoded_data_in[29].qe = encoded_data_in_29_qe;


  // Subregister 30 of Multireg encoded_data_in
  // R[encoded_data_in_30]: V(False)
  logic encoded_data_in_30_qe;
  logic [0:0] encoded_data_in_30_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in30_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_30_flds_we),
    .q_o(encoded_data_in_30_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_30 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_30_we),
    .wd     (encoded_data_in_30_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[30].de),
    .d      (hw2reg.encoded_data_in[30].d),

    // to internal hardware
    .qe     (encoded_data_in_30_flds_we[0]),
    .q      (reg2hw.encoded_data_in[30].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_30_qs)
  );
  assign reg2hw.encoded_data_in[30].qe = encoded_data_in_30_qe;


  // Subregister 31 of Multireg encoded_data_in
  // R[encoded_data_in_31]: V(False)
  logic encoded_data_in_31_qe;
  logic [0:0] encoded_data_in_31_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in31_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_31_flds_we),
    .q_o(encoded_data_in_31_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_31 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_31_we),
    .wd     (encoded_data_in_31_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[31].de),
    .d      (hw2reg.encoded_data_in[31].d),

    // to internal hardware
    .qe     (encoded_data_in_31_flds_we[0]),
    .q      (reg2hw.encoded_data_in[31].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_31_qs)
  );
  assign reg2hw.encoded_data_in[31].qe = encoded_data_in_31_qe;


  // Subregister 32 of Multireg encoded_data_in
  // R[encoded_data_in_32]: V(False)
  logic encoded_data_in_32_qe;
  logic [0:0] encoded_data_in_32_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in32_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_32_flds_we),
    .q_o(encoded_data_in_32_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_32 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_32_we),
    .wd     (encoded_data_in_32_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[32].de),
    .d      (hw2reg.encoded_data_in[32].d),

    // to internal hardware
    .qe     (encoded_data_in_32_flds_we[0]),
    .q      (reg2hw.encoded_data_in[32].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_32_qs)
  );
  assign reg2hw.encoded_data_in[32].qe = encoded_data_in_32_qe;


  // Subregister 33 of Multireg encoded_data_in
  // R[encoded_data_in_33]: V(False)
  logic encoded_data_in_33_qe;
  logic [0:0] encoded_data_in_33_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in33_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_33_flds_we),
    .q_o(encoded_data_in_33_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_33 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_33_we),
    .wd     (encoded_data_in_33_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[33].de),
    .d      (hw2reg.encoded_data_in[33].d),

    // to internal hardware
    .qe     (encoded_data_in_33_flds_we[0]),
    .q      (reg2hw.encoded_data_in[33].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_33_qs)
  );
  assign reg2hw.encoded_data_in[33].qe = encoded_data_in_33_qe;


  // Subregister 34 of Multireg encoded_data_in
  // R[encoded_data_in_34]: V(False)
  logic encoded_data_in_34_qe;
  logic [0:0] encoded_data_in_34_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in34_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_34_flds_we),
    .q_o(encoded_data_in_34_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_34 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_34_we),
    .wd     (encoded_data_in_34_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[34].de),
    .d      (hw2reg.encoded_data_in[34].d),

    // to internal hardware
    .qe     (encoded_data_in_34_flds_we[0]),
    .q      (reg2hw.encoded_data_in[34].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_34_qs)
  );
  assign reg2hw.encoded_data_in[34].qe = encoded_data_in_34_qe;


  // Subregister 35 of Multireg encoded_data_in
  // R[encoded_data_in_35]: V(False)
  logic encoded_data_in_35_qe;
  logic [0:0] encoded_data_in_35_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in35_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_35_flds_we),
    .q_o(encoded_data_in_35_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_35 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_35_we),
    .wd     (encoded_data_in_35_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[35].de),
    .d      (hw2reg.encoded_data_in[35].d),

    // to internal hardware
    .qe     (encoded_data_in_35_flds_we[0]),
    .q      (reg2hw.encoded_data_in[35].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_35_qs)
  );
  assign reg2hw.encoded_data_in[35].qe = encoded_data_in_35_qe;


  // Subregister 36 of Multireg encoded_data_in
  // R[encoded_data_in_36]: V(False)
  logic encoded_data_in_36_qe;
  logic [0:0] encoded_data_in_36_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in36_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_36_flds_we),
    .q_o(encoded_data_in_36_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_36 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_36_we),
    .wd     (encoded_data_in_36_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[36].de),
    .d      (hw2reg.encoded_data_in[36].d),

    // to internal hardware
    .qe     (encoded_data_in_36_flds_we[0]),
    .q      (reg2hw.encoded_data_in[36].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_36_qs)
  );
  assign reg2hw.encoded_data_in[36].qe = encoded_data_in_36_qe;


  // Subregister 37 of Multireg encoded_data_in
  // R[encoded_data_in_37]: V(False)
  logic encoded_data_in_37_qe;
  logic [0:0] encoded_data_in_37_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in37_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_37_flds_we),
    .q_o(encoded_data_in_37_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_37 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_37_we),
    .wd     (encoded_data_in_37_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[37].de),
    .d      (hw2reg.encoded_data_in[37].d),

    // to internal hardware
    .qe     (encoded_data_in_37_flds_we[0]),
    .q      (reg2hw.encoded_data_in[37].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_37_qs)
  );
  assign reg2hw.encoded_data_in[37].qe = encoded_data_in_37_qe;


  // Subregister 38 of Multireg encoded_data_in
  // R[encoded_data_in_38]: V(False)
  logic encoded_data_in_38_qe;
  logic [0:0] encoded_data_in_38_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in38_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_38_flds_we),
    .q_o(encoded_data_in_38_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_38 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_38_we),
    .wd     (encoded_data_in_38_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[38].de),
    .d      (hw2reg.encoded_data_in[38].d),

    // to internal hardware
    .qe     (encoded_data_in_38_flds_we[0]),
    .q      (reg2hw.encoded_data_in[38].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_38_qs)
  );
  assign reg2hw.encoded_data_in[38].qe = encoded_data_in_38_qe;


  // Subregister 39 of Multireg encoded_data_in
  // R[encoded_data_in_39]: V(False)
  logic encoded_data_in_39_qe;
  logic [0:0] encoded_data_in_39_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in39_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_39_flds_we),
    .q_o(encoded_data_in_39_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_39 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_39_we),
    .wd     (encoded_data_in_39_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[39].de),
    .d      (hw2reg.encoded_data_in[39].d),

    // to internal hardware
    .qe     (encoded_data_in_39_flds_we[0]),
    .q      (reg2hw.encoded_data_in[39].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_39_qs)
  );
  assign reg2hw.encoded_data_in[39].qe = encoded_data_in_39_qe;


  // Subregister 40 of Multireg encoded_data_in
  // R[encoded_data_in_40]: V(False)
  logic encoded_data_in_40_qe;
  logic [0:0] encoded_data_in_40_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in40_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_40_flds_we),
    .q_o(encoded_data_in_40_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_40 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_40_we),
    .wd     (encoded_data_in_40_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[40].de),
    .d      (hw2reg.encoded_data_in[40].d),

    // to internal hardware
    .qe     (encoded_data_in_40_flds_we[0]),
    .q      (reg2hw.encoded_data_in[40].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_40_qs)
  );
  assign reg2hw.encoded_data_in[40].qe = encoded_data_in_40_qe;


  // Subregister 41 of Multireg encoded_data_in
  // R[encoded_data_in_41]: V(False)
  logic encoded_data_in_41_qe;
  logic [0:0] encoded_data_in_41_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in41_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_41_flds_we),
    .q_o(encoded_data_in_41_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_41 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_41_we),
    .wd     (encoded_data_in_41_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[41].de),
    .d      (hw2reg.encoded_data_in[41].d),

    // to internal hardware
    .qe     (encoded_data_in_41_flds_we[0]),
    .q      (reg2hw.encoded_data_in[41].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_41_qs)
  );
  assign reg2hw.encoded_data_in[41].qe = encoded_data_in_41_qe;


  // Subregister 42 of Multireg encoded_data_in
  // R[encoded_data_in_42]: V(False)
  logic encoded_data_in_42_qe;
  logic [0:0] encoded_data_in_42_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in42_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_42_flds_we),
    .q_o(encoded_data_in_42_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_42 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_42_we),
    .wd     (encoded_data_in_42_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[42].de),
    .d      (hw2reg.encoded_data_in[42].d),

    // to internal hardware
    .qe     (encoded_data_in_42_flds_we[0]),
    .q      (reg2hw.encoded_data_in[42].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_42_qs)
  );
  assign reg2hw.encoded_data_in[42].qe = encoded_data_in_42_qe;


  // Subregister 43 of Multireg encoded_data_in
  // R[encoded_data_in_43]: V(False)
  logic encoded_data_in_43_qe;
  logic [0:0] encoded_data_in_43_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in43_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_43_flds_we),
    .q_o(encoded_data_in_43_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_43 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_43_we),
    .wd     (encoded_data_in_43_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[43].de),
    .d      (hw2reg.encoded_data_in[43].d),

    // to internal hardware
    .qe     (encoded_data_in_43_flds_we[0]),
    .q      (reg2hw.encoded_data_in[43].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_43_qs)
  );
  assign reg2hw.encoded_data_in[43].qe = encoded_data_in_43_qe;


  // Subregister 44 of Multireg encoded_data_in
  // R[encoded_data_in_44]: V(False)
  logic encoded_data_in_44_qe;
  logic [0:0] encoded_data_in_44_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in44_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_44_flds_we),
    .q_o(encoded_data_in_44_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_44 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_44_we),
    .wd     (encoded_data_in_44_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[44].de),
    .d      (hw2reg.encoded_data_in[44].d),

    // to internal hardware
    .qe     (encoded_data_in_44_flds_we[0]),
    .q      (reg2hw.encoded_data_in[44].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_44_qs)
  );
  assign reg2hw.encoded_data_in[44].qe = encoded_data_in_44_qe;


  // Subregister 45 of Multireg encoded_data_in
  // R[encoded_data_in_45]: V(False)
  logic encoded_data_in_45_qe;
  logic [0:0] encoded_data_in_45_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in45_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_45_flds_we),
    .q_o(encoded_data_in_45_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_45 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_45_we),
    .wd     (encoded_data_in_45_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[45].de),
    .d      (hw2reg.encoded_data_in[45].d),

    // to internal hardware
    .qe     (encoded_data_in_45_flds_we[0]),
    .q      (reg2hw.encoded_data_in[45].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_45_qs)
  );
  assign reg2hw.encoded_data_in[45].qe = encoded_data_in_45_qe;


  // Subregister 46 of Multireg encoded_data_in
  // R[encoded_data_in_46]: V(False)
  logic encoded_data_in_46_qe;
  logic [0:0] encoded_data_in_46_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in46_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_46_flds_we),
    .q_o(encoded_data_in_46_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_46 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_46_we),
    .wd     (encoded_data_in_46_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[46].de),
    .d      (hw2reg.encoded_data_in[46].d),

    // to internal hardware
    .qe     (encoded_data_in_46_flds_we[0]),
    .q      (reg2hw.encoded_data_in[46].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_46_qs)
  );
  assign reg2hw.encoded_data_in[46].qe = encoded_data_in_46_qe;


  // Subregister 47 of Multireg encoded_data_in
  // R[encoded_data_in_47]: V(False)
  logic encoded_data_in_47_qe;
  logic [0:0] encoded_data_in_47_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in47_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_47_flds_we),
    .q_o(encoded_data_in_47_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_47 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_47_we),
    .wd     (encoded_data_in_47_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[47].de),
    .d      (hw2reg.encoded_data_in[47].d),

    // to internal hardware
    .qe     (encoded_data_in_47_flds_we[0]),
    .q      (reg2hw.encoded_data_in[47].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_47_qs)
  );
  assign reg2hw.encoded_data_in[47].qe = encoded_data_in_47_qe;


  // Subregister 48 of Multireg encoded_data_in
  // R[encoded_data_in_48]: V(False)
  logic encoded_data_in_48_qe;
  logic [0:0] encoded_data_in_48_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in48_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_48_flds_we),
    .q_o(encoded_data_in_48_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_48 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_48_we),
    .wd     (encoded_data_in_48_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[48].de),
    .d      (hw2reg.encoded_data_in[48].d),

    // to internal hardware
    .qe     (encoded_data_in_48_flds_we[0]),
    .q      (reg2hw.encoded_data_in[48].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_48_qs)
  );
  assign reg2hw.encoded_data_in[48].qe = encoded_data_in_48_qe;


  // Subregister 49 of Multireg encoded_data_in
  // R[encoded_data_in_49]: V(False)
  logic encoded_data_in_49_qe;
  logic [0:0] encoded_data_in_49_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_encoded_data_in49_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&encoded_data_in_49_flds_we),
    .q_o(encoded_data_in_49_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_encoded_data_in_49 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (encoded_data_in_49_we),
    .wd     (encoded_data_in_49_wd),

    // from internal hardware
    .de     (hw2reg.encoded_data_in[49].de),
    .d      (hw2reg.encoded_data_in[49].d),

    // to internal hardware
    .qe     (encoded_data_in_49_flds_we[0]),
    .q      (reg2hw.encoded_data_in[49].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_in_49_qs)
  );
  assign reg2hw.encoded_data_in[49].qe = encoded_data_in_49_qe;


  // Subregister 0 of Multireg error_pos_out
  // R[error_pos_out_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[0].de),
    .d      (hw2reg.error_pos_out[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_0_qs)
  );


  // Subregister 1 of Multireg error_pos_out
  // R[error_pos_out_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[1].de),
    .d      (hw2reg.error_pos_out[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_1_qs)
  );


  // Subregister 2 of Multireg error_pos_out
  // R[error_pos_out_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[2].de),
    .d      (hw2reg.error_pos_out[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_2_qs)
  );


  // Subregister 3 of Multireg error_pos_out
  // R[error_pos_out_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[3].de),
    .d      (hw2reg.error_pos_out[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_3_qs)
  );


  // Subregister 4 of Multireg error_pos_out
  // R[error_pos_out_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[4].de),
    .d      (hw2reg.error_pos_out[4].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_4_qs)
  );


  // Subregister 5 of Multireg error_pos_out
  // R[error_pos_out_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[5].de),
    .d      (hw2reg.error_pos_out[5].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_5_qs)
  );


  // Subregister 6 of Multireg error_pos_out
  // R[error_pos_out_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[6].de),
    .d      (hw2reg.error_pos_out[6].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_6_qs)
  );


  // Subregister 7 of Multireg error_pos_out
  // R[error_pos_out_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[7].de),
    .d      (hw2reg.error_pos_out[7].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_7_qs)
  );


  // Subregister 8 of Multireg error_pos_out
  // R[error_pos_out_8]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_8 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[8].de),
    .d      (hw2reg.error_pos_out[8].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[8].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_8_qs)
  );


  // Subregister 9 of Multireg error_pos_out
  // R[error_pos_out_9]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_9 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[9].de),
    .d      (hw2reg.error_pos_out[9].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[9].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_9_qs)
  );


  // Subregister 10 of Multireg error_pos_out
  // R[error_pos_out_10]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_10 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[10].de),
    .d      (hw2reg.error_pos_out[10].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[10].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_10_qs)
  );


  // Subregister 11 of Multireg error_pos_out
  // R[error_pos_out_11]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_11 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[11].de),
    .d      (hw2reg.error_pos_out[11].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[11].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_11_qs)
  );


  // Subregister 12 of Multireg error_pos_out
  // R[error_pos_out_12]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_12 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[12].de),
    .d      (hw2reg.error_pos_out[12].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[12].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_12_qs)
  );


  // Subregister 13 of Multireg error_pos_out
  // R[error_pos_out_13]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_13 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[13].de),
    .d      (hw2reg.error_pos_out[13].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[13].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_13_qs)
  );


  // Subregister 14 of Multireg error_pos_out
  // R[error_pos_out_14]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_14 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[14].de),
    .d      (hw2reg.error_pos_out[14].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[14].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_14_qs)
  );


  // Subregister 15 of Multireg error_pos_out
  // R[error_pos_out_15]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_15 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[15].de),
    .d      (hw2reg.error_pos_out[15].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[15].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_15_qs)
  );


  // Subregister 16 of Multireg error_pos_out
  // R[error_pos_out_16]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_16 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[16].de),
    .d      (hw2reg.error_pos_out[16].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[16].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_16_qs)
  );


  // Subregister 17 of Multireg error_pos_out
  // R[error_pos_out_17]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_17 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[17].de),
    .d      (hw2reg.error_pos_out[17].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[17].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_17_qs)
  );


  // Subregister 18 of Multireg error_pos_out
  // R[error_pos_out_18]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_18 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[18].de),
    .d      (hw2reg.error_pos_out[18].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[18].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_18_qs)
  );


  // Subregister 19 of Multireg error_pos_out
  // R[error_pos_out_19]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_19 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[19].de),
    .d      (hw2reg.error_pos_out[19].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[19].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_19_qs)
  );


  // Subregister 20 of Multireg error_pos_out
  // R[error_pos_out_20]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_20 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[20].de),
    .d      (hw2reg.error_pos_out[20].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[20].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_20_qs)
  );


  // Subregister 21 of Multireg error_pos_out
  // R[error_pos_out_21]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_21 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[21].de),
    .d      (hw2reg.error_pos_out[21].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[21].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_21_qs)
  );


  // Subregister 22 of Multireg error_pos_out
  // R[error_pos_out_22]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_22 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[22].de),
    .d      (hw2reg.error_pos_out[22].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[22].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_22_qs)
  );


  // Subregister 23 of Multireg error_pos_out
  // R[error_pos_out_23]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_23 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[23].de),
    .d      (hw2reg.error_pos_out[23].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[23].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_23_qs)
  );


  // Subregister 24 of Multireg error_pos_out
  // R[error_pos_out_24]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_24 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[24].de),
    .d      (hw2reg.error_pos_out[24].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[24].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_24_qs)
  );


  // Subregister 25 of Multireg error_pos_out
  // R[error_pos_out_25]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_25 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[25].de),
    .d      (hw2reg.error_pos_out[25].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[25].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_25_qs)
  );


  // Subregister 26 of Multireg error_pos_out
  // R[error_pos_out_26]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_26 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[26].de),
    .d      (hw2reg.error_pos_out[26].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[26].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_26_qs)
  );


  // Subregister 27 of Multireg error_pos_out
  // R[error_pos_out_27]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_27 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[27].de),
    .d      (hw2reg.error_pos_out[27].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[27].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_27_qs)
  );


  // Subregister 28 of Multireg error_pos_out
  // R[error_pos_out_28]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_28 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[28].de),
    .d      (hw2reg.error_pos_out[28].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[28].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_28_qs)
  );


  // Subregister 29 of Multireg error_pos_out
  // R[error_pos_out_29]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_29 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[29].de),
    .d      (hw2reg.error_pos_out[29].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[29].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_29_qs)
  );


  // Subregister 30 of Multireg error_pos_out
  // R[error_pos_out_30]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_30 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[30].de),
    .d      (hw2reg.error_pos_out[30].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[30].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_30_qs)
  );


  // Subregister 31 of Multireg error_pos_out
  // R[error_pos_out_31]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_31 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[31].de),
    .d      (hw2reg.error_pos_out[31].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[31].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_31_qs)
  );


  // Subregister 32 of Multireg error_pos_out
  // R[error_pos_out_32]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_32 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[32].de),
    .d      (hw2reg.error_pos_out[32].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[32].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_32_qs)
  );


  // Subregister 33 of Multireg error_pos_out
  // R[error_pos_out_33]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_33 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[33].de),
    .d      (hw2reg.error_pos_out[33].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[33].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_33_qs)
  );


  // Subregister 34 of Multireg error_pos_out
  // R[error_pos_out_34]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_34 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[34].de),
    .d      (hw2reg.error_pos_out[34].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[34].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_34_qs)
  );


  // Subregister 35 of Multireg error_pos_out
  // R[error_pos_out_35]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_35 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[35].de),
    .d      (hw2reg.error_pos_out[35].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[35].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_35_qs)
  );


  // Subregister 36 of Multireg error_pos_out
  // R[error_pos_out_36]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_36 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[36].de),
    .d      (hw2reg.error_pos_out[36].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[36].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_36_qs)
  );


  // Subregister 37 of Multireg error_pos_out
  // R[error_pos_out_37]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_37 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[37].de),
    .d      (hw2reg.error_pos_out[37].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[37].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_37_qs)
  );


  // Subregister 38 of Multireg error_pos_out
  // R[error_pos_out_38]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_38 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[38].de),
    .d      (hw2reg.error_pos_out[38].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[38].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_38_qs)
  );


  // Subregister 39 of Multireg error_pos_out
  // R[error_pos_out_39]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_39 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[39].de),
    .d      (hw2reg.error_pos_out[39].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[39].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_39_qs)
  );


  // Subregister 40 of Multireg error_pos_out
  // R[error_pos_out_40]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_40 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[40].de),
    .d      (hw2reg.error_pos_out[40].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[40].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_40_qs)
  );


  // Subregister 41 of Multireg error_pos_out
  // R[error_pos_out_41]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_41 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[41].de),
    .d      (hw2reg.error_pos_out[41].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[41].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_41_qs)
  );


  // Subregister 42 of Multireg error_pos_out
  // R[error_pos_out_42]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_42 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[42].de),
    .d      (hw2reg.error_pos_out[42].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[42].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_42_qs)
  );


  // Subregister 43 of Multireg error_pos_out
  // R[error_pos_out_43]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_43 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[43].de),
    .d      (hw2reg.error_pos_out[43].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[43].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_43_qs)
  );


  // Subregister 44 of Multireg error_pos_out
  // R[error_pos_out_44]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_44 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[44].de),
    .d      (hw2reg.error_pos_out[44].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[44].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_44_qs)
  );


  // Subregister 45 of Multireg error_pos_out
  // R[error_pos_out_45]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_45 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[45].de),
    .d      (hw2reg.error_pos_out[45].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[45].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_45_qs)
  );


  // Subregister 46 of Multireg error_pos_out
  // R[error_pos_out_46]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_46 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[46].de),
    .d      (hw2reg.error_pos_out[46].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[46].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_46_qs)
  );


  // Subregister 47 of Multireg error_pos_out
  // R[error_pos_out_47]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_47 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[47].de),
    .d      (hw2reg.error_pos_out[47].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[47].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_47_qs)
  );


  // Subregister 48 of Multireg error_pos_out
  // R[error_pos_out_48]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_48 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[48].de),
    .d      (hw2reg.error_pos_out[48].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[48].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_48_qs)
  );


  // Subregister 49 of Multireg error_pos_out
  // R[error_pos_out_49]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_error_pos_out_49 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.error_pos_out[49].de),
    .d      (hw2reg.error_pos_out[49].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.error_pos_out[49].q),
    .ds     (),

    // to register interface (read)
    .qs     (error_pos_out_49_qs)
  );



  logic [101:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[  0] = (reg_addr == RS_DECODE_CTRL_SIGNALS_OFFSET);
    addr_hit[  1] = (reg_addr == RS_DECODE_STATE_SIGNALS_OFFSET);
    addr_hit[  2] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_0_OFFSET);
    addr_hit[  3] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_1_OFFSET);
    addr_hit[  4] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_2_OFFSET);
    addr_hit[  5] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_3_OFFSET);
    addr_hit[  6] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_4_OFFSET);
    addr_hit[  7] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_5_OFFSET);
    addr_hit[  8] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_6_OFFSET);
    addr_hit[  9] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_7_OFFSET);
    addr_hit[ 10] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_8_OFFSET);
    addr_hit[ 11] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_9_OFFSET);
    addr_hit[ 12] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_10_OFFSET);
    addr_hit[ 13] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_11_OFFSET);
    addr_hit[ 14] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_12_OFFSET);
    addr_hit[ 15] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_13_OFFSET);
    addr_hit[ 16] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_14_OFFSET);
    addr_hit[ 17] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_15_OFFSET);
    addr_hit[ 18] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_16_OFFSET);
    addr_hit[ 19] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_17_OFFSET);
    addr_hit[ 20] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_18_OFFSET);
    addr_hit[ 21] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_19_OFFSET);
    addr_hit[ 22] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_20_OFFSET);
    addr_hit[ 23] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_21_OFFSET);
    addr_hit[ 24] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_22_OFFSET);
    addr_hit[ 25] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_23_OFFSET);
    addr_hit[ 26] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_24_OFFSET);
    addr_hit[ 27] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_25_OFFSET);
    addr_hit[ 28] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_26_OFFSET);
    addr_hit[ 29] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_27_OFFSET);
    addr_hit[ 30] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_28_OFFSET);
    addr_hit[ 31] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_29_OFFSET);
    addr_hit[ 32] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_30_OFFSET);
    addr_hit[ 33] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_31_OFFSET);
    addr_hit[ 34] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_32_OFFSET);
    addr_hit[ 35] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_33_OFFSET);
    addr_hit[ 36] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_34_OFFSET);
    addr_hit[ 37] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_35_OFFSET);
    addr_hit[ 38] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_36_OFFSET);
    addr_hit[ 39] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_37_OFFSET);
    addr_hit[ 40] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_38_OFFSET);
    addr_hit[ 41] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_39_OFFSET);
    addr_hit[ 42] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_40_OFFSET);
    addr_hit[ 43] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_41_OFFSET);
    addr_hit[ 44] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_42_OFFSET);
    addr_hit[ 45] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_43_OFFSET);
    addr_hit[ 46] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_44_OFFSET);
    addr_hit[ 47] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_45_OFFSET);
    addr_hit[ 48] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_46_OFFSET);
    addr_hit[ 49] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_47_OFFSET);
    addr_hit[ 50] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_48_OFFSET);
    addr_hit[ 51] = (reg_addr == RS_DECODE_ENCODED_DATA_IN_49_OFFSET);
    addr_hit[ 52] = (reg_addr == RS_DECODE_ERROR_POS_OUT_0_OFFSET);
    addr_hit[ 53] = (reg_addr == RS_DECODE_ERROR_POS_OUT_1_OFFSET);
    addr_hit[ 54] = (reg_addr == RS_DECODE_ERROR_POS_OUT_2_OFFSET);
    addr_hit[ 55] = (reg_addr == RS_DECODE_ERROR_POS_OUT_3_OFFSET);
    addr_hit[ 56] = (reg_addr == RS_DECODE_ERROR_POS_OUT_4_OFFSET);
    addr_hit[ 57] = (reg_addr == RS_DECODE_ERROR_POS_OUT_5_OFFSET);
    addr_hit[ 58] = (reg_addr == RS_DECODE_ERROR_POS_OUT_6_OFFSET);
    addr_hit[ 59] = (reg_addr == RS_DECODE_ERROR_POS_OUT_7_OFFSET);
    addr_hit[ 60] = (reg_addr == RS_DECODE_ERROR_POS_OUT_8_OFFSET);
    addr_hit[ 61] = (reg_addr == RS_DECODE_ERROR_POS_OUT_9_OFFSET);
    addr_hit[ 62] = (reg_addr == RS_DECODE_ERROR_POS_OUT_10_OFFSET);
    addr_hit[ 63] = (reg_addr == RS_DECODE_ERROR_POS_OUT_11_OFFSET);
    addr_hit[ 64] = (reg_addr == RS_DECODE_ERROR_POS_OUT_12_OFFSET);
    addr_hit[ 65] = (reg_addr == RS_DECODE_ERROR_POS_OUT_13_OFFSET);
    addr_hit[ 66] = (reg_addr == RS_DECODE_ERROR_POS_OUT_14_OFFSET);
    addr_hit[ 67] = (reg_addr == RS_DECODE_ERROR_POS_OUT_15_OFFSET);
    addr_hit[ 68] = (reg_addr == RS_DECODE_ERROR_POS_OUT_16_OFFSET);
    addr_hit[ 69] = (reg_addr == RS_DECODE_ERROR_POS_OUT_17_OFFSET);
    addr_hit[ 70] = (reg_addr == RS_DECODE_ERROR_POS_OUT_18_OFFSET);
    addr_hit[ 71] = (reg_addr == RS_DECODE_ERROR_POS_OUT_19_OFFSET);
    addr_hit[ 72] = (reg_addr == RS_DECODE_ERROR_POS_OUT_20_OFFSET);
    addr_hit[ 73] = (reg_addr == RS_DECODE_ERROR_POS_OUT_21_OFFSET);
    addr_hit[ 74] = (reg_addr == RS_DECODE_ERROR_POS_OUT_22_OFFSET);
    addr_hit[ 75] = (reg_addr == RS_DECODE_ERROR_POS_OUT_23_OFFSET);
    addr_hit[ 76] = (reg_addr == RS_DECODE_ERROR_POS_OUT_24_OFFSET);
    addr_hit[ 77] = (reg_addr == RS_DECODE_ERROR_POS_OUT_25_OFFSET);
    addr_hit[ 78] = (reg_addr == RS_DECODE_ERROR_POS_OUT_26_OFFSET);
    addr_hit[ 79] = (reg_addr == RS_DECODE_ERROR_POS_OUT_27_OFFSET);
    addr_hit[ 80] = (reg_addr == RS_DECODE_ERROR_POS_OUT_28_OFFSET);
    addr_hit[ 81] = (reg_addr == RS_DECODE_ERROR_POS_OUT_29_OFFSET);
    addr_hit[ 82] = (reg_addr == RS_DECODE_ERROR_POS_OUT_30_OFFSET);
    addr_hit[ 83] = (reg_addr == RS_DECODE_ERROR_POS_OUT_31_OFFSET);
    addr_hit[ 84] = (reg_addr == RS_DECODE_ERROR_POS_OUT_32_OFFSET);
    addr_hit[ 85] = (reg_addr == RS_DECODE_ERROR_POS_OUT_33_OFFSET);
    addr_hit[ 86] = (reg_addr == RS_DECODE_ERROR_POS_OUT_34_OFFSET);
    addr_hit[ 87] = (reg_addr == RS_DECODE_ERROR_POS_OUT_35_OFFSET);
    addr_hit[ 88] = (reg_addr == RS_DECODE_ERROR_POS_OUT_36_OFFSET);
    addr_hit[ 89] = (reg_addr == RS_DECODE_ERROR_POS_OUT_37_OFFSET);
    addr_hit[ 90] = (reg_addr == RS_DECODE_ERROR_POS_OUT_38_OFFSET);
    addr_hit[ 91] = (reg_addr == RS_DECODE_ERROR_POS_OUT_39_OFFSET);
    addr_hit[ 92] = (reg_addr == RS_DECODE_ERROR_POS_OUT_40_OFFSET);
    addr_hit[ 93] = (reg_addr == RS_DECODE_ERROR_POS_OUT_41_OFFSET);
    addr_hit[ 94] = (reg_addr == RS_DECODE_ERROR_POS_OUT_42_OFFSET);
    addr_hit[ 95] = (reg_addr == RS_DECODE_ERROR_POS_OUT_43_OFFSET);
    addr_hit[ 96] = (reg_addr == RS_DECODE_ERROR_POS_OUT_44_OFFSET);
    addr_hit[ 97] = (reg_addr == RS_DECODE_ERROR_POS_OUT_45_OFFSET);
    addr_hit[ 98] = (reg_addr == RS_DECODE_ERROR_POS_OUT_46_OFFSET);
    addr_hit[ 99] = (reg_addr == RS_DECODE_ERROR_POS_OUT_47_OFFSET);
    addr_hit[100] = (reg_addr == RS_DECODE_ERROR_POS_OUT_48_OFFSET);
    addr_hit[101] = (reg_addr == RS_DECODE_ERROR_POS_OUT_49_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[  0] & (|(RS_DECODE_PERMIT[  0] & ~reg_be))) |
               (addr_hit[  1] & (|(RS_DECODE_PERMIT[  1] & ~reg_be))) |
               (addr_hit[  2] & (|(RS_DECODE_PERMIT[  2] & ~reg_be))) |
               (addr_hit[  3] & (|(RS_DECODE_PERMIT[  3] & ~reg_be))) |
               (addr_hit[  4] & (|(RS_DECODE_PERMIT[  4] & ~reg_be))) |
               (addr_hit[  5] & (|(RS_DECODE_PERMIT[  5] & ~reg_be))) |
               (addr_hit[  6] & (|(RS_DECODE_PERMIT[  6] & ~reg_be))) |
               (addr_hit[  7] & (|(RS_DECODE_PERMIT[  7] & ~reg_be))) |
               (addr_hit[  8] & (|(RS_DECODE_PERMIT[  8] & ~reg_be))) |
               (addr_hit[  9] & (|(RS_DECODE_PERMIT[  9] & ~reg_be))) |
               (addr_hit[ 10] & (|(RS_DECODE_PERMIT[ 10] & ~reg_be))) |
               (addr_hit[ 11] & (|(RS_DECODE_PERMIT[ 11] & ~reg_be))) |
               (addr_hit[ 12] & (|(RS_DECODE_PERMIT[ 12] & ~reg_be))) |
               (addr_hit[ 13] & (|(RS_DECODE_PERMIT[ 13] & ~reg_be))) |
               (addr_hit[ 14] & (|(RS_DECODE_PERMIT[ 14] & ~reg_be))) |
               (addr_hit[ 15] & (|(RS_DECODE_PERMIT[ 15] & ~reg_be))) |
               (addr_hit[ 16] & (|(RS_DECODE_PERMIT[ 16] & ~reg_be))) |
               (addr_hit[ 17] & (|(RS_DECODE_PERMIT[ 17] & ~reg_be))) |
               (addr_hit[ 18] & (|(RS_DECODE_PERMIT[ 18] & ~reg_be))) |
               (addr_hit[ 19] & (|(RS_DECODE_PERMIT[ 19] & ~reg_be))) |
               (addr_hit[ 20] & (|(RS_DECODE_PERMIT[ 20] & ~reg_be))) |
               (addr_hit[ 21] & (|(RS_DECODE_PERMIT[ 21] & ~reg_be))) |
               (addr_hit[ 22] & (|(RS_DECODE_PERMIT[ 22] & ~reg_be))) |
               (addr_hit[ 23] & (|(RS_DECODE_PERMIT[ 23] & ~reg_be))) |
               (addr_hit[ 24] & (|(RS_DECODE_PERMIT[ 24] & ~reg_be))) |
               (addr_hit[ 25] & (|(RS_DECODE_PERMIT[ 25] & ~reg_be))) |
               (addr_hit[ 26] & (|(RS_DECODE_PERMIT[ 26] & ~reg_be))) |
               (addr_hit[ 27] & (|(RS_DECODE_PERMIT[ 27] & ~reg_be))) |
               (addr_hit[ 28] & (|(RS_DECODE_PERMIT[ 28] & ~reg_be))) |
               (addr_hit[ 29] & (|(RS_DECODE_PERMIT[ 29] & ~reg_be))) |
               (addr_hit[ 30] & (|(RS_DECODE_PERMIT[ 30] & ~reg_be))) |
               (addr_hit[ 31] & (|(RS_DECODE_PERMIT[ 31] & ~reg_be))) |
               (addr_hit[ 32] & (|(RS_DECODE_PERMIT[ 32] & ~reg_be))) |
               (addr_hit[ 33] & (|(RS_DECODE_PERMIT[ 33] & ~reg_be))) |
               (addr_hit[ 34] & (|(RS_DECODE_PERMIT[ 34] & ~reg_be))) |
               (addr_hit[ 35] & (|(RS_DECODE_PERMIT[ 35] & ~reg_be))) |
               (addr_hit[ 36] & (|(RS_DECODE_PERMIT[ 36] & ~reg_be))) |
               (addr_hit[ 37] & (|(RS_DECODE_PERMIT[ 37] & ~reg_be))) |
               (addr_hit[ 38] & (|(RS_DECODE_PERMIT[ 38] & ~reg_be))) |
               (addr_hit[ 39] & (|(RS_DECODE_PERMIT[ 39] & ~reg_be))) |
               (addr_hit[ 40] & (|(RS_DECODE_PERMIT[ 40] & ~reg_be))) |
               (addr_hit[ 41] & (|(RS_DECODE_PERMIT[ 41] & ~reg_be))) |
               (addr_hit[ 42] & (|(RS_DECODE_PERMIT[ 42] & ~reg_be))) |
               (addr_hit[ 43] & (|(RS_DECODE_PERMIT[ 43] & ~reg_be))) |
               (addr_hit[ 44] & (|(RS_DECODE_PERMIT[ 44] & ~reg_be))) |
               (addr_hit[ 45] & (|(RS_DECODE_PERMIT[ 45] & ~reg_be))) |
               (addr_hit[ 46] & (|(RS_DECODE_PERMIT[ 46] & ~reg_be))) |
               (addr_hit[ 47] & (|(RS_DECODE_PERMIT[ 47] & ~reg_be))) |
               (addr_hit[ 48] & (|(RS_DECODE_PERMIT[ 48] & ~reg_be))) |
               (addr_hit[ 49] & (|(RS_DECODE_PERMIT[ 49] & ~reg_be))) |
               (addr_hit[ 50] & (|(RS_DECODE_PERMIT[ 50] & ~reg_be))) |
               (addr_hit[ 51] & (|(RS_DECODE_PERMIT[ 51] & ~reg_be))) |
               (addr_hit[ 52] & (|(RS_DECODE_PERMIT[ 52] & ~reg_be))) |
               (addr_hit[ 53] & (|(RS_DECODE_PERMIT[ 53] & ~reg_be))) |
               (addr_hit[ 54] & (|(RS_DECODE_PERMIT[ 54] & ~reg_be))) |
               (addr_hit[ 55] & (|(RS_DECODE_PERMIT[ 55] & ~reg_be))) |
               (addr_hit[ 56] & (|(RS_DECODE_PERMIT[ 56] & ~reg_be))) |
               (addr_hit[ 57] & (|(RS_DECODE_PERMIT[ 57] & ~reg_be))) |
               (addr_hit[ 58] & (|(RS_DECODE_PERMIT[ 58] & ~reg_be))) |
               (addr_hit[ 59] & (|(RS_DECODE_PERMIT[ 59] & ~reg_be))) |
               (addr_hit[ 60] & (|(RS_DECODE_PERMIT[ 60] & ~reg_be))) |
               (addr_hit[ 61] & (|(RS_DECODE_PERMIT[ 61] & ~reg_be))) |
               (addr_hit[ 62] & (|(RS_DECODE_PERMIT[ 62] & ~reg_be))) |
               (addr_hit[ 63] & (|(RS_DECODE_PERMIT[ 63] & ~reg_be))) |
               (addr_hit[ 64] & (|(RS_DECODE_PERMIT[ 64] & ~reg_be))) |
               (addr_hit[ 65] & (|(RS_DECODE_PERMIT[ 65] & ~reg_be))) |
               (addr_hit[ 66] & (|(RS_DECODE_PERMIT[ 66] & ~reg_be))) |
               (addr_hit[ 67] & (|(RS_DECODE_PERMIT[ 67] & ~reg_be))) |
               (addr_hit[ 68] & (|(RS_DECODE_PERMIT[ 68] & ~reg_be))) |
               (addr_hit[ 69] & (|(RS_DECODE_PERMIT[ 69] & ~reg_be))) |
               (addr_hit[ 70] & (|(RS_DECODE_PERMIT[ 70] & ~reg_be))) |
               (addr_hit[ 71] & (|(RS_DECODE_PERMIT[ 71] & ~reg_be))) |
               (addr_hit[ 72] & (|(RS_DECODE_PERMIT[ 72] & ~reg_be))) |
               (addr_hit[ 73] & (|(RS_DECODE_PERMIT[ 73] & ~reg_be))) |
               (addr_hit[ 74] & (|(RS_DECODE_PERMIT[ 74] & ~reg_be))) |
               (addr_hit[ 75] & (|(RS_DECODE_PERMIT[ 75] & ~reg_be))) |
               (addr_hit[ 76] & (|(RS_DECODE_PERMIT[ 76] & ~reg_be))) |
               (addr_hit[ 77] & (|(RS_DECODE_PERMIT[ 77] & ~reg_be))) |
               (addr_hit[ 78] & (|(RS_DECODE_PERMIT[ 78] & ~reg_be))) |
               (addr_hit[ 79] & (|(RS_DECODE_PERMIT[ 79] & ~reg_be))) |
               (addr_hit[ 80] & (|(RS_DECODE_PERMIT[ 80] & ~reg_be))) |
               (addr_hit[ 81] & (|(RS_DECODE_PERMIT[ 81] & ~reg_be))) |
               (addr_hit[ 82] & (|(RS_DECODE_PERMIT[ 82] & ~reg_be))) |
               (addr_hit[ 83] & (|(RS_DECODE_PERMIT[ 83] & ~reg_be))) |
               (addr_hit[ 84] & (|(RS_DECODE_PERMIT[ 84] & ~reg_be))) |
               (addr_hit[ 85] & (|(RS_DECODE_PERMIT[ 85] & ~reg_be))) |
               (addr_hit[ 86] & (|(RS_DECODE_PERMIT[ 86] & ~reg_be))) |
               (addr_hit[ 87] & (|(RS_DECODE_PERMIT[ 87] & ~reg_be))) |
               (addr_hit[ 88] & (|(RS_DECODE_PERMIT[ 88] & ~reg_be))) |
               (addr_hit[ 89] & (|(RS_DECODE_PERMIT[ 89] & ~reg_be))) |
               (addr_hit[ 90] & (|(RS_DECODE_PERMIT[ 90] & ~reg_be))) |
               (addr_hit[ 91] & (|(RS_DECODE_PERMIT[ 91] & ~reg_be))) |
               (addr_hit[ 92] & (|(RS_DECODE_PERMIT[ 92] & ~reg_be))) |
               (addr_hit[ 93] & (|(RS_DECODE_PERMIT[ 93] & ~reg_be))) |
               (addr_hit[ 94] & (|(RS_DECODE_PERMIT[ 94] & ~reg_be))) |
               (addr_hit[ 95] & (|(RS_DECODE_PERMIT[ 95] & ~reg_be))) |
               (addr_hit[ 96] & (|(RS_DECODE_PERMIT[ 96] & ~reg_be))) |
               (addr_hit[ 97] & (|(RS_DECODE_PERMIT[ 97] & ~reg_be))) |
               (addr_hit[ 98] & (|(RS_DECODE_PERMIT[ 98] & ~reg_be))) |
               (addr_hit[ 99] & (|(RS_DECODE_PERMIT[ 99] & ~reg_be))) |
               (addr_hit[100] & (|(RS_DECODE_PERMIT[100] & ~reg_be))) |
               (addr_hit[101] & (|(RS_DECODE_PERMIT[101] & ~reg_be)))));
  end

  // Generate write-enables
  assign ctrl_signals_we = addr_hit[0] & reg_we & !reg_error;

  assign ctrl_signals_decode_en_wd = reg_wdata[0];

  assign ctrl_signals_clrn_wd = reg_wdata[1];
  assign encoded_data_in_0_we = addr_hit[2] & reg_we & !reg_error;

  assign encoded_data_in_0_wd = reg_wdata[31:0];
  assign encoded_data_in_1_we = addr_hit[3] & reg_we & !reg_error;

  assign encoded_data_in_1_wd = reg_wdata[31:0];
  assign encoded_data_in_2_we = addr_hit[4] & reg_we & !reg_error;

  assign encoded_data_in_2_wd = reg_wdata[31:0];
  assign encoded_data_in_3_we = addr_hit[5] & reg_we & !reg_error;

  assign encoded_data_in_3_wd = reg_wdata[31:0];
  assign encoded_data_in_4_we = addr_hit[6] & reg_we & !reg_error;

  assign encoded_data_in_4_wd = reg_wdata[31:0];
  assign encoded_data_in_5_we = addr_hit[7] & reg_we & !reg_error;

  assign encoded_data_in_5_wd = reg_wdata[31:0];
  assign encoded_data_in_6_we = addr_hit[8] & reg_we & !reg_error;

  assign encoded_data_in_6_wd = reg_wdata[31:0];
  assign encoded_data_in_7_we = addr_hit[9] & reg_we & !reg_error;

  assign encoded_data_in_7_wd = reg_wdata[31:0];
  assign encoded_data_in_8_we = addr_hit[10] & reg_we & !reg_error;

  assign encoded_data_in_8_wd = reg_wdata[31:0];
  assign encoded_data_in_9_we = addr_hit[11] & reg_we & !reg_error;

  assign encoded_data_in_9_wd = reg_wdata[31:0];
  assign encoded_data_in_10_we = addr_hit[12] & reg_we & !reg_error;

  assign encoded_data_in_10_wd = reg_wdata[31:0];
  assign encoded_data_in_11_we = addr_hit[13] & reg_we & !reg_error;

  assign encoded_data_in_11_wd = reg_wdata[31:0];
  assign encoded_data_in_12_we = addr_hit[14] & reg_we & !reg_error;

  assign encoded_data_in_12_wd = reg_wdata[31:0];
  assign encoded_data_in_13_we = addr_hit[15] & reg_we & !reg_error;

  assign encoded_data_in_13_wd = reg_wdata[31:0];
  assign encoded_data_in_14_we = addr_hit[16] & reg_we & !reg_error;

  assign encoded_data_in_14_wd = reg_wdata[31:0];
  assign encoded_data_in_15_we = addr_hit[17] & reg_we & !reg_error;

  assign encoded_data_in_15_wd = reg_wdata[31:0];
  assign encoded_data_in_16_we = addr_hit[18] & reg_we & !reg_error;

  assign encoded_data_in_16_wd = reg_wdata[31:0];
  assign encoded_data_in_17_we = addr_hit[19] & reg_we & !reg_error;

  assign encoded_data_in_17_wd = reg_wdata[31:0];
  assign encoded_data_in_18_we = addr_hit[20] & reg_we & !reg_error;

  assign encoded_data_in_18_wd = reg_wdata[31:0];
  assign encoded_data_in_19_we = addr_hit[21] & reg_we & !reg_error;

  assign encoded_data_in_19_wd = reg_wdata[31:0];
  assign encoded_data_in_20_we = addr_hit[22] & reg_we & !reg_error;

  assign encoded_data_in_20_wd = reg_wdata[31:0];
  assign encoded_data_in_21_we = addr_hit[23] & reg_we & !reg_error;

  assign encoded_data_in_21_wd = reg_wdata[31:0];
  assign encoded_data_in_22_we = addr_hit[24] & reg_we & !reg_error;

  assign encoded_data_in_22_wd = reg_wdata[31:0];
  assign encoded_data_in_23_we = addr_hit[25] & reg_we & !reg_error;

  assign encoded_data_in_23_wd = reg_wdata[31:0];
  assign encoded_data_in_24_we = addr_hit[26] & reg_we & !reg_error;

  assign encoded_data_in_24_wd = reg_wdata[31:0];
  assign encoded_data_in_25_we = addr_hit[27] & reg_we & !reg_error;

  assign encoded_data_in_25_wd = reg_wdata[31:0];
  assign encoded_data_in_26_we = addr_hit[28] & reg_we & !reg_error;

  assign encoded_data_in_26_wd = reg_wdata[31:0];
  assign encoded_data_in_27_we = addr_hit[29] & reg_we & !reg_error;

  assign encoded_data_in_27_wd = reg_wdata[31:0];
  assign encoded_data_in_28_we = addr_hit[30] & reg_we & !reg_error;

  assign encoded_data_in_28_wd = reg_wdata[31:0];
  assign encoded_data_in_29_we = addr_hit[31] & reg_we & !reg_error;

  assign encoded_data_in_29_wd = reg_wdata[31:0];
  assign encoded_data_in_30_we = addr_hit[32] & reg_we & !reg_error;

  assign encoded_data_in_30_wd = reg_wdata[31:0];
  assign encoded_data_in_31_we = addr_hit[33] & reg_we & !reg_error;

  assign encoded_data_in_31_wd = reg_wdata[31:0];
  assign encoded_data_in_32_we = addr_hit[34] & reg_we & !reg_error;

  assign encoded_data_in_32_wd = reg_wdata[31:0];
  assign encoded_data_in_33_we = addr_hit[35] & reg_we & !reg_error;

  assign encoded_data_in_33_wd = reg_wdata[31:0];
  assign encoded_data_in_34_we = addr_hit[36] & reg_we & !reg_error;

  assign encoded_data_in_34_wd = reg_wdata[31:0];
  assign encoded_data_in_35_we = addr_hit[37] & reg_we & !reg_error;

  assign encoded_data_in_35_wd = reg_wdata[31:0];
  assign encoded_data_in_36_we = addr_hit[38] & reg_we & !reg_error;

  assign encoded_data_in_36_wd = reg_wdata[31:0];
  assign encoded_data_in_37_we = addr_hit[39] & reg_we & !reg_error;

  assign encoded_data_in_37_wd = reg_wdata[31:0];
  assign encoded_data_in_38_we = addr_hit[40] & reg_we & !reg_error;

  assign encoded_data_in_38_wd = reg_wdata[31:0];
  assign encoded_data_in_39_we = addr_hit[41] & reg_we & !reg_error;

  assign encoded_data_in_39_wd = reg_wdata[31:0];
  assign encoded_data_in_40_we = addr_hit[42] & reg_we & !reg_error;

  assign encoded_data_in_40_wd = reg_wdata[31:0];
  assign encoded_data_in_41_we = addr_hit[43] & reg_we & !reg_error;

  assign encoded_data_in_41_wd = reg_wdata[31:0];
  assign encoded_data_in_42_we = addr_hit[44] & reg_we & !reg_error;

  assign encoded_data_in_42_wd = reg_wdata[31:0];
  assign encoded_data_in_43_we = addr_hit[45] & reg_we & !reg_error;

  assign encoded_data_in_43_wd = reg_wdata[31:0];
  assign encoded_data_in_44_we = addr_hit[46] & reg_we & !reg_error;

  assign encoded_data_in_44_wd = reg_wdata[31:0];
  assign encoded_data_in_45_we = addr_hit[47] & reg_we & !reg_error;

  assign encoded_data_in_45_wd = reg_wdata[31:0];
  assign encoded_data_in_46_we = addr_hit[48] & reg_we & !reg_error;

  assign encoded_data_in_46_wd = reg_wdata[31:0];
  assign encoded_data_in_47_we = addr_hit[49] & reg_we & !reg_error;

  assign encoded_data_in_47_wd = reg_wdata[31:0];
  assign encoded_data_in_48_we = addr_hit[50] & reg_we & !reg_error;

  assign encoded_data_in_48_wd = reg_wdata[31:0];
  assign encoded_data_in_49_we = addr_hit[51] & reg_we & !reg_error;

  assign encoded_data_in_49_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = ctrl_signals_we;
    reg_we_check[1] = 1'b0;
    reg_we_check[2] = encoded_data_in_0_we;
    reg_we_check[3] = encoded_data_in_1_we;
    reg_we_check[4] = encoded_data_in_2_we;
    reg_we_check[5] = encoded_data_in_3_we;
    reg_we_check[6] = encoded_data_in_4_we;
    reg_we_check[7] = encoded_data_in_5_we;
    reg_we_check[8] = encoded_data_in_6_we;
    reg_we_check[9] = encoded_data_in_7_we;
    reg_we_check[10] = encoded_data_in_8_we;
    reg_we_check[11] = encoded_data_in_9_we;
    reg_we_check[12] = encoded_data_in_10_we;
    reg_we_check[13] = encoded_data_in_11_we;
    reg_we_check[14] = encoded_data_in_12_we;
    reg_we_check[15] = encoded_data_in_13_we;
    reg_we_check[16] = encoded_data_in_14_we;
    reg_we_check[17] = encoded_data_in_15_we;
    reg_we_check[18] = encoded_data_in_16_we;
    reg_we_check[19] = encoded_data_in_17_we;
    reg_we_check[20] = encoded_data_in_18_we;
    reg_we_check[21] = encoded_data_in_19_we;
    reg_we_check[22] = encoded_data_in_20_we;
    reg_we_check[23] = encoded_data_in_21_we;
    reg_we_check[24] = encoded_data_in_22_we;
    reg_we_check[25] = encoded_data_in_23_we;
    reg_we_check[26] = encoded_data_in_24_we;
    reg_we_check[27] = encoded_data_in_25_we;
    reg_we_check[28] = encoded_data_in_26_we;
    reg_we_check[29] = encoded_data_in_27_we;
    reg_we_check[30] = encoded_data_in_28_we;
    reg_we_check[31] = encoded_data_in_29_we;
    reg_we_check[32] = encoded_data_in_30_we;
    reg_we_check[33] = encoded_data_in_31_we;
    reg_we_check[34] = encoded_data_in_32_we;
    reg_we_check[35] = encoded_data_in_33_we;
    reg_we_check[36] = encoded_data_in_34_we;
    reg_we_check[37] = encoded_data_in_35_we;
    reg_we_check[38] = encoded_data_in_36_we;
    reg_we_check[39] = encoded_data_in_37_we;
    reg_we_check[40] = encoded_data_in_38_we;
    reg_we_check[41] = encoded_data_in_39_we;
    reg_we_check[42] = encoded_data_in_40_we;
    reg_we_check[43] = encoded_data_in_41_we;
    reg_we_check[44] = encoded_data_in_42_we;
    reg_we_check[45] = encoded_data_in_43_we;
    reg_we_check[46] = encoded_data_in_44_we;
    reg_we_check[47] = encoded_data_in_45_we;
    reg_we_check[48] = encoded_data_in_46_we;
    reg_we_check[49] = encoded_data_in_47_we;
    reg_we_check[50] = encoded_data_in_48_we;
    reg_we_check[51] = encoded_data_in_49_we;
    reg_we_check[52] = 1'b0;
    reg_we_check[53] = 1'b0;
    reg_we_check[54] = 1'b0;
    reg_we_check[55] = 1'b0;
    reg_we_check[56] = 1'b0;
    reg_we_check[57] = 1'b0;
    reg_we_check[58] = 1'b0;
    reg_we_check[59] = 1'b0;
    reg_we_check[60] = 1'b0;
    reg_we_check[61] = 1'b0;
    reg_we_check[62] = 1'b0;
    reg_we_check[63] = 1'b0;
    reg_we_check[64] = 1'b0;
    reg_we_check[65] = 1'b0;
    reg_we_check[66] = 1'b0;
    reg_we_check[67] = 1'b0;
    reg_we_check[68] = 1'b0;
    reg_we_check[69] = 1'b0;
    reg_we_check[70] = 1'b0;
    reg_we_check[71] = 1'b0;
    reg_we_check[72] = 1'b0;
    reg_we_check[73] = 1'b0;
    reg_we_check[74] = 1'b0;
    reg_we_check[75] = 1'b0;
    reg_we_check[76] = 1'b0;
    reg_we_check[77] = 1'b0;
    reg_we_check[78] = 1'b0;
    reg_we_check[79] = 1'b0;
    reg_we_check[80] = 1'b0;
    reg_we_check[81] = 1'b0;
    reg_we_check[82] = 1'b0;
    reg_we_check[83] = 1'b0;
    reg_we_check[84] = 1'b0;
    reg_we_check[85] = 1'b0;
    reg_we_check[86] = 1'b0;
    reg_we_check[87] = 1'b0;
    reg_we_check[88] = 1'b0;
    reg_we_check[89] = 1'b0;
    reg_we_check[90] = 1'b0;
    reg_we_check[91] = 1'b0;
    reg_we_check[92] = 1'b0;
    reg_we_check[93] = 1'b0;
    reg_we_check[94] = 1'b0;
    reg_we_check[95] = 1'b0;
    reg_we_check[96] = 1'b0;
    reg_we_check[97] = 1'b0;
    reg_we_check[98] = 1'b0;
    reg_we_check[99] = 1'b0;
    reg_we_check[100] = 1'b0;
    reg_we_check[101] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = ctrl_signals_decode_en_qs;
        reg_rdata_next[1] = ctrl_signals_clrn_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = state_signals_output_valid_bit_qs;
        reg_rdata_next[1] = state_signals_ready_bit_qs;
        reg_rdata_next[2] = state_signals_with_error_bit_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = encoded_data_in_0_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = encoded_data_in_1_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = encoded_data_in_2_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = encoded_data_in_3_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = encoded_data_in_4_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = encoded_data_in_5_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = encoded_data_in_6_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = encoded_data_in_7_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = encoded_data_in_8_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = encoded_data_in_9_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = encoded_data_in_10_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = encoded_data_in_11_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = encoded_data_in_12_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = encoded_data_in_13_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = encoded_data_in_14_qs;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = encoded_data_in_15_qs;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = encoded_data_in_16_qs;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = encoded_data_in_17_qs;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = encoded_data_in_18_qs;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = encoded_data_in_19_qs;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = encoded_data_in_20_qs;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = encoded_data_in_21_qs;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = encoded_data_in_22_qs;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = encoded_data_in_23_qs;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = encoded_data_in_24_qs;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = encoded_data_in_25_qs;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = encoded_data_in_26_qs;
      end

      addr_hit[29]: begin
        reg_rdata_next[31:0] = encoded_data_in_27_qs;
      end

      addr_hit[30]: begin
        reg_rdata_next[31:0] = encoded_data_in_28_qs;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = encoded_data_in_29_qs;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = encoded_data_in_30_qs;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = encoded_data_in_31_qs;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = encoded_data_in_32_qs;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = encoded_data_in_33_qs;
      end

      addr_hit[36]: begin
        reg_rdata_next[31:0] = encoded_data_in_34_qs;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = encoded_data_in_35_qs;
      end

      addr_hit[38]: begin
        reg_rdata_next[31:0] = encoded_data_in_36_qs;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = encoded_data_in_37_qs;
      end

      addr_hit[40]: begin
        reg_rdata_next[31:0] = encoded_data_in_38_qs;
      end

      addr_hit[41]: begin
        reg_rdata_next[31:0] = encoded_data_in_39_qs;
      end

      addr_hit[42]: begin
        reg_rdata_next[31:0] = encoded_data_in_40_qs;
      end

      addr_hit[43]: begin
        reg_rdata_next[31:0] = encoded_data_in_41_qs;
      end

      addr_hit[44]: begin
        reg_rdata_next[31:0] = encoded_data_in_42_qs;
      end

      addr_hit[45]: begin
        reg_rdata_next[31:0] = encoded_data_in_43_qs;
      end

      addr_hit[46]: begin
        reg_rdata_next[31:0] = encoded_data_in_44_qs;
      end

      addr_hit[47]: begin
        reg_rdata_next[31:0] = encoded_data_in_45_qs;
      end

      addr_hit[48]: begin
        reg_rdata_next[31:0] = encoded_data_in_46_qs;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = encoded_data_in_47_qs;
      end

      addr_hit[50]: begin
        reg_rdata_next[31:0] = encoded_data_in_48_qs;
      end

      addr_hit[51]: begin
        reg_rdata_next[31:0] = encoded_data_in_49_qs;
      end

      addr_hit[52]: begin
        reg_rdata_next[31:0] = error_pos_out_0_qs;
      end

      addr_hit[53]: begin
        reg_rdata_next[31:0] = error_pos_out_1_qs;
      end

      addr_hit[54]: begin
        reg_rdata_next[31:0] = error_pos_out_2_qs;
      end

      addr_hit[55]: begin
        reg_rdata_next[31:0] = error_pos_out_3_qs;
      end

      addr_hit[56]: begin
        reg_rdata_next[31:0] = error_pos_out_4_qs;
      end

      addr_hit[57]: begin
        reg_rdata_next[31:0] = error_pos_out_5_qs;
      end

      addr_hit[58]: begin
        reg_rdata_next[31:0] = error_pos_out_6_qs;
      end

      addr_hit[59]: begin
        reg_rdata_next[31:0] = error_pos_out_7_qs;
      end

      addr_hit[60]: begin
        reg_rdata_next[31:0] = error_pos_out_8_qs;
      end

      addr_hit[61]: begin
        reg_rdata_next[31:0] = error_pos_out_9_qs;
      end

      addr_hit[62]: begin
        reg_rdata_next[31:0] = error_pos_out_10_qs;
      end

      addr_hit[63]: begin
        reg_rdata_next[31:0] = error_pos_out_11_qs;
      end

      addr_hit[64]: begin
        reg_rdata_next[31:0] = error_pos_out_12_qs;
      end

      addr_hit[65]: begin
        reg_rdata_next[31:0] = error_pos_out_13_qs;
      end

      addr_hit[66]: begin
        reg_rdata_next[31:0] = error_pos_out_14_qs;
      end

      addr_hit[67]: begin
        reg_rdata_next[31:0] = error_pos_out_15_qs;
      end

      addr_hit[68]: begin
        reg_rdata_next[31:0] = error_pos_out_16_qs;
      end

      addr_hit[69]: begin
        reg_rdata_next[31:0] = error_pos_out_17_qs;
      end

      addr_hit[70]: begin
        reg_rdata_next[31:0] = error_pos_out_18_qs;
      end

      addr_hit[71]: begin
        reg_rdata_next[31:0] = error_pos_out_19_qs;
      end

      addr_hit[72]: begin
        reg_rdata_next[31:0] = error_pos_out_20_qs;
      end

      addr_hit[73]: begin
        reg_rdata_next[31:0] = error_pos_out_21_qs;
      end

      addr_hit[74]: begin
        reg_rdata_next[31:0] = error_pos_out_22_qs;
      end

      addr_hit[75]: begin
        reg_rdata_next[31:0] = error_pos_out_23_qs;
      end

      addr_hit[76]: begin
        reg_rdata_next[31:0] = error_pos_out_24_qs;
      end

      addr_hit[77]: begin
        reg_rdata_next[31:0] = error_pos_out_25_qs;
      end

      addr_hit[78]: begin
        reg_rdata_next[31:0] = error_pos_out_26_qs;
      end

      addr_hit[79]: begin
        reg_rdata_next[31:0] = error_pos_out_27_qs;
      end

      addr_hit[80]: begin
        reg_rdata_next[31:0] = error_pos_out_28_qs;
      end

      addr_hit[81]: begin
        reg_rdata_next[31:0] = error_pos_out_29_qs;
      end

      addr_hit[82]: begin
        reg_rdata_next[31:0] = error_pos_out_30_qs;
      end

      addr_hit[83]: begin
        reg_rdata_next[31:0] = error_pos_out_31_qs;
      end

      addr_hit[84]: begin
        reg_rdata_next[31:0] = error_pos_out_32_qs;
      end

      addr_hit[85]: begin
        reg_rdata_next[31:0] = error_pos_out_33_qs;
      end

      addr_hit[86]: begin
        reg_rdata_next[31:0] = error_pos_out_34_qs;
      end

      addr_hit[87]: begin
        reg_rdata_next[31:0] = error_pos_out_35_qs;
      end

      addr_hit[88]: begin
        reg_rdata_next[31:0] = error_pos_out_36_qs;
      end

      addr_hit[89]: begin
        reg_rdata_next[31:0] = error_pos_out_37_qs;
      end

      addr_hit[90]: begin
        reg_rdata_next[31:0] = error_pos_out_38_qs;
      end

      addr_hit[91]: begin
        reg_rdata_next[31:0] = error_pos_out_39_qs;
      end

      addr_hit[92]: begin
        reg_rdata_next[31:0] = error_pos_out_40_qs;
      end

      addr_hit[93]: begin
        reg_rdata_next[31:0] = error_pos_out_41_qs;
      end

      addr_hit[94]: begin
        reg_rdata_next[31:0] = error_pos_out_42_qs;
      end

      addr_hit[95]: begin
        reg_rdata_next[31:0] = error_pos_out_43_qs;
      end

      addr_hit[96]: begin
        reg_rdata_next[31:0] = error_pos_out_44_qs;
      end

      addr_hit[97]: begin
        reg_rdata_next[31:0] = error_pos_out_45_qs;
      end

      addr_hit[98]: begin
        reg_rdata_next[31:0] = error_pos_out_46_qs;
      end

      addr_hit[99]: begin
        reg_rdata_next[31:0] = error_pos_out_47_qs;
      end

      addr_hit[100]: begin
        reg_rdata_next[31:0] = error_pos_out_48_qs;
      end

      addr_hit[101]: begin
        reg_rdata_next[31:0] = error_pos_out_49_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


`include "prim_assert.sv"

module rs_decode
  import rs_decode_reg_pkg::*;
(
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  input  logic                                      scan_mode,
  // Bus interface
  input  tlul_pkg::tl_h2d_t                         tl_i,
  output tlul_pkg::tl_d2h_t                         tl_o
);

  rs_decode_reg2hw_t               reg2hw;
  rs_decode_hw2reg_t               hw2reg;
  //wire                       ready_out;

  rs_decode_reg_top  u_rs_decode_reg_top (
    .clk_i                             ( clk_i           ),
    .rst_ni                            ( rst_ni          ),
    .tl_i                              ( tl_i            ),
    .hw2reg                            ( hw2reg          ),
    .devmode_i                         ( 1'b1            ),

    .tl_o                              ( tl_o            ),
    .reg2hw                            ( reg2hw          ),
    .intg_err_o                        (                 )
);

assign hw2reg.ctrl_signals.decode_en.de = 1'd0;
assign hw2reg.ctrl_signals.clrn.de = 1'd0;
always_comb begin
  for (int i = 0; i < 50; i++) begin
    hw2reg.encoded_data_in[i].de = 1'd0;
  end
end


  rs_decode_wrapper  u_rs_decode_wrapper (
    .clk                     ( clk_i        ),
    .rst_n                   ( rst_ni       ),
    .decode_en               ( reg2hw.ctrl_signals.decode_en.q),
    .clrn                    ( reg2hw.ctrl_signals.clrn.q ),
    .scan_mode               (scan_mode),
    .encoded_data            ( {reg2hw.encoded_data_in[49].q,reg2hw.encoded_data_in[48].q,reg2hw.encoded_data_in[47].q,reg2hw.encoded_data_in[46].q,reg2hw.encoded_data_in[45].q,reg2hw.encoded_data_in[44].q,reg2hw.encoded_data_in[43].q,reg2hw.encoded_data_in[42].q,reg2hw.encoded_data_in[41].q,reg2hw.encoded_data_in[40].q,reg2hw.encoded_data_in[39].q,reg2hw.encoded_data_in[38].q,reg2hw.encoded_data_in[37].q,reg2hw.encoded_data_in[36].q,reg2hw.encoded_data_in[35].q,reg2hw.encoded_data_in[34].q,reg2hw.encoded_data_in[33].q,reg2hw.encoded_data_in[32].q,reg2hw.encoded_data_in[31].q,reg2hw.encoded_data_in[30].q,reg2hw.encoded_data_in[29].q,reg2hw.encoded_data_in[28].q,reg2hw.encoded_data_in[27].q,reg2hw.encoded_data_in[26].q,reg2hw.encoded_data_in[25].q,reg2hw.encoded_data_in[24].q,reg2hw.encoded_data_in[23].q,reg2hw.encoded_data_in[22].q,reg2hw.encoded_data_in[21].q,reg2hw.encoded_data_in[20].q,reg2hw.encoded_data_in[19].q,reg2hw.encoded_data_in[18].q,reg2hw.encoded_data_in[17].q,reg2hw.encoded_data_in[16].q,reg2hw.encoded_data_in[15].q,reg2hw.encoded_data_in[14].q,reg2hw.encoded_data_in[13].q,reg2hw.encoded_data_in[12].q,reg2hw.encoded_data_in[11].q,reg2hw.encoded_data_in[10].q,reg2hw.encoded_data_in[9].q,reg2hw.encoded_data_in[8].q,reg2hw.encoded_data_in[7].q,reg2hw.encoded_data_in[6].q,reg2hw.encoded_data_in[5].q,reg2hw.encoded_data_in[4].q,reg2hw.encoded_data_in[3].q,reg2hw.encoded_data_in[2].q,reg2hw.encoded_data_in[1].q,reg2hw.encoded_data_in[0].q} ),

    .error_pos               ( {hw2reg.error_pos_out[49].d,hw2reg.error_pos_out[48].d,hw2reg.error_pos_out[47].d,hw2reg.error_pos_out[46].d,hw2reg.error_pos_out[45].d,hw2reg.error_pos_out[44].d,hw2reg.error_pos_out[43].d,hw2reg.error_pos_out[42].d,hw2reg.error_pos_out[41].d,hw2reg.error_pos_out[40].d,hw2reg.error_pos_out[39].d,hw2reg.error_pos_out[38].d,hw2reg.error_pos_out[37].d,hw2reg.error_pos_out[36].d,hw2reg.error_pos_out[35].d,hw2reg.error_pos_out[34].d,hw2reg.error_pos_out[33].d,hw2reg.error_pos_out[32].d,hw2reg.error_pos_out[31].d,hw2reg.error_pos_out[30].d,hw2reg.error_pos_out[29].d,hw2reg.error_pos_out[28].d,hw2reg.error_pos_out[27].d,hw2reg.error_pos_out[26].d,hw2reg.error_pos_out[25].d,hw2reg.error_pos_out[24].d,hw2reg.error_pos_out[23].d,hw2reg.error_pos_out[22].d,hw2reg.error_pos_out[21].d,hw2reg.error_pos_out[20].d,hw2reg.error_pos_out[19].d,hw2reg.error_pos_out[18].d,hw2reg.error_pos_out[17].d,hw2reg.error_pos_out[16].d,hw2reg.error_pos_out[15].d,hw2reg.error_pos_out[14].d,hw2reg.error_pos_out[13].d,hw2reg.error_pos_out[12].d,hw2reg.error_pos_out[11].d,hw2reg.error_pos_out[10].d,hw2reg.error_pos_out[9].d,hw2reg.error_pos_out[8].d,hw2reg.error_pos_out[7].d,hw2reg.error_pos_out[6].d,hw2reg.error_pos_out[5].d,hw2reg.error_pos_out[4].d,hw2reg.error_pos_out[3].d,hw2reg.error_pos_out[2].d,hw2reg.error_pos_out[1].d,hw2reg.error_pos_out[0].d} ),
    .output_valid            ( hw2reg.state_signals.output_valid_bit.d ),
    .ready                   ( hw2reg.state_signals.ready_bit.d ),
    .with_error              ( hw2reg.state_signals.with_error_bit.d ),
    .ready_re                ( hw2reg.state_signals.ready_bit.de ),
    .output_valid_re         ( hw2reg.state_signals.output_valid_bit.de ),
    .error_pos_re            ( {hw2reg.error_pos_out[49].de,hw2reg.error_pos_out[48].de,hw2reg.error_pos_out[47].de,hw2reg.error_pos_out[46].de,hw2reg.error_pos_out[45].de,hw2reg.error_pos_out[44].de,hw2reg.error_pos_out[43].de,hw2reg.error_pos_out[42].de,hw2reg.error_pos_out[41].de,hw2reg.error_pos_out[40].de,hw2reg.error_pos_out[39].de,hw2reg.error_pos_out[38].de,hw2reg.error_pos_out[37].de,hw2reg.error_pos_out[36].de,hw2reg.error_pos_out[35].de,hw2reg.error_pos_out[34].de,hw2reg.error_pos_out[33].de,hw2reg.error_pos_out[32].de,hw2reg.error_pos_out[31].de,hw2reg.error_pos_out[30].de,hw2reg.error_pos_out[29].de,hw2reg.error_pos_out[28].de,hw2reg.error_pos_out[27].de,hw2reg.error_pos_out[26].de,hw2reg.error_pos_out[25].de,hw2reg.error_pos_out[24].de,hw2reg.error_pos_out[23].de,hw2reg.error_pos_out[22].de,hw2reg.error_pos_out[21].de,hw2reg.error_pos_out[20].de,hw2reg.error_pos_out[19].de,hw2reg.error_pos_out[18].de,hw2reg.error_pos_out[17].de,hw2reg.error_pos_out[16].de,hw2reg.error_pos_out[15].de,hw2reg.error_pos_out[14].de,hw2reg.error_pos_out[13].de,hw2reg.error_pos_out[12].de,hw2reg.error_pos_out[11].de,hw2reg.error_pos_out[10].de,hw2reg.error_pos_out[9].de,hw2reg.error_pos_out[8].de,hw2reg.error_pos_out[7].de,hw2reg.error_pos_out[6].de,hw2reg.error_pos_out[5].de,hw2reg.error_pos_out[4].de,hw2reg.error_pos_out[3].de,hw2reg.error_pos_out[2].de,hw2reg.error_pos_out[1].de,hw2reg.error_pos_out[0].de} ),
    .with_error_re           ( hw2reg.state_signals.with_error_bit.de )
); 

endmodule




module rs_decode_wrapper(
    input clk,
    input rst_n, // Active low reset
    input decode_en,
    input clrn,
    input scan_mode,
    input [200*8-1:0] encoded_data,
    output reg [200*8-1:0] error_pos,
    output reg output_valid,
    output reg ready,
    output  with_error,  //output reg  with_error 
    
    output  ready_re,
    output  output_valid_re,
    output  [49:0] error_pos_re,
    output  with_error_re
);

// State declaration
localparam [1:0]
    IDLE = 2'b00,
    DECODE = 2'b01,
    COLLECT_ERROR = 2'b10,
    COMPLETE = 2'b11;

// Internal signals
reg [7:0] received;
reg dec_ena;
wire [7:0] error;
wire valid;
reg [11:0] bit_count;
reg [1:0] state, next_state;
reg [7:0] decode_counter; // Counter to maintain dec_ena for k clock cycles

localparam [7:0] k = 8'd200;

assign ready_re = 1'b1;
assign output_valid_re = output_valid;
assign with_error_re = 1'b1;
assign error_pos_re = {50{output_valid}};

// Instantiate the rsdec decoder module
rsdec x2 (
    .x(received),
    .error(error),
    .with_error(with_error), // Assuming not used, connect it properly if required
    .enable(dec_ena), // Connect dec_ena signal
    .valid(valid),
    .k(k),
    .clk(clk),
    .clrn(rst_n & (clrn | scan_mode))
    // Other connections to rsdec if needed
);

// State machine transition and output logic
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= IDLE;
        bit_count <= 0;
        error_pos <= 0;
        output_valid <= 0;
        decode_counter <= 0;
        dec_ena <= 0;
        ready <= 1;
    end else if (!clrn) begin
        state <= IDLE;
        bit_count <= 0;
        error_pos <= 0;
        output_valid <= 0;
        decode_counter <= 0;
        dec_ena <= 0;
        ready <= 1;
    end else begin
        case (state)
            IDLE: begin
                if (decode_en) begin
                    state <= DECODE;
                    dec_ena <= 0; // Enable the decoder
                    decode_counter <= 0; // Reset the counter
                    bit_count <= 0;
                    ready <= 0;
                end
            end
            DECODE: begin
                if (decode_counter >= (k)) begin
                    dec_ena <= 0;
                end else begin
                    dec_ena <= 1;
                    received <= encoded_data[decode_counter*8 +: 8]; // Grab the next byte of input data
                    decode_counter <= decode_counter + 1; // Increment counter
                end

                if (!dec_ena && with_error) begin
                    state <= COLLECT_ERROR;
                    decode_counter <= 0;
                end
            end
            COLLECT_ERROR: begin
                if (valid) begin
                    error_pos[bit_count*8 +: 8] <= error; // Collect error data
                    bit_count <= bit_count + 1; // Increment bit_count to point to the next byte
                    if (bit_count >= k-1) begin // Check if all bytes processed
                        state <= COMPLETE;
                    end
                end else begin
                    state <= COLLECT_ERROR; // Transition to complete once valid goes low
                end
            end
            COMPLETE: begin
                output_valid <= 1; // Indicate that the output data is valid
                state <= IDLE; // Reset to idle state for the next operation
                bit_count <= 0; // Reset bit_count for the next operation
                ready <= 1;
            end
            default: state <= IDLE;
        endcase
    end
end

endmodule



// -------------------------------------------------------------------------
//Reed-Solomon Encoder
//Copyright (C) Tue Apr  2 17:06:57 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module rs_enc_m0 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[5] ^ x[6];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3] ^ x[4];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[4] ^ x[5] ^ x[7];
	end
endmodule

module rs_enc_m1 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[4] ^ x[5];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[6];
		y[2] = x[0] ^ x[7];
		y[3] = x[1];
		y[4] = x[0] ^ x[2];
		y[5] = x[0] ^ x[1] ^ x[3];
		y[6] = x[1] ^ x[2] ^ x[4];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[4];
	end
endmodule

module rs_enc_m2 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[1] = x[0] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[3] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[4] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
	end
endmodule

module rs_enc_m3 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3];
		y[3] = x[1] ^ x[2] ^ x[4];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[5];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[6];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[1] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rs_enc_m4 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[5] ^ x[7];
		y[1] = x[2] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[5] = x[2] ^ x[3] ^ x[4] ^ x[6];
		y[6] = x[0] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[0] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rs_enc_m5 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[4];
		y[1] = x[0] ^ x[2] ^ x[4] ^ x[5];
		y[2] = x[3] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[1] ^ x[2] ^ x[6] ^ x[7];
		y[6] = x[0] ^ x[2] ^ x[3] ^ x[7];
		y[7] = x[0] ^ x[3];
	end
endmodule

module rs_enc_m6 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[3] ^ x[4];
		y[2] = x[2] ^ x[6] ^ x[7];
		y[3] = x[3] ^ x[7];
		y[4] = x[0] ^ x[4];
		y[5] = x[0] ^ x[1] ^ x[5];
		y[6] = x[1] ^ x[2] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
	end
endmodule

module rs_enc_m7 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[2] = x[4] ^ x[7];
		y[3] = x[0] ^ x[5];
		y[4] = x[0] ^ x[1] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[3];
		y[7] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rs_enc_m8 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[6];
		y[1] = x[2] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[3] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[4] ^ x[7];
		y[4] = x[2] ^ x[3] ^ x[5];
		y[5] = x[3] ^ x[4] ^ x[6];
		y[6] = x[0] ^ x[4] ^ x[5] ^ x[7];
		y[7] = x[0] ^ x[5];
	end
endmodule

module rs_enc_m9 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[5] ^ x[7];
		y[1] = x[1] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[4] ^ x[5] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[3] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
		y[6] = x[1] ^ x[3] ^ x[4] ^ x[5];
		y[7] = x[0] ^ x[1] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rs_enc_m10 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[4] ^ x[7];
		y[1] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[7];
		y[4] = x[1] ^ x[3] ^ x[4];
		y[5] = x[0] ^ x[2] ^ x[4] ^ x[5];
		y[6] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[3] ^ x[6];
	end
endmodule

module rs_enc_m11 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[1] = x[2] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[4];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[5];
		y[4] = x[1] ^ x[2] ^ x[4] ^ x[6];
		y[5] = x[2] ^ x[3] ^ x[5] ^ x[7];
		y[6] = x[0] ^ x[3] ^ x[4] ^ x[6];
		y[7] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6];
	end
endmodule

module rs_enc_m12 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4];
		y[2] = x[2] ^ x[4] ^ x[5];
		y[3] = x[3] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[5] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[7];
	end
endmodule

module rs_enc_m13 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[2] ^ x[3] ^ x[6] ^ x[7];
		y[1] = x[2] ^ x[4] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[5] ^ x[6];
		y[3] = x[1] ^ x[3] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[4] ^ x[7];
		y[5] = x[1] ^ x[3] ^ x[5];
		y[6] = x[0] ^ x[2] ^ x[4] ^ x[6];
		y[7] = x[1] ^ x[2] ^ x[5] ^ x[6];
	end
endmodule

module rs_enc_m14 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[5];
		y[1] = x[1] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[4] ^ x[7];
		y[5] = x[2] ^ x[3] ^ x[5];
		y[6] = x[3] ^ x[4] ^ x[6];
		y[7] = x[4] ^ x[7];
	end
endmodule

module rs_enc_m15 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[1] = x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[4] = x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6];
	end
endmodule

module rs_enc_m16 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[1];
		y[2] = x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[5] ^ x[6] ^ x[7];
		y[5] = x[6] ^ x[7];
		y[6] = x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
	end
endmodule

module rs_enc_m17 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[5];
		y[1] = x[1] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[6] ^ x[7];
		y[4] = x[1] ^ x[2] ^ x[4] ^ x[7];
		y[5] = x[2] ^ x[3] ^ x[5];
		y[6] = x[3] ^ x[4] ^ x[6];
		y[7] = x[4] ^ x[7];
	end
endmodule

module rs_enc_m18 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3] ^ x[5];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[3] ^ x[5] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[4] ^ x[7];
	end
endmodule

module rs_enc_m19 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[1] = x[3] ^ x[4] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[6];
		y[3] = x[2] ^ x[3] ^ x[7];
		y[4] = x[0] ^ x[3] ^ x[4];
		y[5] = x[0] ^ x[1] ^ x[4] ^ x[5];
		y[6] = x[1] ^ x[2] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
	end
endmodule

module rs_enc_m20 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[6];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[5] ^ x[7];
	end
endmodule

module rs_enc_m21 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[3] ^ x[5];
		y[2] = x[2] ^ x[4] ^ x[5] ^ x[7];
		y[3] = x[0] ^ x[3] ^ x[5] ^ x[6];
		y[4] = x[1] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[2] ^ x[5] ^ x[7];
		y[6] = x[1] ^ x[3] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[4] ^ x[5] ^ x[6];
	end
endmodule

module rs_enc_m22 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[7];
		y[1] = x[3] ^ x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2];
		y[3] = x[1] ^ x[2] ^ x[3];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4];
		y[5] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5];
		y[6] = x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[6];
	end
endmodule

module rs_enc_m23 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6];
		y[1] = x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[3];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[4];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5];
		y[5] = x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5] ^ x[7];
	end
endmodule

module rs_enc_m24 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[1] = x[2] ^ x[3] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[5];
		y[3] = x[1] ^ x[2] ^ x[6];
		y[4] = x[2] ^ x[3] ^ x[7];
		y[5] = x[0] ^ x[3] ^ x[4];
		y[6] = x[0] ^ x[1] ^ x[4] ^ x[5];
		y[7] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
	end
endmodule

module rs_enc_m25 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[7];
		y[1] = x[3] ^ x[4] ^ x[5] ^ x[7];
		y[2] = x[1] ^ x[2] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[2] ^ x[3] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[4] ^ x[5];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6];
		y[7] = x[0] ^ x[1] ^ x[3] ^ x[6];
	end
endmodule

module rs_enc_m26 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[3] ^ x[5];
		y[1] = x[3] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[7];
		y[7] = x[2] ^ x[4];
	end
endmodule

module rs_enc_m27 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[3];
		y[1] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4];
		y[2] = x[2] ^ x[4] ^ x[5];
		y[3] = x[3] ^ x[5] ^ x[6];
		y[4] = x[0] ^ x[4] ^ x[6] ^ x[7];
		y[5] = x[0] ^ x[1] ^ x[5] ^ x[7];
		y[6] = x[0] ^ x[1] ^ x[2] ^ x[6];
		y[7] = x[0] ^ x[2] ^ x[7];
	end
endmodule

module rs_enc_m28 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6] ^ x[7];
		y[1] = x[0] ^ x[4] ^ x[6];
		y[2] = x[0] ^ x[2] ^ x[3] ^ x[5] ^ x[6];
		y[3] = x[1] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[1] ^ x[3] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[4] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[6];
	end
endmodule

module rs_enc_m29 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[1] ^ x[2] ^ x[3] ^ x[5];
		y[1] = x[0] ^ x[1] ^ x[4] ^ x[5] ^ x[6];
		y[2] = x[0] ^ x[3] ^ x[6] ^ x[7];
		y[3] = x[0] ^ x[1] ^ x[4] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[5];
		y[5] = x[1] ^ x[2] ^ x[3] ^ x[6];
		y[6] = x[2] ^ x[3] ^ x[4] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[4];
	end
endmodule

module rs_enc_m30 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[3] ^ x[5] ^ x[7];
		y[1] = x[0] ^ x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6];
		y[3] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[4] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[5] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[6] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[2] ^ x[4] ^ x[6];
	end
endmodule

module rs_enc_m31 (y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;
	always @ (x)
	begin
		y[0] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[6];
		y[1] = x[4] ^ x[6] ^ x[7];
		y[2] = x[0] ^ x[1] ^ x[2] ^ x[3] ^ x[5] ^ x[6] ^ x[7];
		y[3] = x[1] ^ x[2] ^ x[3] ^ x[4] ^ x[6] ^ x[7];
		y[4] = x[0] ^ x[2] ^ x[3] ^ x[4] ^ x[5] ^ x[7];
		y[5] = x[1] ^ x[3] ^ x[4] ^ x[5] ^ x[6];
		y[6] = x[2] ^ x[4] ^ x[5] ^ x[6] ^ x[7];
		y[7] = x[0] ^ x[1] ^ x[2] ^ x[5] ^ x[7];
	end
endmodule

module rs_enc (y, x, enable, data, clk, clrn);
	input [7:0] x;
	input clk, clrn, enable, data;
	output [7:0] y;
	reg [7:0] y;

	wire [7:0] scale0;
	wire [7:0] scale1;
	wire [7:0] scale2;
	wire [7:0] scale3;
	wire [7:0] scale4;
	wire [7:0] scale5;
	wire [7:0] scale6;
	wire [7:0] scale7;
	wire [7:0] scale8;
	wire [7:0] scale9;
	wire [7:0] scale10;
	wire [7:0] scale11;
	wire [7:0] scale12;
	wire [7:0] scale13;
	wire [7:0] scale14;
	wire [7:0] scale15;
	wire [7:0] scale16;
	wire [7:0] scale17;
	wire [7:0] scale18;
	wire [7:0] scale19;
	wire [7:0] scale20;
	wire [7:0] scale21;
	wire [7:0] scale22;
	wire [7:0] scale23;
	wire [7:0] scale24;
	wire [7:0] scale25;
	wire [7:0] scale26;
	wire [7:0] scale27;
	wire [7:0] scale28;
	wire [7:0] scale29;
	wire [7:0] scale30;
	wire [7:0] scale31;
	reg [7:0] mem0;
	reg [7:0] mem1;
	reg [7:0] mem2;
	reg [7:0] mem3;
	reg [7:0] mem4;
	reg [7:0] mem5;
	reg [7:0] mem6;
	reg [7:0] mem7;
	reg [7:0] mem8;
	reg [7:0] mem9;
	reg [7:0] mem10;
	reg [7:0] mem11;
	reg [7:0] mem12;
	reg [7:0] mem13;
	reg [7:0] mem14;
	reg [7:0] mem15;
	reg [7:0] mem16;
	reg [7:0] mem17;
	reg [7:0] mem18;
	reg [7:0] mem19;
	reg [7:0] mem20;
	reg [7:0] mem21;
	reg [7:0] mem22;
	reg [7:0] mem23;
	reg [7:0] mem24;
	reg [7:0] mem25;
	reg [7:0] mem26;
	reg [7:0] mem27;
	reg [7:0] mem28;
	reg [7:0] mem29;
	reg [7:0] mem30;
	reg [7:0] mem31;
	reg [7:0] feedback;

	rs_enc_m0 m0 (scale0, feedback);
	rs_enc_m1 m1 (scale1, feedback);
	rs_enc_m2 m2 (scale2, feedback);
	rs_enc_m3 m3 (scale3, feedback);
	rs_enc_m4 m4 (scale4, feedback);
	rs_enc_m5 m5 (scale5, feedback);
	rs_enc_m6 m6 (scale6, feedback);
	rs_enc_m7 m7 (scale7, feedback);
	rs_enc_m8 m8 (scale8, feedback);
	rs_enc_m9 m9 (scale9, feedback);
	rs_enc_m10 m10 (scale10, feedback);
	rs_enc_m11 m11 (scale11, feedback);
	rs_enc_m12 m12 (scale12, feedback);
	rs_enc_m13 m13 (scale13, feedback);
	rs_enc_m14 m14 (scale14, feedback);
	rs_enc_m15 m15 (scale15, feedback);
	rs_enc_m16 m16 (scale16, feedback);
	rs_enc_m17 m17 (scale17, feedback);
	rs_enc_m18 m18 (scale18, feedback);
	rs_enc_m19 m19 (scale19, feedback);
	rs_enc_m20 m20 (scale20, feedback);
	rs_enc_m21 m21 (scale21, feedback);
	rs_enc_m22 m22 (scale22, feedback);
	rs_enc_m23 m23 (scale23, feedback);
	rs_enc_m24 m24 (scale24, feedback);
	rs_enc_m25 m25 (scale25, feedback);
	rs_enc_m26 m26 (scale26, feedback);
	rs_enc_m27 m27 (scale27, feedback);
	rs_enc_m28 m28 (scale28, feedback);
	rs_enc_m29 m29 (scale29, feedback);
	rs_enc_m30 m30 (scale30, feedback);
	rs_enc_m31 m31 (scale31, feedback);

	always @ (posedge clk or negedge clrn)
	begin
		if (~clrn)
		begin
			mem0 <= 0;
			mem1 <= 0;
			mem2 <= 0;
			mem3 <= 0;
			mem4 <= 0;
			mem5 <= 0;
			mem6 <= 0;
			mem7 <= 0;
			mem8 <= 0;
			mem9 <= 0;
			mem10 <= 0;
			mem11 <= 0;
			mem12 <= 0;
			mem13 <= 0;
			mem14 <= 0;
			mem15 <= 0;
			mem16 <= 0;
			mem17 <= 0;
			mem18 <= 0;
			mem19 <= 0;
			mem20 <= 0;
			mem21 <= 0;
			mem22 <= 0;
			mem23 <= 0;
			mem24 <= 0;
			mem25 <= 0;
			mem26 <= 0;
			mem27 <= 0;
			mem28 <= 0;
			mem29 <= 0;
			mem30 <= 0;
			mem31 <= 0;
		end
		else if (enable)
		begin
			mem31 <= mem30 ^ scale31;
			mem30 <= mem29 ^ scale30;
			mem29 <= mem28 ^ scale29;
			mem28 <= mem27 ^ scale28;
			mem27 <= mem26 ^ scale27;
			mem26 <= mem25 ^ scale26;
			mem25 <= mem24 ^ scale25;
			mem24 <= mem23 ^ scale24;
			mem23 <= mem22 ^ scale23;
			mem22 <= mem21 ^ scale22;
			mem21 <= mem20 ^ scale21;
			mem20 <= mem19 ^ scale20;
			mem19 <= mem18 ^ scale19;
			mem18 <= mem17 ^ scale18;
			mem17 <= mem16 ^ scale17;
			mem16 <= mem15 ^ scale16;
			mem15 <= mem14 ^ scale15;
			mem14 <= mem13 ^ scale14;
			mem13 <= mem12 ^ scale13;
			mem12 <= mem11 ^ scale12;
			mem11 <= mem10 ^ scale11;
			mem10 <= mem9 ^ scale10;
			mem9 <= mem8 ^ scale9;
			mem8 <= mem7 ^ scale8;
			mem7 <= mem6 ^ scale7;
			mem6 <= mem5 ^ scale6;
			mem5 <= mem4 ^ scale5;
			mem4 <= mem3 ^ scale4;
			mem3 <= mem2 ^ scale3;
			mem2 <= mem1 ^ scale2;
			mem1 <= mem0 ^ scale1;
			mem0 <= scale0;
		end
	end

	always @ (data or x or mem31)
		if (data) feedback = x ^ mem31;
		else feedback = 0;

	always @ (data or x or mem31)
		if (data) y = x;
		else y = mem31;

endmodule


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package rs_encode_reg_pkg;

  // Param list
  parameter int NumRegs_Data_in = 42;
  parameter int NumRegs_encoded_data = 50;

  // Address widths within the block
  parameter int BlockAw = 9;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    struct packed {
      logic        q;
      logic        qe;
    } encode_en;
    struct packed {
      logic        q;
      logic        qe;
    } clrn;
  } rs_encode_reg2hw_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        q;
    } valid_bit;
    struct packed {
      logic        q;
    } ready_bit;
  } rs_encode_reg2hw_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] q;
    logic        qe;
  } rs_encode_reg2hw_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] q;
  } rs_encode_reg2hw_encoded_data_out_mreg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } encode_en;
    struct packed {
      logic        d;
      logic        de;
    } clrn;
  } rs_encode_hw2reg_ctrl_signals_reg_t;

  typedef struct packed {
    struct packed {
      logic        d;
      logic        de;
    } valid_bit;
    struct packed {
      logic        d;
      logic        de;
    } ready_bit;
  } rs_encode_hw2reg_state_signals_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } rs_encode_hw2reg_data_in_mreg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } rs_encode_hw2reg_encoded_data_out_mreg_t;

  // Register -> HW type
  typedef struct packed {
    rs_encode_reg2hw_ctrl_signals_reg_t ctrl_signals; // [2991:2988]
    rs_encode_reg2hw_state_signals_reg_t state_signals; // [2987:2986]
    rs_encode_reg2hw_data_in_mreg_t [41:0] data_in; // [2985:1600]
    rs_encode_reg2hw_encoded_data_out_mreg_t [49:0] encoded_data_out; // [1599:0]
  } rs_encode_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    rs_encode_hw2reg_ctrl_signals_reg_t ctrl_signals; // [3043:3040]
    rs_encode_hw2reg_state_signals_reg_t state_signals; // [3039:3036]
    rs_encode_hw2reg_data_in_mreg_t [41:0] data_in; // [3035:1650]
    rs_encode_hw2reg_encoded_data_out_mreg_t [49:0] encoded_data_out; // [1649:0]
  } rs_encode_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] RS_ENCODE_CTRL_SIGNALS_OFFSET = 9'h 0;
  parameter logic [BlockAw-1:0] RS_ENCODE_STATE_SIGNALS_OFFSET = 9'h 4;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_0_OFFSET = 9'h 8;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_1_OFFSET = 9'h c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_2_OFFSET = 9'h 10;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_3_OFFSET = 9'h 14;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_4_OFFSET = 9'h 18;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_5_OFFSET = 9'h 1c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_6_OFFSET = 9'h 20;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_7_OFFSET = 9'h 24;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_8_OFFSET = 9'h 28;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_9_OFFSET = 9'h 2c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_10_OFFSET = 9'h 30;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_11_OFFSET = 9'h 34;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_12_OFFSET = 9'h 38;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_13_OFFSET = 9'h 3c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_14_OFFSET = 9'h 40;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_15_OFFSET = 9'h 44;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_16_OFFSET = 9'h 48;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_17_OFFSET = 9'h 4c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_18_OFFSET = 9'h 50;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_19_OFFSET = 9'h 54;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_20_OFFSET = 9'h 58;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_21_OFFSET = 9'h 5c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_22_OFFSET = 9'h 60;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_23_OFFSET = 9'h 64;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_24_OFFSET = 9'h 68;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_25_OFFSET = 9'h 6c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_26_OFFSET = 9'h 70;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_27_OFFSET = 9'h 74;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_28_OFFSET = 9'h 78;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_29_OFFSET = 9'h 7c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_30_OFFSET = 9'h 80;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_31_OFFSET = 9'h 84;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_32_OFFSET = 9'h 88;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_33_OFFSET = 9'h 8c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_34_OFFSET = 9'h 90;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_35_OFFSET = 9'h 94;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_36_OFFSET = 9'h 98;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_37_OFFSET = 9'h 9c;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_38_OFFSET = 9'h a0;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_39_OFFSET = 9'h a4;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_40_OFFSET = 9'h a8;
  parameter logic [BlockAw-1:0] RS_ENCODE_DATA_IN_41_OFFSET = 9'h ac;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_0_OFFSET = 9'h b0;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_1_OFFSET = 9'h b4;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_2_OFFSET = 9'h b8;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_3_OFFSET = 9'h bc;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_4_OFFSET = 9'h c0;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_5_OFFSET = 9'h c4;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_6_OFFSET = 9'h c8;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_7_OFFSET = 9'h cc;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_8_OFFSET = 9'h d0;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_9_OFFSET = 9'h d4;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_10_OFFSET = 9'h d8;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_11_OFFSET = 9'h dc;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_12_OFFSET = 9'h e0;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_13_OFFSET = 9'h e4;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_14_OFFSET = 9'h e8;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_15_OFFSET = 9'h ec;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_16_OFFSET = 9'h f0;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_17_OFFSET = 9'h f4;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_18_OFFSET = 9'h f8;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_19_OFFSET = 9'h fc;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_20_OFFSET = 9'h 100;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_21_OFFSET = 9'h 104;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_22_OFFSET = 9'h 108;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_23_OFFSET = 9'h 10c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_24_OFFSET = 9'h 110;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_25_OFFSET = 9'h 114;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_26_OFFSET = 9'h 118;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_27_OFFSET = 9'h 11c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_28_OFFSET = 9'h 120;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_29_OFFSET = 9'h 124;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_30_OFFSET = 9'h 128;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_31_OFFSET = 9'h 12c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_32_OFFSET = 9'h 130;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_33_OFFSET = 9'h 134;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_34_OFFSET = 9'h 138;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_35_OFFSET = 9'h 13c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_36_OFFSET = 9'h 140;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_37_OFFSET = 9'h 144;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_38_OFFSET = 9'h 148;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_39_OFFSET = 9'h 14c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_40_OFFSET = 9'h 150;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_41_OFFSET = 9'h 154;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_42_OFFSET = 9'h 158;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_43_OFFSET = 9'h 15c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_44_OFFSET = 9'h 160;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_45_OFFSET = 9'h 164;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_46_OFFSET = 9'h 168;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_47_OFFSET = 9'h 16c;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_48_OFFSET = 9'h 170;
  parameter logic [BlockAw-1:0] RS_ENCODE_ENCODED_DATA_OUT_49_OFFSET = 9'h 174;

  // Register index
  typedef enum int {
    RS_ENCODE_CTRL_SIGNALS,
    RS_ENCODE_STATE_SIGNALS,
    RS_ENCODE_DATA_IN_0,
    RS_ENCODE_DATA_IN_1,
    RS_ENCODE_DATA_IN_2,
    RS_ENCODE_DATA_IN_3,
    RS_ENCODE_DATA_IN_4,
    RS_ENCODE_DATA_IN_5,
    RS_ENCODE_DATA_IN_6,
    RS_ENCODE_DATA_IN_7,
    RS_ENCODE_DATA_IN_8,
    RS_ENCODE_DATA_IN_9,
    RS_ENCODE_DATA_IN_10,
    RS_ENCODE_DATA_IN_11,
    RS_ENCODE_DATA_IN_12,
    RS_ENCODE_DATA_IN_13,
    RS_ENCODE_DATA_IN_14,
    RS_ENCODE_DATA_IN_15,
    RS_ENCODE_DATA_IN_16,
    RS_ENCODE_DATA_IN_17,
    RS_ENCODE_DATA_IN_18,
    RS_ENCODE_DATA_IN_19,
    RS_ENCODE_DATA_IN_20,
    RS_ENCODE_DATA_IN_21,
    RS_ENCODE_DATA_IN_22,
    RS_ENCODE_DATA_IN_23,
    RS_ENCODE_DATA_IN_24,
    RS_ENCODE_DATA_IN_25,
    RS_ENCODE_DATA_IN_26,
    RS_ENCODE_DATA_IN_27,
    RS_ENCODE_DATA_IN_28,
    RS_ENCODE_DATA_IN_29,
    RS_ENCODE_DATA_IN_30,
    RS_ENCODE_DATA_IN_31,
    RS_ENCODE_DATA_IN_32,
    RS_ENCODE_DATA_IN_33,
    RS_ENCODE_DATA_IN_34,
    RS_ENCODE_DATA_IN_35,
    RS_ENCODE_DATA_IN_36,
    RS_ENCODE_DATA_IN_37,
    RS_ENCODE_DATA_IN_38,
    RS_ENCODE_DATA_IN_39,
    RS_ENCODE_DATA_IN_40,
    RS_ENCODE_DATA_IN_41,
    RS_ENCODE_ENCODED_DATA_OUT_0,
    RS_ENCODE_ENCODED_DATA_OUT_1,
    RS_ENCODE_ENCODED_DATA_OUT_2,
    RS_ENCODE_ENCODED_DATA_OUT_3,
    RS_ENCODE_ENCODED_DATA_OUT_4,
    RS_ENCODE_ENCODED_DATA_OUT_5,
    RS_ENCODE_ENCODED_DATA_OUT_6,
    RS_ENCODE_ENCODED_DATA_OUT_7,
    RS_ENCODE_ENCODED_DATA_OUT_8,
    RS_ENCODE_ENCODED_DATA_OUT_9,
    RS_ENCODE_ENCODED_DATA_OUT_10,
    RS_ENCODE_ENCODED_DATA_OUT_11,
    RS_ENCODE_ENCODED_DATA_OUT_12,
    RS_ENCODE_ENCODED_DATA_OUT_13,
    RS_ENCODE_ENCODED_DATA_OUT_14,
    RS_ENCODE_ENCODED_DATA_OUT_15,
    RS_ENCODE_ENCODED_DATA_OUT_16,
    RS_ENCODE_ENCODED_DATA_OUT_17,
    RS_ENCODE_ENCODED_DATA_OUT_18,
    RS_ENCODE_ENCODED_DATA_OUT_19,
    RS_ENCODE_ENCODED_DATA_OUT_20,
    RS_ENCODE_ENCODED_DATA_OUT_21,
    RS_ENCODE_ENCODED_DATA_OUT_22,
    RS_ENCODE_ENCODED_DATA_OUT_23,
    RS_ENCODE_ENCODED_DATA_OUT_24,
    RS_ENCODE_ENCODED_DATA_OUT_25,
    RS_ENCODE_ENCODED_DATA_OUT_26,
    RS_ENCODE_ENCODED_DATA_OUT_27,
    RS_ENCODE_ENCODED_DATA_OUT_28,
    RS_ENCODE_ENCODED_DATA_OUT_29,
    RS_ENCODE_ENCODED_DATA_OUT_30,
    RS_ENCODE_ENCODED_DATA_OUT_31,
    RS_ENCODE_ENCODED_DATA_OUT_32,
    RS_ENCODE_ENCODED_DATA_OUT_33,
    RS_ENCODE_ENCODED_DATA_OUT_34,
    RS_ENCODE_ENCODED_DATA_OUT_35,
    RS_ENCODE_ENCODED_DATA_OUT_36,
    RS_ENCODE_ENCODED_DATA_OUT_37,
    RS_ENCODE_ENCODED_DATA_OUT_38,
    RS_ENCODE_ENCODED_DATA_OUT_39,
    RS_ENCODE_ENCODED_DATA_OUT_40,
    RS_ENCODE_ENCODED_DATA_OUT_41,
    RS_ENCODE_ENCODED_DATA_OUT_42,
    RS_ENCODE_ENCODED_DATA_OUT_43,
    RS_ENCODE_ENCODED_DATA_OUT_44,
    RS_ENCODE_ENCODED_DATA_OUT_45,
    RS_ENCODE_ENCODED_DATA_OUT_46,
    RS_ENCODE_ENCODED_DATA_OUT_47,
    RS_ENCODE_ENCODED_DATA_OUT_48,
    RS_ENCODE_ENCODED_DATA_OUT_49
  } rs_encode_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] RS_ENCODE_PERMIT [94] = '{
    4'b 0001, // index[ 0] RS_ENCODE_CTRL_SIGNALS
    4'b 0001, // index[ 1] RS_ENCODE_STATE_SIGNALS
    4'b 1111, // index[ 2] RS_ENCODE_DATA_IN_0
    4'b 1111, // index[ 3] RS_ENCODE_DATA_IN_1
    4'b 1111, // index[ 4] RS_ENCODE_DATA_IN_2
    4'b 1111, // index[ 5] RS_ENCODE_DATA_IN_3
    4'b 1111, // index[ 6] RS_ENCODE_DATA_IN_4
    4'b 1111, // index[ 7] RS_ENCODE_DATA_IN_5
    4'b 1111, // index[ 8] RS_ENCODE_DATA_IN_6
    4'b 1111, // index[ 9] RS_ENCODE_DATA_IN_7
    4'b 1111, // index[10] RS_ENCODE_DATA_IN_8
    4'b 1111, // index[11] RS_ENCODE_DATA_IN_9
    4'b 1111, // index[12] RS_ENCODE_DATA_IN_10
    4'b 1111, // index[13] RS_ENCODE_DATA_IN_11
    4'b 1111, // index[14] RS_ENCODE_DATA_IN_12
    4'b 1111, // index[15] RS_ENCODE_DATA_IN_13
    4'b 1111, // index[16] RS_ENCODE_DATA_IN_14
    4'b 1111, // index[17] RS_ENCODE_DATA_IN_15
    4'b 1111, // index[18] RS_ENCODE_DATA_IN_16
    4'b 1111, // index[19] RS_ENCODE_DATA_IN_17
    4'b 1111, // index[20] RS_ENCODE_DATA_IN_18
    4'b 1111, // index[21] RS_ENCODE_DATA_IN_19
    4'b 1111, // index[22] RS_ENCODE_DATA_IN_20
    4'b 1111, // index[23] RS_ENCODE_DATA_IN_21
    4'b 1111, // index[24] RS_ENCODE_DATA_IN_22
    4'b 1111, // index[25] RS_ENCODE_DATA_IN_23
    4'b 1111, // index[26] RS_ENCODE_DATA_IN_24
    4'b 1111, // index[27] RS_ENCODE_DATA_IN_25
    4'b 1111, // index[28] RS_ENCODE_DATA_IN_26
    4'b 1111, // index[29] RS_ENCODE_DATA_IN_27
    4'b 1111, // index[30] RS_ENCODE_DATA_IN_28
    4'b 1111, // index[31] RS_ENCODE_DATA_IN_29
    4'b 1111, // index[32] RS_ENCODE_DATA_IN_30
    4'b 1111, // index[33] RS_ENCODE_DATA_IN_31
    4'b 1111, // index[34] RS_ENCODE_DATA_IN_32
    4'b 1111, // index[35] RS_ENCODE_DATA_IN_33
    4'b 1111, // index[36] RS_ENCODE_DATA_IN_34
    4'b 1111, // index[37] RS_ENCODE_DATA_IN_35
    4'b 1111, // index[38] RS_ENCODE_DATA_IN_36
    4'b 1111, // index[39] RS_ENCODE_DATA_IN_37
    4'b 1111, // index[40] RS_ENCODE_DATA_IN_38
    4'b 1111, // index[41] RS_ENCODE_DATA_IN_39
    4'b 1111, // index[42] RS_ENCODE_DATA_IN_40
    4'b 1111, // index[43] RS_ENCODE_DATA_IN_41
    4'b 1111, // index[44] RS_ENCODE_ENCODED_DATA_OUT_0
    4'b 1111, // index[45] RS_ENCODE_ENCODED_DATA_OUT_1
    4'b 1111, // index[46] RS_ENCODE_ENCODED_DATA_OUT_2
    4'b 1111, // index[47] RS_ENCODE_ENCODED_DATA_OUT_3
    4'b 1111, // index[48] RS_ENCODE_ENCODED_DATA_OUT_4
    4'b 1111, // index[49] RS_ENCODE_ENCODED_DATA_OUT_5
    4'b 1111, // index[50] RS_ENCODE_ENCODED_DATA_OUT_6
    4'b 1111, // index[51] RS_ENCODE_ENCODED_DATA_OUT_7
    4'b 1111, // index[52] RS_ENCODE_ENCODED_DATA_OUT_8
    4'b 1111, // index[53] RS_ENCODE_ENCODED_DATA_OUT_9
    4'b 1111, // index[54] RS_ENCODE_ENCODED_DATA_OUT_10
    4'b 1111, // index[55] RS_ENCODE_ENCODED_DATA_OUT_11
    4'b 1111, // index[56] RS_ENCODE_ENCODED_DATA_OUT_12
    4'b 1111, // index[57] RS_ENCODE_ENCODED_DATA_OUT_13
    4'b 1111, // index[58] RS_ENCODE_ENCODED_DATA_OUT_14
    4'b 1111, // index[59] RS_ENCODE_ENCODED_DATA_OUT_15
    4'b 1111, // index[60] RS_ENCODE_ENCODED_DATA_OUT_16
    4'b 1111, // index[61] RS_ENCODE_ENCODED_DATA_OUT_17
    4'b 1111, // index[62] RS_ENCODE_ENCODED_DATA_OUT_18
    4'b 1111, // index[63] RS_ENCODE_ENCODED_DATA_OUT_19
    4'b 1111, // index[64] RS_ENCODE_ENCODED_DATA_OUT_20
    4'b 1111, // index[65] RS_ENCODE_ENCODED_DATA_OUT_21
    4'b 1111, // index[66] RS_ENCODE_ENCODED_DATA_OUT_22
    4'b 1111, // index[67] RS_ENCODE_ENCODED_DATA_OUT_23
    4'b 1111, // index[68] RS_ENCODE_ENCODED_DATA_OUT_24
    4'b 1111, // index[69] RS_ENCODE_ENCODED_DATA_OUT_25
    4'b 1111, // index[70] RS_ENCODE_ENCODED_DATA_OUT_26
    4'b 1111, // index[71] RS_ENCODE_ENCODED_DATA_OUT_27
    4'b 1111, // index[72] RS_ENCODE_ENCODED_DATA_OUT_28
    4'b 1111, // index[73] RS_ENCODE_ENCODED_DATA_OUT_29
    4'b 1111, // index[74] RS_ENCODE_ENCODED_DATA_OUT_30
    4'b 1111, // index[75] RS_ENCODE_ENCODED_DATA_OUT_31
    4'b 1111, // index[76] RS_ENCODE_ENCODED_DATA_OUT_32
    4'b 1111, // index[77] RS_ENCODE_ENCODED_DATA_OUT_33
    4'b 1111, // index[78] RS_ENCODE_ENCODED_DATA_OUT_34
    4'b 1111, // index[79] RS_ENCODE_ENCODED_DATA_OUT_35
    4'b 1111, // index[80] RS_ENCODE_ENCODED_DATA_OUT_36
    4'b 1111, // index[81] RS_ENCODE_ENCODED_DATA_OUT_37
    4'b 1111, // index[82] RS_ENCODE_ENCODED_DATA_OUT_38
    4'b 1111, // index[83] RS_ENCODE_ENCODED_DATA_OUT_39
    4'b 1111, // index[84] RS_ENCODE_ENCODED_DATA_OUT_40
    4'b 1111, // index[85] RS_ENCODE_ENCODED_DATA_OUT_41
    4'b 1111, // index[86] RS_ENCODE_ENCODED_DATA_OUT_42
    4'b 1111, // index[87] RS_ENCODE_ENCODED_DATA_OUT_43
    4'b 1111, // index[88] RS_ENCODE_ENCODED_DATA_OUT_44
    4'b 1111, // index[89] RS_ENCODE_ENCODED_DATA_OUT_45
    4'b 1111, // index[90] RS_ENCODE_ENCODED_DATA_OUT_46
    4'b 1111, // index[91] RS_ENCODE_ENCODED_DATA_OUT_47
    4'b 1111, // index[92] RS_ENCODE_ENCODED_DATA_OUT_48
    4'b 1111  // index[93] RS_ENCODE_ENCODED_DATA_OUT_49
  };

endpackage


// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`

`include "prim_assert.sv"

module rs_encode_reg_top (
  input clk_i,
  input rst_ni,
  input  tlul_pkg::tl_h2d_t tl_i,
  output tlul_pkg::tl_d2h_t tl_o,
  // To HW
  output rs_encode_reg_pkg::rs_encode_reg2hw_t reg2hw, // Write
  input  rs_encode_reg_pkg::rs_encode_hw2reg_t hw2reg, // Read

  // Integrity check errors
  output logic intg_err_o,

  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import rs_encode_reg_pkg::* ;

  localparam int AW = 9;
  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;
  logic reg_busy;

  tlul_pkg::tl_h2d_t tl_reg_h2d;
  tlul_pkg::tl_d2h_t tl_reg_d2h;


  // incoming payload check
  logic intg_err;
  tlul_cmd_intg_chk u_chk (
    .tl_i(tl_i),
    .err_o(intg_err)
  );

  // also check for spurious write enables
  logic reg_we_err;
  logic [93:0] reg_we_check;
  prim_reg_we_check #(
    .OneHotWidth(94)
  ) u_prim_reg_we_check (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .oh_i  (reg_we_check),
    .en_i  (reg_we && !addrmiss),
    .err_o (reg_we_err)
  );

  logic err_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      err_q <= '0;
    end else if (intg_err || reg_we_err) begin
      err_q <= 1'b1;
    end
  end

  // integrity error output is permanent and should be used for alert generation
  // register errors are transactional
  assign intg_err_o = err_q | intg_err | reg_we_err;

  // outgoing integrity generation
  tlul_pkg::tl_d2h_t tl_o_pre;
  tlul_rsp_intg_gen #(
    .EnableRspIntgGen(1),
    .EnableDataIntgGen(1)
  ) u_rsp_intg_gen (
    .tl_i(tl_o_pre),
    .tl_o(tl_o)
  );

  assign tl_reg_h2d = tl_i;
  assign tl_o_pre   = tl_reg_d2h;

  tlul_adapter_reg #(
    .RegAw(AW),
    .RegDw(DW),
    .EnableDataIntgGen(0)
  ) u_reg_if (
    .clk_i  (clk_i),
    .rst_ni (rst_ni),

    .tl_i (tl_reg_h2d),
    .tl_o (tl_reg_d2h),

    .en_ifetch_i(prim_mubi_pkg::MuBi4False),
    .intg_error_o(),

    .we_o    (reg_we),
    .re_o    (reg_re),
    .addr_o  (reg_addr),
    .wdata_o (reg_wdata),
    .be_o    (reg_be),
    .busy_i  (reg_busy),
    .rdata_i (reg_rdata),
    .error_i (reg_error)
  );

  // cdc oversampling signals

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err | intg_err;

  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic ctrl_signals_we;
  logic ctrl_signals_encode_en_qs;
  logic ctrl_signals_encode_en_wd;
  logic ctrl_signals_clrn_qs;
  logic ctrl_signals_clrn_wd;
  logic state_signals_valid_bit_qs;
  logic state_signals_ready_bit_qs;
  logic data_in_0_we;
  logic [31:0] data_in_0_qs;
  logic [31:0] data_in_0_wd;
  logic data_in_1_we;
  logic [31:0] data_in_1_qs;
  logic [31:0] data_in_1_wd;
  logic data_in_2_we;
  logic [31:0] data_in_2_qs;
  logic [31:0] data_in_2_wd;
  logic data_in_3_we;
  logic [31:0] data_in_3_qs;
  logic [31:0] data_in_3_wd;
  logic data_in_4_we;
  logic [31:0] data_in_4_qs;
  logic [31:0] data_in_4_wd;
  logic data_in_5_we;
  logic [31:0] data_in_5_qs;
  logic [31:0] data_in_5_wd;
  logic data_in_6_we;
  logic [31:0] data_in_6_qs;
  logic [31:0] data_in_6_wd;
  logic data_in_7_we;
  logic [31:0] data_in_7_qs;
  logic [31:0] data_in_7_wd;
  logic data_in_8_we;
  logic [31:0] data_in_8_qs;
  logic [31:0] data_in_8_wd;
  logic data_in_9_we;
  logic [31:0] data_in_9_qs;
  logic [31:0] data_in_9_wd;
  logic data_in_10_we;
  logic [31:0] data_in_10_qs;
  logic [31:0] data_in_10_wd;
  logic data_in_11_we;
  logic [31:0] data_in_11_qs;
  logic [31:0] data_in_11_wd;
  logic data_in_12_we;
  logic [31:0] data_in_12_qs;
  logic [31:0] data_in_12_wd;
  logic data_in_13_we;
  logic [31:0] data_in_13_qs;
  logic [31:0] data_in_13_wd;
  logic data_in_14_we;
  logic [31:0] data_in_14_qs;
  logic [31:0] data_in_14_wd;
  logic data_in_15_we;
  logic [31:0] data_in_15_qs;
  logic [31:0] data_in_15_wd;
  logic data_in_16_we;
  logic [31:0] data_in_16_qs;
  logic [31:0] data_in_16_wd;
  logic data_in_17_we;
  logic [31:0] data_in_17_qs;
  logic [31:0] data_in_17_wd;
  logic data_in_18_we;
  logic [31:0] data_in_18_qs;
  logic [31:0] data_in_18_wd;
  logic data_in_19_we;
  logic [31:0] data_in_19_qs;
  logic [31:0] data_in_19_wd;
  logic data_in_20_we;
  logic [31:0] data_in_20_qs;
  logic [31:0] data_in_20_wd;
  logic data_in_21_we;
  logic [31:0] data_in_21_qs;
  logic [31:0] data_in_21_wd;
  logic data_in_22_we;
  logic [31:0] data_in_22_qs;
  logic [31:0] data_in_22_wd;
  logic data_in_23_we;
  logic [31:0] data_in_23_qs;
  logic [31:0] data_in_23_wd;
  logic data_in_24_we;
  logic [31:0] data_in_24_qs;
  logic [31:0] data_in_24_wd;
  logic data_in_25_we;
  logic [31:0] data_in_25_qs;
  logic [31:0] data_in_25_wd;
  logic data_in_26_we;
  logic [31:0] data_in_26_qs;
  logic [31:0] data_in_26_wd;
  logic data_in_27_we;
  logic [31:0] data_in_27_qs;
  logic [31:0] data_in_27_wd;
  logic data_in_28_we;
  logic [31:0] data_in_28_qs;
  logic [31:0] data_in_28_wd;
  logic data_in_29_we;
  logic [31:0] data_in_29_qs;
  logic [31:0] data_in_29_wd;
  logic data_in_30_we;
  logic [31:0] data_in_30_qs;
  logic [31:0] data_in_30_wd;
  logic data_in_31_we;
  logic [31:0] data_in_31_qs;
  logic [31:0] data_in_31_wd;
  logic data_in_32_we;
  logic [31:0] data_in_32_qs;
  logic [31:0] data_in_32_wd;
  logic data_in_33_we;
  logic [31:0] data_in_33_qs;
  logic [31:0] data_in_33_wd;
  logic data_in_34_we;
  logic [31:0] data_in_34_qs;
  logic [31:0] data_in_34_wd;
  logic data_in_35_we;
  logic [31:0] data_in_35_qs;
  logic [31:0] data_in_35_wd;
  logic data_in_36_we;
  logic [31:0] data_in_36_qs;
  logic [31:0] data_in_36_wd;
  logic data_in_37_we;
  logic [31:0] data_in_37_qs;
  logic [31:0] data_in_37_wd;
  logic data_in_38_we;
  logic [31:0] data_in_38_qs;
  logic [31:0] data_in_38_wd;
  logic data_in_39_we;
  logic [31:0] data_in_39_qs;
  logic [31:0] data_in_39_wd;
  logic data_in_40_we;
  logic [31:0] data_in_40_qs;
  logic [31:0] data_in_40_wd;
  logic data_in_41_we;
  logic [31:0] data_in_41_qs;
  logic [31:0] data_in_41_wd;
  logic [31:0] encoded_data_out_0_qs;
  logic [31:0] encoded_data_out_1_qs;
  logic [31:0] encoded_data_out_2_qs;
  logic [31:0] encoded_data_out_3_qs;
  logic [31:0] encoded_data_out_4_qs;
  logic [31:0] encoded_data_out_5_qs;
  logic [31:0] encoded_data_out_6_qs;
  logic [31:0] encoded_data_out_7_qs;
  logic [31:0] encoded_data_out_8_qs;
  logic [31:0] encoded_data_out_9_qs;
  logic [31:0] encoded_data_out_10_qs;
  logic [31:0] encoded_data_out_11_qs;
  logic [31:0] encoded_data_out_12_qs;
  logic [31:0] encoded_data_out_13_qs;
  logic [31:0] encoded_data_out_14_qs;
  logic [31:0] encoded_data_out_15_qs;
  logic [31:0] encoded_data_out_16_qs;
  logic [31:0] encoded_data_out_17_qs;
  logic [31:0] encoded_data_out_18_qs;
  logic [31:0] encoded_data_out_19_qs;
  logic [31:0] encoded_data_out_20_qs;
  logic [31:0] encoded_data_out_21_qs;
  logic [31:0] encoded_data_out_22_qs;
  logic [31:0] encoded_data_out_23_qs;
  logic [31:0] encoded_data_out_24_qs;
  logic [31:0] encoded_data_out_25_qs;
  logic [31:0] encoded_data_out_26_qs;
  logic [31:0] encoded_data_out_27_qs;
  logic [31:0] encoded_data_out_28_qs;
  logic [31:0] encoded_data_out_29_qs;
  logic [31:0] encoded_data_out_30_qs;
  logic [31:0] encoded_data_out_31_qs;
  logic [31:0] encoded_data_out_32_qs;
  logic [31:0] encoded_data_out_33_qs;
  logic [31:0] encoded_data_out_34_qs;
  logic [31:0] encoded_data_out_35_qs;
  logic [31:0] encoded_data_out_36_qs;
  logic [31:0] encoded_data_out_37_qs;
  logic [31:0] encoded_data_out_38_qs;
  logic [31:0] encoded_data_out_39_qs;
  logic [31:0] encoded_data_out_40_qs;
  logic [31:0] encoded_data_out_41_qs;
  logic [31:0] encoded_data_out_42_qs;
  logic [31:0] encoded_data_out_43_qs;
  logic [31:0] encoded_data_out_44_qs;
  logic [31:0] encoded_data_out_45_qs;
  logic [31:0] encoded_data_out_46_qs;
  logic [31:0] encoded_data_out_47_qs;
  logic [31:0] encoded_data_out_48_qs;
  logic [31:0] encoded_data_out_49_qs;

  // Register instances
  // R[ctrl_signals]: V(False)
  logic ctrl_signals_qe;
  logic [1:0] ctrl_signals_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_ctrl_signals0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&ctrl_signals_flds_we),
    .q_o(ctrl_signals_qe)
  );
  //   F[encode_en]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h0)
  ) u_ctrl_signals_encode_en (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_encode_en_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.encode_en.de),
    .d      (hw2reg.ctrl_signals.encode_en.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[0]),
    .q      (reg2hw.ctrl_signals.encode_en.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_encode_en_qs)
  );
  assign reg2hw.ctrl_signals.encode_en.qe = ctrl_signals_qe;

  //   F[clrn]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (1'h1)
  ) u_ctrl_signals_clrn (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (ctrl_signals_we),
    .wd     (ctrl_signals_clrn_wd),

    // from internal hardware
    .de     (hw2reg.ctrl_signals.clrn.de),
    .d      (hw2reg.ctrl_signals.clrn.d),

    // to internal hardware
    .qe     (ctrl_signals_flds_we[1]),
    .q      (reg2hw.ctrl_signals.clrn.q),
    .ds     (),

    // to register interface (read)
    .qs     (ctrl_signals_clrn_qs)
  );
  assign reg2hw.ctrl_signals.clrn.qe = ctrl_signals_qe;


  // R[state_signals]: V(False)
  //   F[valid_bit]: 0:0
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_valid_bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.valid_bit.de),
    .d      (hw2reg.state_signals.valid_bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.valid_bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_valid_bit_qs)
  );

  //   F[ready_bit]: 1:1
  prim_subreg #(
    .DW      (1),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (1'h0)
  ) u_state_signals_ready_bit (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.state_signals.ready_bit.de),
    .d      (hw2reg.state_signals.ready_bit.d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.state_signals.ready_bit.q),
    .ds     (),

    // to register interface (read)
    .qs     (state_signals_ready_bit_qs)
  );


  // Subregister 0 of Multireg data_in
  // R[data_in_0]: V(False)
  logic data_in_0_qe;
  logic [0:0] data_in_0_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in0_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_0_flds_we),
    .q_o(data_in_0_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_0_we),
    .wd     (data_in_0_wd),

    // from internal hardware
    .de     (hw2reg.data_in[0].de),
    .d      (hw2reg.data_in[0].d),

    // to internal hardware
    .qe     (data_in_0_flds_we[0]),
    .q      (reg2hw.data_in[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_0_qs)
  );
  assign reg2hw.data_in[0].qe = data_in_0_qe;


  // Subregister 1 of Multireg data_in
  // R[data_in_1]: V(False)
  logic data_in_1_qe;
  logic [0:0] data_in_1_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in1_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_1_flds_we),
    .q_o(data_in_1_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_1_we),
    .wd     (data_in_1_wd),

    // from internal hardware
    .de     (hw2reg.data_in[1].de),
    .d      (hw2reg.data_in[1].d),

    // to internal hardware
    .qe     (data_in_1_flds_we[0]),
    .q      (reg2hw.data_in[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_1_qs)
  );
  assign reg2hw.data_in[1].qe = data_in_1_qe;


  // Subregister 2 of Multireg data_in
  // R[data_in_2]: V(False)
  logic data_in_2_qe;
  logic [0:0] data_in_2_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in2_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_2_flds_we),
    .q_o(data_in_2_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_2_we),
    .wd     (data_in_2_wd),

    // from internal hardware
    .de     (hw2reg.data_in[2].de),
    .d      (hw2reg.data_in[2].d),

    // to internal hardware
    .qe     (data_in_2_flds_we[0]),
    .q      (reg2hw.data_in[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_2_qs)
  );
  assign reg2hw.data_in[2].qe = data_in_2_qe;


  // Subregister 3 of Multireg data_in
  // R[data_in_3]: V(False)
  logic data_in_3_qe;
  logic [0:0] data_in_3_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in3_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_3_flds_we),
    .q_o(data_in_3_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_3_we),
    .wd     (data_in_3_wd),

    // from internal hardware
    .de     (hw2reg.data_in[3].de),
    .d      (hw2reg.data_in[3].d),

    // to internal hardware
    .qe     (data_in_3_flds_we[0]),
    .q      (reg2hw.data_in[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_3_qs)
  );
  assign reg2hw.data_in[3].qe = data_in_3_qe;


  // Subregister 4 of Multireg data_in
  // R[data_in_4]: V(False)
  logic data_in_4_qe;
  logic [0:0] data_in_4_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in4_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_4_flds_we),
    .q_o(data_in_4_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_4_we),
    .wd     (data_in_4_wd),

    // from internal hardware
    .de     (hw2reg.data_in[4].de),
    .d      (hw2reg.data_in[4].d),

    // to internal hardware
    .qe     (data_in_4_flds_we[0]),
    .q      (reg2hw.data_in[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_4_qs)
  );
  assign reg2hw.data_in[4].qe = data_in_4_qe;


  // Subregister 5 of Multireg data_in
  // R[data_in_5]: V(False)
  logic data_in_5_qe;
  logic [0:0] data_in_5_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in5_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_5_flds_we),
    .q_o(data_in_5_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_5_we),
    .wd     (data_in_5_wd),

    // from internal hardware
    .de     (hw2reg.data_in[5].de),
    .d      (hw2reg.data_in[5].d),

    // to internal hardware
    .qe     (data_in_5_flds_we[0]),
    .q      (reg2hw.data_in[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_5_qs)
  );
  assign reg2hw.data_in[5].qe = data_in_5_qe;


  // Subregister 6 of Multireg data_in
  // R[data_in_6]: V(False)
  logic data_in_6_qe;
  logic [0:0] data_in_6_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in6_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_6_flds_we),
    .q_o(data_in_6_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_6_we),
    .wd     (data_in_6_wd),

    // from internal hardware
    .de     (hw2reg.data_in[6].de),
    .d      (hw2reg.data_in[6].d),

    // to internal hardware
    .qe     (data_in_6_flds_we[0]),
    .q      (reg2hw.data_in[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_6_qs)
  );
  assign reg2hw.data_in[6].qe = data_in_6_qe;


  // Subregister 7 of Multireg data_in
  // R[data_in_7]: V(False)
  logic data_in_7_qe;
  logic [0:0] data_in_7_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in7_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_7_flds_we),
    .q_o(data_in_7_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_7_we),
    .wd     (data_in_7_wd),

    // from internal hardware
    .de     (hw2reg.data_in[7].de),
    .d      (hw2reg.data_in[7].d),

    // to internal hardware
    .qe     (data_in_7_flds_we[0]),
    .q      (reg2hw.data_in[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_7_qs)
  );
  assign reg2hw.data_in[7].qe = data_in_7_qe;


  // Subregister 8 of Multireg data_in
  // R[data_in_8]: V(False)
  logic data_in_8_qe;
  logic [0:0] data_in_8_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in8_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_8_flds_we),
    .q_o(data_in_8_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_8 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_8_we),
    .wd     (data_in_8_wd),

    // from internal hardware
    .de     (hw2reg.data_in[8].de),
    .d      (hw2reg.data_in[8].d),

    // to internal hardware
    .qe     (data_in_8_flds_we[0]),
    .q      (reg2hw.data_in[8].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_8_qs)
  );
  assign reg2hw.data_in[8].qe = data_in_8_qe;


  // Subregister 9 of Multireg data_in
  // R[data_in_9]: V(False)
  logic data_in_9_qe;
  logic [0:0] data_in_9_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in9_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_9_flds_we),
    .q_o(data_in_9_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_9 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_9_we),
    .wd     (data_in_9_wd),

    // from internal hardware
    .de     (hw2reg.data_in[9].de),
    .d      (hw2reg.data_in[9].d),

    // to internal hardware
    .qe     (data_in_9_flds_we[0]),
    .q      (reg2hw.data_in[9].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_9_qs)
  );
  assign reg2hw.data_in[9].qe = data_in_9_qe;


  // Subregister 10 of Multireg data_in
  // R[data_in_10]: V(False)
  logic data_in_10_qe;
  logic [0:0] data_in_10_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in10_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_10_flds_we),
    .q_o(data_in_10_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_10 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_10_we),
    .wd     (data_in_10_wd),

    // from internal hardware
    .de     (hw2reg.data_in[10].de),
    .d      (hw2reg.data_in[10].d),

    // to internal hardware
    .qe     (data_in_10_flds_we[0]),
    .q      (reg2hw.data_in[10].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_10_qs)
  );
  assign reg2hw.data_in[10].qe = data_in_10_qe;


  // Subregister 11 of Multireg data_in
  // R[data_in_11]: V(False)
  logic data_in_11_qe;
  logic [0:0] data_in_11_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in11_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_11_flds_we),
    .q_o(data_in_11_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_11 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_11_we),
    .wd     (data_in_11_wd),

    // from internal hardware
    .de     (hw2reg.data_in[11].de),
    .d      (hw2reg.data_in[11].d),

    // to internal hardware
    .qe     (data_in_11_flds_we[0]),
    .q      (reg2hw.data_in[11].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_11_qs)
  );
  assign reg2hw.data_in[11].qe = data_in_11_qe;


  // Subregister 12 of Multireg data_in
  // R[data_in_12]: V(False)
  logic data_in_12_qe;
  logic [0:0] data_in_12_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in12_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_12_flds_we),
    .q_o(data_in_12_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_12 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_12_we),
    .wd     (data_in_12_wd),

    // from internal hardware
    .de     (hw2reg.data_in[12].de),
    .d      (hw2reg.data_in[12].d),

    // to internal hardware
    .qe     (data_in_12_flds_we[0]),
    .q      (reg2hw.data_in[12].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_12_qs)
  );
  assign reg2hw.data_in[12].qe = data_in_12_qe;


  // Subregister 13 of Multireg data_in
  // R[data_in_13]: V(False)
  logic data_in_13_qe;
  logic [0:0] data_in_13_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in13_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_13_flds_we),
    .q_o(data_in_13_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_13 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_13_we),
    .wd     (data_in_13_wd),

    // from internal hardware
    .de     (hw2reg.data_in[13].de),
    .d      (hw2reg.data_in[13].d),

    // to internal hardware
    .qe     (data_in_13_flds_we[0]),
    .q      (reg2hw.data_in[13].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_13_qs)
  );
  assign reg2hw.data_in[13].qe = data_in_13_qe;


  // Subregister 14 of Multireg data_in
  // R[data_in_14]: V(False)
  logic data_in_14_qe;
  logic [0:0] data_in_14_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in14_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_14_flds_we),
    .q_o(data_in_14_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_14 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_14_we),
    .wd     (data_in_14_wd),

    // from internal hardware
    .de     (hw2reg.data_in[14].de),
    .d      (hw2reg.data_in[14].d),

    // to internal hardware
    .qe     (data_in_14_flds_we[0]),
    .q      (reg2hw.data_in[14].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_14_qs)
  );
  assign reg2hw.data_in[14].qe = data_in_14_qe;


  // Subregister 15 of Multireg data_in
  // R[data_in_15]: V(False)
  logic data_in_15_qe;
  logic [0:0] data_in_15_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in15_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_15_flds_we),
    .q_o(data_in_15_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_15 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_15_we),
    .wd     (data_in_15_wd),

    // from internal hardware
    .de     (hw2reg.data_in[15].de),
    .d      (hw2reg.data_in[15].d),

    // to internal hardware
    .qe     (data_in_15_flds_we[0]),
    .q      (reg2hw.data_in[15].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_15_qs)
  );
  assign reg2hw.data_in[15].qe = data_in_15_qe;


  // Subregister 16 of Multireg data_in
  // R[data_in_16]: V(False)
  logic data_in_16_qe;
  logic [0:0] data_in_16_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in16_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_16_flds_we),
    .q_o(data_in_16_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_16 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_16_we),
    .wd     (data_in_16_wd),

    // from internal hardware
    .de     (hw2reg.data_in[16].de),
    .d      (hw2reg.data_in[16].d),

    // to internal hardware
    .qe     (data_in_16_flds_we[0]),
    .q      (reg2hw.data_in[16].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_16_qs)
  );
  assign reg2hw.data_in[16].qe = data_in_16_qe;


  // Subregister 17 of Multireg data_in
  // R[data_in_17]: V(False)
  logic data_in_17_qe;
  logic [0:0] data_in_17_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in17_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_17_flds_we),
    .q_o(data_in_17_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_17 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_17_we),
    .wd     (data_in_17_wd),

    // from internal hardware
    .de     (hw2reg.data_in[17].de),
    .d      (hw2reg.data_in[17].d),

    // to internal hardware
    .qe     (data_in_17_flds_we[0]),
    .q      (reg2hw.data_in[17].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_17_qs)
  );
  assign reg2hw.data_in[17].qe = data_in_17_qe;


  // Subregister 18 of Multireg data_in
  // R[data_in_18]: V(False)
  logic data_in_18_qe;
  logic [0:0] data_in_18_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in18_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_18_flds_we),
    .q_o(data_in_18_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_18 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_18_we),
    .wd     (data_in_18_wd),

    // from internal hardware
    .de     (hw2reg.data_in[18].de),
    .d      (hw2reg.data_in[18].d),

    // to internal hardware
    .qe     (data_in_18_flds_we[0]),
    .q      (reg2hw.data_in[18].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_18_qs)
  );
  assign reg2hw.data_in[18].qe = data_in_18_qe;


  // Subregister 19 of Multireg data_in
  // R[data_in_19]: V(False)
  logic data_in_19_qe;
  logic [0:0] data_in_19_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in19_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_19_flds_we),
    .q_o(data_in_19_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_19 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_19_we),
    .wd     (data_in_19_wd),

    // from internal hardware
    .de     (hw2reg.data_in[19].de),
    .d      (hw2reg.data_in[19].d),

    // to internal hardware
    .qe     (data_in_19_flds_we[0]),
    .q      (reg2hw.data_in[19].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_19_qs)
  );
  assign reg2hw.data_in[19].qe = data_in_19_qe;


  // Subregister 20 of Multireg data_in
  // R[data_in_20]: V(False)
  logic data_in_20_qe;
  logic [0:0] data_in_20_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in20_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_20_flds_we),
    .q_o(data_in_20_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_20 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_20_we),
    .wd     (data_in_20_wd),

    // from internal hardware
    .de     (hw2reg.data_in[20].de),
    .d      (hw2reg.data_in[20].d),

    // to internal hardware
    .qe     (data_in_20_flds_we[0]),
    .q      (reg2hw.data_in[20].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_20_qs)
  );
  assign reg2hw.data_in[20].qe = data_in_20_qe;


  // Subregister 21 of Multireg data_in
  // R[data_in_21]: V(False)
  logic data_in_21_qe;
  logic [0:0] data_in_21_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in21_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_21_flds_we),
    .q_o(data_in_21_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_21 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_21_we),
    .wd     (data_in_21_wd),

    // from internal hardware
    .de     (hw2reg.data_in[21].de),
    .d      (hw2reg.data_in[21].d),

    // to internal hardware
    .qe     (data_in_21_flds_we[0]),
    .q      (reg2hw.data_in[21].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_21_qs)
  );
  assign reg2hw.data_in[21].qe = data_in_21_qe;


  // Subregister 22 of Multireg data_in
  // R[data_in_22]: V(False)
  logic data_in_22_qe;
  logic [0:0] data_in_22_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in22_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_22_flds_we),
    .q_o(data_in_22_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_22 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_22_we),
    .wd     (data_in_22_wd),

    // from internal hardware
    .de     (hw2reg.data_in[22].de),
    .d      (hw2reg.data_in[22].d),

    // to internal hardware
    .qe     (data_in_22_flds_we[0]),
    .q      (reg2hw.data_in[22].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_22_qs)
  );
  assign reg2hw.data_in[22].qe = data_in_22_qe;


  // Subregister 23 of Multireg data_in
  // R[data_in_23]: V(False)
  logic data_in_23_qe;
  logic [0:0] data_in_23_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in23_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_23_flds_we),
    .q_o(data_in_23_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_23 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_23_we),
    .wd     (data_in_23_wd),

    // from internal hardware
    .de     (hw2reg.data_in[23].de),
    .d      (hw2reg.data_in[23].d),

    // to internal hardware
    .qe     (data_in_23_flds_we[0]),
    .q      (reg2hw.data_in[23].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_23_qs)
  );
  assign reg2hw.data_in[23].qe = data_in_23_qe;


  // Subregister 24 of Multireg data_in
  // R[data_in_24]: V(False)
  logic data_in_24_qe;
  logic [0:0] data_in_24_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in24_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_24_flds_we),
    .q_o(data_in_24_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_24 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_24_we),
    .wd     (data_in_24_wd),

    // from internal hardware
    .de     (hw2reg.data_in[24].de),
    .d      (hw2reg.data_in[24].d),

    // to internal hardware
    .qe     (data_in_24_flds_we[0]),
    .q      (reg2hw.data_in[24].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_24_qs)
  );
  assign reg2hw.data_in[24].qe = data_in_24_qe;


  // Subregister 25 of Multireg data_in
  // R[data_in_25]: V(False)
  logic data_in_25_qe;
  logic [0:0] data_in_25_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in25_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_25_flds_we),
    .q_o(data_in_25_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_25 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_25_we),
    .wd     (data_in_25_wd),

    // from internal hardware
    .de     (hw2reg.data_in[25].de),
    .d      (hw2reg.data_in[25].d),

    // to internal hardware
    .qe     (data_in_25_flds_we[0]),
    .q      (reg2hw.data_in[25].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_25_qs)
  );
  assign reg2hw.data_in[25].qe = data_in_25_qe;


  // Subregister 26 of Multireg data_in
  // R[data_in_26]: V(False)
  logic data_in_26_qe;
  logic [0:0] data_in_26_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in26_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_26_flds_we),
    .q_o(data_in_26_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_26 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_26_we),
    .wd     (data_in_26_wd),

    // from internal hardware
    .de     (hw2reg.data_in[26].de),
    .d      (hw2reg.data_in[26].d),

    // to internal hardware
    .qe     (data_in_26_flds_we[0]),
    .q      (reg2hw.data_in[26].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_26_qs)
  );
  assign reg2hw.data_in[26].qe = data_in_26_qe;


  // Subregister 27 of Multireg data_in
  // R[data_in_27]: V(False)
  logic data_in_27_qe;
  logic [0:0] data_in_27_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in27_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_27_flds_we),
    .q_o(data_in_27_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_27 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_27_we),
    .wd     (data_in_27_wd),

    // from internal hardware
    .de     (hw2reg.data_in[27].de),
    .d      (hw2reg.data_in[27].d),

    // to internal hardware
    .qe     (data_in_27_flds_we[0]),
    .q      (reg2hw.data_in[27].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_27_qs)
  );
  assign reg2hw.data_in[27].qe = data_in_27_qe;


  // Subregister 28 of Multireg data_in
  // R[data_in_28]: V(False)
  logic data_in_28_qe;
  logic [0:0] data_in_28_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in28_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_28_flds_we),
    .q_o(data_in_28_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_28 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_28_we),
    .wd     (data_in_28_wd),

    // from internal hardware
    .de     (hw2reg.data_in[28].de),
    .d      (hw2reg.data_in[28].d),

    // to internal hardware
    .qe     (data_in_28_flds_we[0]),
    .q      (reg2hw.data_in[28].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_28_qs)
  );
  assign reg2hw.data_in[28].qe = data_in_28_qe;


  // Subregister 29 of Multireg data_in
  // R[data_in_29]: V(False)
  logic data_in_29_qe;
  logic [0:0] data_in_29_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in29_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_29_flds_we),
    .q_o(data_in_29_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_29 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_29_we),
    .wd     (data_in_29_wd),

    // from internal hardware
    .de     (hw2reg.data_in[29].de),
    .d      (hw2reg.data_in[29].d),

    // to internal hardware
    .qe     (data_in_29_flds_we[0]),
    .q      (reg2hw.data_in[29].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_29_qs)
  );
  assign reg2hw.data_in[29].qe = data_in_29_qe;


  // Subregister 30 of Multireg data_in
  // R[data_in_30]: V(False)
  logic data_in_30_qe;
  logic [0:0] data_in_30_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in30_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_30_flds_we),
    .q_o(data_in_30_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_30 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_30_we),
    .wd     (data_in_30_wd),

    // from internal hardware
    .de     (hw2reg.data_in[30].de),
    .d      (hw2reg.data_in[30].d),

    // to internal hardware
    .qe     (data_in_30_flds_we[0]),
    .q      (reg2hw.data_in[30].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_30_qs)
  );
  assign reg2hw.data_in[30].qe = data_in_30_qe;


  // Subregister 31 of Multireg data_in
  // R[data_in_31]: V(False)
  logic data_in_31_qe;
  logic [0:0] data_in_31_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in31_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_31_flds_we),
    .q_o(data_in_31_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_31 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_31_we),
    .wd     (data_in_31_wd),

    // from internal hardware
    .de     (hw2reg.data_in[31].de),
    .d      (hw2reg.data_in[31].d),

    // to internal hardware
    .qe     (data_in_31_flds_we[0]),
    .q      (reg2hw.data_in[31].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_31_qs)
  );
  assign reg2hw.data_in[31].qe = data_in_31_qe;


  // Subregister 32 of Multireg data_in
  // R[data_in_32]: V(False)
  logic data_in_32_qe;
  logic [0:0] data_in_32_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in32_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_32_flds_we),
    .q_o(data_in_32_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_32 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_32_we),
    .wd     (data_in_32_wd),

    // from internal hardware
    .de     (hw2reg.data_in[32].de),
    .d      (hw2reg.data_in[32].d),

    // to internal hardware
    .qe     (data_in_32_flds_we[0]),
    .q      (reg2hw.data_in[32].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_32_qs)
  );
  assign reg2hw.data_in[32].qe = data_in_32_qe;


  // Subregister 33 of Multireg data_in
  // R[data_in_33]: V(False)
  logic data_in_33_qe;
  logic [0:0] data_in_33_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in33_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_33_flds_we),
    .q_o(data_in_33_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_33 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_33_we),
    .wd     (data_in_33_wd),

    // from internal hardware
    .de     (hw2reg.data_in[33].de),
    .d      (hw2reg.data_in[33].d),

    // to internal hardware
    .qe     (data_in_33_flds_we[0]),
    .q      (reg2hw.data_in[33].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_33_qs)
  );
  assign reg2hw.data_in[33].qe = data_in_33_qe;


  // Subregister 34 of Multireg data_in
  // R[data_in_34]: V(False)
  logic data_in_34_qe;
  logic [0:0] data_in_34_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in34_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_34_flds_we),
    .q_o(data_in_34_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_34 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_34_we),
    .wd     (data_in_34_wd),

    // from internal hardware
    .de     (hw2reg.data_in[34].de),
    .d      (hw2reg.data_in[34].d),

    // to internal hardware
    .qe     (data_in_34_flds_we[0]),
    .q      (reg2hw.data_in[34].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_34_qs)
  );
  assign reg2hw.data_in[34].qe = data_in_34_qe;


  // Subregister 35 of Multireg data_in
  // R[data_in_35]: V(False)
  logic data_in_35_qe;
  logic [0:0] data_in_35_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in35_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_35_flds_we),
    .q_o(data_in_35_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_35 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_35_we),
    .wd     (data_in_35_wd),

    // from internal hardware
    .de     (hw2reg.data_in[35].de),
    .d      (hw2reg.data_in[35].d),

    // to internal hardware
    .qe     (data_in_35_flds_we[0]),
    .q      (reg2hw.data_in[35].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_35_qs)
  );
  assign reg2hw.data_in[35].qe = data_in_35_qe;


  // Subregister 36 of Multireg data_in
  // R[data_in_36]: V(False)
  logic data_in_36_qe;
  logic [0:0] data_in_36_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in36_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_36_flds_we),
    .q_o(data_in_36_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_36 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_36_we),
    .wd     (data_in_36_wd),

    // from internal hardware
    .de     (hw2reg.data_in[36].de),
    .d      (hw2reg.data_in[36].d),

    // to internal hardware
    .qe     (data_in_36_flds_we[0]),
    .q      (reg2hw.data_in[36].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_36_qs)
  );
  assign reg2hw.data_in[36].qe = data_in_36_qe;


  // Subregister 37 of Multireg data_in
  // R[data_in_37]: V(False)
  logic data_in_37_qe;
  logic [0:0] data_in_37_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in37_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_37_flds_we),
    .q_o(data_in_37_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_37 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_37_we),
    .wd     (data_in_37_wd),

    // from internal hardware
    .de     (hw2reg.data_in[37].de),
    .d      (hw2reg.data_in[37].d),

    // to internal hardware
    .qe     (data_in_37_flds_we[0]),
    .q      (reg2hw.data_in[37].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_37_qs)
  );
  assign reg2hw.data_in[37].qe = data_in_37_qe;


  // Subregister 38 of Multireg data_in
  // R[data_in_38]: V(False)
  logic data_in_38_qe;
  logic [0:0] data_in_38_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in38_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_38_flds_we),
    .q_o(data_in_38_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_38 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_38_we),
    .wd     (data_in_38_wd),

    // from internal hardware
    .de     (hw2reg.data_in[38].de),
    .d      (hw2reg.data_in[38].d),

    // to internal hardware
    .qe     (data_in_38_flds_we[0]),
    .q      (reg2hw.data_in[38].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_38_qs)
  );
  assign reg2hw.data_in[38].qe = data_in_38_qe;


  // Subregister 39 of Multireg data_in
  // R[data_in_39]: V(False)
  logic data_in_39_qe;
  logic [0:0] data_in_39_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in39_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_39_flds_we),
    .q_o(data_in_39_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_39 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_39_we),
    .wd     (data_in_39_wd),

    // from internal hardware
    .de     (hw2reg.data_in[39].de),
    .d      (hw2reg.data_in[39].d),

    // to internal hardware
    .qe     (data_in_39_flds_we[0]),
    .q      (reg2hw.data_in[39].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_39_qs)
  );
  assign reg2hw.data_in[39].qe = data_in_39_qe;


  // Subregister 40 of Multireg data_in
  // R[data_in_40]: V(False)
  logic data_in_40_qe;
  logic [0:0] data_in_40_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in40_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_40_flds_we),
    .q_o(data_in_40_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_40 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_40_we),
    .wd     (data_in_40_wd),

    // from internal hardware
    .de     (hw2reg.data_in[40].de),
    .d      (hw2reg.data_in[40].d),

    // to internal hardware
    .qe     (data_in_40_flds_we[0]),
    .q      (reg2hw.data_in[40].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_40_qs)
  );
  assign reg2hw.data_in[40].qe = data_in_40_qe;


  // Subregister 41 of Multireg data_in
  // R[data_in_41]: V(False)
  logic data_in_41_qe;
  logic [0:0] data_in_41_flds_we;
  prim_flop #(
    .Width(1),
    .ResetValue(0)
  ) u_data_in41_qe (
    .clk_i(clk_i),
    .rst_ni(rst_ni),
    .d_i(&data_in_41_flds_we),
    .q_o(data_in_41_qe)
  );
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRW),
    .RESVAL  (32'h0)
  ) u_data_in_41 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (data_in_41_we),
    .wd     (data_in_41_wd),

    // from internal hardware
    .de     (hw2reg.data_in[41].de),
    .d      (hw2reg.data_in[41].d),

    // to internal hardware
    .qe     (data_in_41_flds_we[0]),
    .q      (reg2hw.data_in[41].q),
    .ds     (),

    // to register interface (read)
    .qs     (data_in_41_qs)
  );
  assign reg2hw.data_in[41].qe = data_in_41_qe;


  // Subregister 0 of Multireg encoded_data_out
  // R[encoded_data_out_0]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_0 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[0].de),
    .d      (hw2reg.encoded_data_out[0].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[0].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_0_qs)
  );


  // Subregister 1 of Multireg encoded_data_out
  // R[encoded_data_out_1]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_1 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[1].de),
    .d      (hw2reg.encoded_data_out[1].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[1].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_1_qs)
  );


  // Subregister 2 of Multireg encoded_data_out
  // R[encoded_data_out_2]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_2 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[2].de),
    .d      (hw2reg.encoded_data_out[2].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[2].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_2_qs)
  );


  // Subregister 3 of Multireg encoded_data_out
  // R[encoded_data_out_3]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_3 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[3].de),
    .d      (hw2reg.encoded_data_out[3].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[3].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_3_qs)
  );


  // Subregister 4 of Multireg encoded_data_out
  // R[encoded_data_out_4]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_4 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[4].de),
    .d      (hw2reg.encoded_data_out[4].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[4].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_4_qs)
  );


  // Subregister 5 of Multireg encoded_data_out
  // R[encoded_data_out_5]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_5 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[5].de),
    .d      (hw2reg.encoded_data_out[5].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[5].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_5_qs)
  );


  // Subregister 6 of Multireg encoded_data_out
  // R[encoded_data_out_6]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_6 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[6].de),
    .d      (hw2reg.encoded_data_out[6].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[6].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_6_qs)
  );


  // Subregister 7 of Multireg encoded_data_out
  // R[encoded_data_out_7]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_7 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[7].de),
    .d      (hw2reg.encoded_data_out[7].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[7].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_7_qs)
  );


  // Subregister 8 of Multireg encoded_data_out
  // R[encoded_data_out_8]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_8 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[8].de),
    .d      (hw2reg.encoded_data_out[8].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[8].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_8_qs)
  );


  // Subregister 9 of Multireg encoded_data_out
  // R[encoded_data_out_9]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_9 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[9].de),
    .d      (hw2reg.encoded_data_out[9].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[9].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_9_qs)
  );


  // Subregister 10 of Multireg encoded_data_out
  // R[encoded_data_out_10]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_10 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[10].de),
    .d      (hw2reg.encoded_data_out[10].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[10].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_10_qs)
  );


  // Subregister 11 of Multireg encoded_data_out
  // R[encoded_data_out_11]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_11 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[11].de),
    .d      (hw2reg.encoded_data_out[11].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[11].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_11_qs)
  );


  // Subregister 12 of Multireg encoded_data_out
  // R[encoded_data_out_12]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_12 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[12].de),
    .d      (hw2reg.encoded_data_out[12].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[12].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_12_qs)
  );


  // Subregister 13 of Multireg encoded_data_out
  // R[encoded_data_out_13]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_13 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[13].de),
    .d      (hw2reg.encoded_data_out[13].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[13].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_13_qs)
  );


  // Subregister 14 of Multireg encoded_data_out
  // R[encoded_data_out_14]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_14 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[14].de),
    .d      (hw2reg.encoded_data_out[14].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[14].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_14_qs)
  );


  // Subregister 15 of Multireg encoded_data_out
  // R[encoded_data_out_15]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_15 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[15].de),
    .d      (hw2reg.encoded_data_out[15].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[15].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_15_qs)
  );


  // Subregister 16 of Multireg encoded_data_out
  // R[encoded_data_out_16]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_16 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[16].de),
    .d      (hw2reg.encoded_data_out[16].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[16].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_16_qs)
  );


  // Subregister 17 of Multireg encoded_data_out
  // R[encoded_data_out_17]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_17 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[17].de),
    .d      (hw2reg.encoded_data_out[17].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[17].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_17_qs)
  );


  // Subregister 18 of Multireg encoded_data_out
  // R[encoded_data_out_18]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_18 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[18].de),
    .d      (hw2reg.encoded_data_out[18].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[18].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_18_qs)
  );


  // Subregister 19 of Multireg encoded_data_out
  // R[encoded_data_out_19]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_19 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[19].de),
    .d      (hw2reg.encoded_data_out[19].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[19].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_19_qs)
  );


  // Subregister 20 of Multireg encoded_data_out
  // R[encoded_data_out_20]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_20 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[20].de),
    .d      (hw2reg.encoded_data_out[20].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[20].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_20_qs)
  );


  // Subregister 21 of Multireg encoded_data_out
  // R[encoded_data_out_21]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_21 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[21].de),
    .d      (hw2reg.encoded_data_out[21].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[21].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_21_qs)
  );


  // Subregister 22 of Multireg encoded_data_out
  // R[encoded_data_out_22]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_22 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[22].de),
    .d      (hw2reg.encoded_data_out[22].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[22].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_22_qs)
  );


  // Subregister 23 of Multireg encoded_data_out
  // R[encoded_data_out_23]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_23 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[23].de),
    .d      (hw2reg.encoded_data_out[23].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[23].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_23_qs)
  );


  // Subregister 24 of Multireg encoded_data_out
  // R[encoded_data_out_24]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_24 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[24].de),
    .d      (hw2reg.encoded_data_out[24].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[24].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_24_qs)
  );


  // Subregister 25 of Multireg encoded_data_out
  // R[encoded_data_out_25]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_25 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[25].de),
    .d      (hw2reg.encoded_data_out[25].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[25].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_25_qs)
  );


  // Subregister 26 of Multireg encoded_data_out
  // R[encoded_data_out_26]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_26 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[26].de),
    .d      (hw2reg.encoded_data_out[26].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[26].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_26_qs)
  );


  // Subregister 27 of Multireg encoded_data_out
  // R[encoded_data_out_27]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_27 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[27].de),
    .d      (hw2reg.encoded_data_out[27].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[27].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_27_qs)
  );


  // Subregister 28 of Multireg encoded_data_out
  // R[encoded_data_out_28]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_28 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[28].de),
    .d      (hw2reg.encoded_data_out[28].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[28].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_28_qs)
  );


  // Subregister 29 of Multireg encoded_data_out
  // R[encoded_data_out_29]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_29 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[29].de),
    .d      (hw2reg.encoded_data_out[29].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[29].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_29_qs)
  );


  // Subregister 30 of Multireg encoded_data_out
  // R[encoded_data_out_30]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_30 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[30].de),
    .d      (hw2reg.encoded_data_out[30].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[30].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_30_qs)
  );


  // Subregister 31 of Multireg encoded_data_out
  // R[encoded_data_out_31]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_31 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[31].de),
    .d      (hw2reg.encoded_data_out[31].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[31].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_31_qs)
  );


  // Subregister 32 of Multireg encoded_data_out
  // R[encoded_data_out_32]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_32 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[32].de),
    .d      (hw2reg.encoded_data_out[32].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[32].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_32_qs)
  );


  // Subregister 33 of Multireg encoded_data_out
  // R[encoded_data_out_33]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_33 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[33].de),
    .d      (hw2reg.encoded_data_out[33].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[33].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_33_qs)
  );


  // Subregister 34 of Multireg encoded_data_out
  // R[encoded_data_out_34]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_34 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[34].de),
    .d      (hw2reg.encoded_data_out[34].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[34].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_34_qs)
  );


  // Subregister 35 of Multireg encoded_data_out
  // R[encoded_data_out_35]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_35 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[35].de),
    .d      (hw2reg.encoded_data_out[35].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[35].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_35_qs)
  );


  // Subregister 36 of Multireg encoded_data_out
  // R[encoded_data_out_36]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_36 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[36].de),
    .d      (hw2reg.encoded_data_out[36].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[36].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_36_qs)
  );


  // Subregister 37 of Multireg encoded_data_out
  // R[encoded_data_out_37]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_37 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[37].de),
    .d      (hw2reg.encoded_data_out[37].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[37].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_37_qs)
  );


  // Subregister 38 of Multireg encoded_data_out
  // R[encoded_data_out_38]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_38 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[38].de),
    .d      (hw2reg.encoded_data_out[38].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[38].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_38_qs)
  );


  // Subregister 39 of Multireg encoded_data_out
  // R[encoded_data_out_39]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_39 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[39].de),
    .d      (hw2reg.encoded_data_out[39].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[39].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_39_qs)
  );


  // Subregister 40 of Multireg encoded_data_out
  // R[encoded_data_out_40]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_40 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[40].de),
    .d      (hw2reg.encoded_data_out[40].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[40].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_40_qs)
  );


  // Subregister 41 of Multireg encoded_data_out
  // R[encoded_data_out_41]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_41 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[41].de),
    .d      (hw2reg.encoded_data_out[41].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[41].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_41_qs)
  );


  // Subregister 42 of Multireg encoded_data_out
  // R[encoded_data_out_42]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_42 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[42].de),
    .d      (hw2reg.encoded_data_out[42].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[42].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_42_qs)
  );


  // Subregister 43 of Multireg encoded_data_out
  // R[encoded_data_out_43]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_43 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[43].de),
    .d      (hw2reg.encoded_data_out[43].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[43].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_43_qs)
  );


  // Subregister 44 of Multireg encoded_data_out
  // R[encoded_data_out_44]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_44 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[44].de),
    .d      (hw2reg.encoded_data_out[44].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[44].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_44_qs)
  );


  // Subregister 45 of Multireg encoded_data_out
  // R[encoded_data_out_45]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_45 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[45].de),
    .d      (hw2reg.encoded_data_out[45].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[45].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_45_qs)
  );


  // Subregister 46 of Multireg encoded_data_out
  // R[encoded_data_out_46]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_46 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[46].de),
    .d      (hw2reg.encoded_data_out[46].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[46].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_46_qs)
  );


  // Subregister 47 of Multireg encoded_data_out
  // R[encoded_data_out_47]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_47 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[47].de),
    .d      (hw2reg.encoded_data_out[47].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[47].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_47_qs)
  );


  // Subregister 48 of Multireg encoded_data_out
  // R[encoded_data_out_48]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_48 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[48].de),
    .d      (hw2reg.encoded_data_out[48].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[48].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_48_qs)
  );


  // Subregister 49 of Multireg encoded_data_out
  // R[encoded_data_out_49]: V(False)
  prim_subreg #(
    .DW      (32),
    .SwAccess(prim_subreg_pkg::SwAccessRO),
    .RESVAL  (32'h0)
  ) u_encoded_data_out_49 (
    .clk_i   (clk_i),
    .rst_ni  (rst_ni),

    // from register interface
    .we     (1'b0),
    .wd     ('0),

    // from internal hardware
    .de     (hw2reg.encoded_data_out[49].de),
    .d      (hw2reg.encoded_data_out[49].d),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.encoded_data_out[49].q),
    .ds     (),

    // to register interface (read)
    .qs     (encoded_data_out_49_qs)
  );



  logic [93:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == RS_ENCODE_CTRL_SIGNALS_OFFSET);
    addr_hit[ 1] = (reg_addr == RS_ENCODE_STATE_SIGNALS_OFFSET);
    addr_hit[ 2] = (reg_addr == RS_ENCODE_DATA_IN_0_OFFSET);
    addr_hit[ 3] = (reg_addr == RS_ENCODE_DATA_IN_1_OFFSET);
    addr_hit[ 4] = (reg_addr == RS_ENCODE_DATA_IN_2_OFFSET);
    addr_hit[ 5] = (reg_addr == RS_ENCODE_DATA_IN_3_OFFSET);
    addr_hit[ 6] = (reg_addr == RS_ENCODE_DATA_IN_4_OFFSET);
    addr_hit[ 7] = (reg_addr == RS_ENCODE_DATA_IN_5_OFFSET);
    addr_hit[ 8] = (reg_addr == RS_ENCODE_DATA_IN_6_OFFSET);
    addr_hit[ 9] = (reg_addr == RS_ENCODE_DATA_IN_7_OFFSET);
    addr_hit[10] = (reg_addr == RS_ENCODE_DATA_IN_8_OFFSET);
    addr_hit[11] = (reg_addr == RS_ENCODE_DATA_IN_9_OFFSET);
    addr_hit[12] = (reg_addr == RS_ENCODE_DATA_IN_10_OFFSET);
    addr_hit[13] = (reg_addr == RS_ENCODE_DATA_IN_11_OFFSET);
    addr_hit[14] = (reg_addr == RS_ENCODE_DATA_IN_12_OFFSET);
    addr_hit[15] = (reg_addr == RS_ENCODE_DATA_IN_13_OFFSET);
    addr_hit[16] = (reg_addr == RS_ENCODE_DATA_IN_14_OFFSET);
    addr_hit[17] = (reg_addr == RS_ENCODE_DATA_IN_15_OFFSET);
    addr_hit[18] = (reg_addr == RS_ENCODE_DATA_IN_16_OFFSET);
    addr_hit[19] = (reg_addr == RS_ENCODE_DATA_IN_17_OFFSET);
    addr_hit[20] = (reg_addr == RS_ENCODE_DATA_IN_18_OFFSET);
    addr_hit[21] = (reg_addr == RS_ENCODE_DATA_IN_19_OFFSET);
    addr_hit[22] = (reg_addr == RS_ENCODE_DATA_IN_20_OFFSET);
    addr_hit[23] = (reg_addr == RS_ENCODE_DATA_IN_21_OFFSET);
    addr_hit[24] = (reg_addr == RS_ENCODE_DATA_IN_22_OFFSET);
    addr_hit[25] = (reg_addr == RS_ENCODE_DATA_IN_23_OFFSET);
    addr_hit[26] = (reg_addr == RS_ENCODE_DATA_IN_24_OFFSET);
    addr_hit[27] = (reg_addr == RS_ENCODE_DATA_IN_25_OFFSET);
    addr_hit[28] = (reg_addr == RS_ENCODE_DATA_IN_26_OFFSET);
    addr_hit[29] = (reg_addr == RS_ENCODE_DATA_IN_27_OFFSET);
    addr_hit[30] = (reg_addr == RS_ENCODE_DATA_IN_28_OFFSET);
    addr_hit[31] = (reg_addr == RS_ENCODE_DATA_IN_29_OFFSET);
    addr_hit[32] = (reg_addr == RS_ENCODE_DATA_IN_30_OFFSET);
    addr_hit[33] = (reg_addr == RS_ENCODE_DATA_IN_31_OFFSET);
    addr_hit[34] = (reg_addr == RS_ENCODE_DATA_IN_32_OFFSET);
    addr_hit[35] = (reg_addr == RS_ENCODE_DATA_IN_33_OFFSET);
    addr_hit[36] = (reg_addr == RS_ENCODE_DATA_IN_34_OFFSET);
    addr_hit[37] = (reg_addr == RS_ENCODE_DATA_IN_35_OFFSET);
    addr_hit[38] = (reg_addr == RS_ENCODE_DATA_IN_36_OFFSET);
    addr_hit[39] = (reg_addr == RS_ENCODE_DATA_IN_37_OFFSET);
    addr_hit[40] = (reg_addr == RS_ENCODE_DATA_IN_38_OFFSET);
    addr_hit[41] = (reg_addr == RS_ENCODE_DATA_IN_39_OFFSET);
    addr_hit[42] = (reg_addr == RS_ENCODE_DATA_IN_40_OFFSET);
    addr_hit[43] = (reg_addr == RS_ENCODE_DATA_IN_41_OFFSET);
    addr_hit[44] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_0_OFFSET);
    addr_hit[45] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_1_OFFSET);
    addr_hit[46] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_2_OFFSET);
    addr_hit[47] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_3_OFFSET);
    addr_hit[48] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_4_OFFSET);
    addr_hit[49] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_5_OFFSET);
    addr_hit[50] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_6_OFFSET);
    addr_hit[51] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_7_OFFSET);
    addr_hit[52] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_8_OFFSET);
    addr_hit[53] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_9_OFFSET);
    addr_hit[54] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_10_OFFSET);
    addr_hit[55] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_11_OFFSET);
    addr_hit[56] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_12_OFFSET);
    addr_hit[57] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_13_OFFSET);
    addr_hit[58] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_14_OFFSET);
    addr_hit[59] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_15_OFFSET);
    addr_hit[60] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_16_OFFSET);
    addr_hit[61] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_17_OFFSET);
    addr_hit[62] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_18_OFFSET);
    addr_hit[63] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_19_OFFSET);
    addr_hit[64] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_20_OFFSET);
    addr_hit[65] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_21_OFFSET);
    addr_hit[66] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_22_OFFSET);
    addr_hit[67] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_23_OFFSET);
    addr_hit[68] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_24_OFFSET);
    addr_hit[69] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_25_OFFSET);
    addr_hit[70] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_26_OFFSET);
    addr_hit[71] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_27_OFFSET);
    addr_hit[72] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_28_OFFSET);
    addr_hit[73] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_29_OFFSET);
    addr_hit[74] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_30_OFFSET);
    addr_hit[75] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_31_OFFSET);
    addr_hit[76] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_32_OFFSET);
    addr_hit[77] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_33_OFFSET);
    addr_hit[78] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_34_OFFSET);
    addr_hit[79] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_35_OFFSET);
    addr_hit[80] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_36_OFFSET);
    addr_hit[81] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_37_OFFSET);
    addr_hit[82] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_38_OFFSET);
    addr_hit[83] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_39_OFFSET);
    addr_hit[84] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_40_OFFSET);
    addr_hit[85] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_41_OFFSET);
    addr_hit[86] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_42_OFFSET);
    addr_hit[87] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_43_OFFSET);
    addr_hit[88] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_44_OFFSET);
    addr_hit[89] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_45_OFFSET);
    addr_hit[90] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_46_OFFSET);
    addr_hit[91] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_47_OFFSET);
    addr_hit[92] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_48_OFFSET);
    addr_hit[93] = (reg_addr == RS_ENCODE_ENCODED_DATA_OUT_49_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(RS_ENCODE_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(RS_ENCODE_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(RS_ENCODE_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(RS_ENCODE_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(RS_ENCODE_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(RS_ENCODE_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(RS_ENCODE_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(RS_ENCODE_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(RS_ENCODE_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(RS_ENCODE_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(RS_ENCODE_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(RS_ENCODE_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(RS_ENCODE_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(RS_ENCODE_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(RS_ENCODE_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(RS_ENCODE_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(RS_ENCODE_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(RS_ENCODE_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(RS_ENCODE_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(RS_ENCODE_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(RS_ENCODE_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(RS_ENCODE_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(RS_ENCODE_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(RS_ENCODE_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(RS_ENCODE_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(RS_ENCODE_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(RS_ENCODE_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(RS_ENCODE_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(RS_ENCODE_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(RS_ENCODE_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(RS_ENCODE_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(RS_ENCODE_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(RS_ENCODE_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(RS_ENCODE_PERMIT[33] & ~reg_be))) |
               (addr_hit[34] & (|(RS_ENCODE_PERMIT[34] & ~reg_be))) |
               (addr_hit[35] & (|(RS_ENCODE_PERMIT[35] & ~reg_be))) |
               (addr_hit[36] & (|(RS_ENCODE_PERMIT[36] & ~reg_be))) |
               (addr_hit[37] & (|(RS_ENCODE_PERMIT[37] & ~reg_be))) |
               (addr_hit[38] & (|(RS_ENCODE_PERMIT[38] & ~reg_be))) |
               (addr_hit[39] & (|(RS_ENCODE_PERMIT[39] & ~reg_be))) |
               (addr_hit[40] & (|(RS_ENCODE_PERMIT[40] & ~reg_be))) |
               (addr_hit[41] & (|(RS_ENCODE_PERMIT[41] & ~reg_be))) |
               (addr_hit[42] & (|(RS_ENCODE_PERMIT[42] & ~reg_be))) |
               (addr_hit[43] & (|(RS_ENCODE_PERMIT[43] & ~reg_be))) |
               (addr_hit[44] & (|(RS_ENCODE_PERMIT[44] & ~reg_be))) |
               (addr_hit[45] & (|(RS_ENCODE_PERMIT[45] & ~reg_be))) |
               (addr_hit[46] & (|(RS_ENCODE_PERMIT[46] & ~reg_be))) |
               (addr_hit[47] & (|(RS_ENCODE_PERMIT[47] & ~reg_be))) |
               (addr_hit[48] & (|(RS_ENCODE_PERMIT[48] & ~reg_be))) |
               (addr_hit[49] & (|(RS_ENCODE_PERMIT[49] & ~reg_be))) |
               (addr_hit[50] & (|(RS_ENCODE_PERMIT[50] & ~reg_be))) |
               (addr_hit[51] & (|(RS_ENCODE_PERMIT[51] & ~reg_be))) |
               (addr_hit[52] & (|(RS_ENCODE_PERMIT[52] & ~reg_be))) |
               (addr_hit[53] & (|(RS_ENCODE_PERMIT[53] & ~reg_be))) |
               (addr_hit[54] & (|(RS_ENCODE_PERMIT[54] & ~reg_be))) |
               (addr_hit[55] & (|(RS_ENCODE_PERMIT[55] & ~reg_be))) |
               (addr_hit[56] & (|(RS_ENCODE_PERMIT[56] & ~reg_be))) |
               (addr_hit[57] & (|(RS_ENCODE_PERMIT[57] & ~reg_be))) |
               (addr_hit[58] & (|(RS_ENCODE_PERMIT[58] & ~reg_be))) |
               (addr_hit[59] & (|(RS_ENCODE_PERMIT[59] & ~reg_be))) |
               (addr_hit[60] & (|(RS_ENCODE_PERMIT[60] & ~reg_be))) |
               (addr_hit[61] & (|(RS_ENCODE_PERMIT[61] & ~reg_be))) |
               (addr_hit[62] & (|(RS_ENCODE_PERMIT[62] & ~reg_be))) |
               (addr_hit[63] & (|(RS_ENCODE_PERMIT[63] & ~reg_be))) |
               (addr_hit[64] & (|(RS_ENCODE_PERMIT[64] & ~reg_be))) |
               (addr_hit[65] & (|(RS_ENCODE_PERMIT[65] & ~reg_be))) |
               (addr_hit[66] & (|(RS_ENCODE_PERMIT[66] & ~reg_be))) |
               (addr_hit[67] & (|(RS_ENCODE_PERMIT[67] & ~reg_be))) |
               (addr_hit[68] & (|(RS_ENCODE_PERMIT[68] & ~reg_be))) |
               (addr_hit[69] & (|(RS_ENCODE_PERMIT[69] & ~reg_be))) |
               (addr_hit[70] & (|(RS_ENCODE_PERMIT[70] & ~reg_be))) |
               (addr_hit[71] & (|(RS_ENCODE_PERMIT[71] & ~reg_be))) |
               (addr_hit[72] & (|(RS_ENCODE_PERMIT[72] & ~reg_be))) |
               (addr_hit[73] & (|(RS_ENCODE_PERMIT[73] & ~reg_be))) |
               (addr_hit[74] & (|(RS_ENCODE_PERMIT[74] & ~reg_be))) |
               (addr_hit[75] & (|(RS_ENCODE_PERMIT[75] & ~reg_be))) |
               (addr_hit[76] & (|(RS_ENCODE_PERMIT[76] & ~reg_be))) |
               (addr_hit[77] & (|(RS_ENCODE_PERMIT[77] & ~reg_be))) |
               (addr_hit[78] & (|(RS_ENCODE_PERMIT[78] & ~reg_be))) |
               (addr_hit[79] & (|(RS_ENCODE_PERMIT[79] & ~reg_be))) |
               (addr_hit[80] & (|(RS_ENCODE_PERMIT[80] & ~reg_be))) |
               (addr_hit[81] & (|(RS_ENCODE_PERMIT[81] & ~reg_be))) |
               (addr_hit[82] & (|(RS_ENCODE_PERMIT[82] & ~reg_be))) |
               (addr_hit[83] & (|(RS_ENCODE_PERMIT[83] & ~reg_be))) |
               (addr_hit[84] & (|(RS_ENCODE_PERMIT[84] & ~reg_be))) |
               (addr_hit[85] & (|(RS_ENCODE_PERMIT[85] & ~reg_be))) |
               (addr_hit[86] & (|(RS_ENCODE_PERMIT[86] & ~reg_be))) |
               (addr_hit[87] & (|(RS_ENCODE_PERMIT[87] & ~reg_be))) |
               (addr_hit[88] & (|(RS_ENCODE_PERMIT[88] & ~reg_be))) |
               (addr_hit[89] & (|(RS_ENCODE_PERMIT[89] & ~reg_be))) |
               (addr_hit[90] & (|(RS_ENCODE_PERMIT[90] & ~reg_be))) |
               (addr_hit[91] & (|(RS_ENCODE_PERMIT[91] & ~reg_be))) |
               (addr_hit[92] & (|(RS_ENCODE_PERMIT[92] & ~reg_be))) |
               (addr_hit[93] & (|(RS_ENCODE_PERMIT[93] & ~reg_be)))));
  end

  // Generate write-enables
  assign ctrl_signals_we = addr_hit[0] & reg_we & !reg_error;

  assign ctrl_signals_encode_en_wd = reg_wdata[0];

  assign ctrl_signals_clrn_wd = reg_wdata[1];
  assign data_in_0_we = addr_hit[2] & reg_we & !reg_error;

  assign data_in_0_wd = reg_wdata[31:0];
  assign data_in_1_we = addr_hit[3] & reg_we & !reg_error;

  assign data_in_1_wd = reg_wdata[31:0];
  assign data_in_2_we = addr_hit[4] & reg_we & !reg_error;

  assign data_in_2_wd = reg_wdata[31:0];
  assign data_in_3_we = addr_hit[5] & reg_we & !reg_error;

  assign data_in_3_wd = reg_wdata[31:0];
  assign data_in_4_we = addr_hit[6] & reg_we & !reg_error;

  assign data_in_4_wd = reg_wdata[31:0];
  assign data_in_5_we = addr_hit[7] & reg_we & !reg_error;

  assign data_in_5_wd = reg_wdata[31:0];
  assign data_in_6_we = addr_hit[8] & reg_we & !reg_error;

  assign data_in_6_wd = reg_wdata[31:0];
  assign data_in_7_we = addr_hit[9] & reg_we & !reg_error;

  assign data_in_7_wd = reg_wdata[31:0];
  assign data_in_8_we = addr_hit[10] & reg_we & !reg_error;

  assign data_in_8_wd = reg_wdata[31:0];
  assign data_in_9_we = addr_hit[11] & reg_we & !reg_error;

  assign data_in_9_wd = reg_wdata[31:0];
  assign data_in_10_we = addr_hit[12] & reg_we & !reg_error;

  assign data_in_10_wd = reg_wdata[31:0];
  assign data_in_11_we = addr_hit[13] & reg_we & !reg_error;

  assign data_in_11_wd = reg_wdata[31:0];
  assign data_in_12_we = addr_hit[14] & reg_we & !reg_error;

  assign data_in_12_wd = reg_wdata[31:0];
  assign data_in_13_we = addr_hit[15] & reg_we & !reg_error;

  assign data_in_13_wd = reg_wdata[31:0];
  assign data_in_14_we = addr_hit[16] & reg_we & !reg_error;

  assign data_in_14_wd = reg_wdata[31:0];
  assign data_in_15_we = addr_hit[17] & reg_we & !reg_error;

  assign data_in_15_wd = reg_wdata[31:0];
  assign data_in_16_we = addr_hit[18] & reg_we & !reg_error;

  assign data_in_16_wd = reg_wdata[31:0];
  assign data_in_17_we = addr_hit[19] & reg_we & !reg_error;

  assign data_in_17_wd = reg_wdata[31:0];
  assign data_in_18_we = addr_hit[20] & reg_we & !reg_error;

  assign data_in_18_wd = reg_wdata[31:0];
  assign data_in_19_we = addr_hit[21] & reg_we & !reg_error;

  assign data_in_19_wd = reg_wdata[31:0];
  assign data_in_20_we = addr_hit[22] & reg_we & !reg_error;

  assign data_in_20_wd = reg_wdata[31:0];
  assign data_in_21_we = addr_hit[23] & reg_we & !reg_error;

  assign data_in_21_wd = reg_wdata[31:0];
  assign data_in_22_we = addr_hit[24] & reg_we & !reg_error;

  assign data_in_22_wd = reg_wdata[31:0];
  assign data_in_23_we = addr_hit[25] & reg_we & !reg_error;

  assign data_in_23_wd = reg_wdata[31:0];
  assign data_in_24_we = addr_hit[26] & reg_we & !reg_error;

  assign data_in_24_wd = reg_wdata[31:0];
  assign data_in_25_we = addr_hit[27] & reg_we & !reg_error;

  assign data_in_25_wd = reg_wdata[31:0];
  assign data_in_26_we = addr_hit[28] & reg_we & !reg_error;

  assign data_in_26_wd = reg_wdata[31:0];
  assign data_in_27_we = addr_hit[29] & reg_we & !reg_error;

  assign data_in_27_wd = reg_wdata[31:0];
  assign data_in_28_we = addr_hit[30] & reg_we & !reg_error;

  assign data_in_28_wd = reg_wdata[31:0];
  assign data_in_29_we = addr_hit[31] & reg_we & !reg_error;

  assign data_in_29_wd = reg_wdata[31:0];
  assign data_in_30_we = addr_hit[32] & reg_we & !reg_error;

  assign data_in_30_wd = reg_wdata[31:0];
  assign data_in_31_we = addr_hit[33] & reg_we & !reg_error;

  assign data_in_31_wd = reg_wdata[31:0];
  assign data_in_32_we = addr_hit[34] & reg_we & !reg_error;

  assign data_in_32_wd = reg_wdata[31:0];
  assign data_in_33_we = addr_hit[35] & reg_we & !reg_error;

  assign data_in_33_wd = reg_wdata[31:0];
  assign data_in_34_we = addr_hit[36] & reg_we & !reg_error;

  assign data_in_34_wd = reg_wdata[31:0];
  assign data_in_35_we = addr_hit[37] & reg_we & !reg_error;

  assign data_in_35_wd = reg_wdata[31:0];
  assign data_in_36_we = addr_hit[38] & reg_we & !reg_error;

  assign data_in_36_wd = reg_wdata[31:0];
  assign data_in_37_we = addr_hit[39] & reg_we & !reg_error;

  assign data_in_37_wd = reg_wdata[31:0];
  assign data_in_38_we = addr_hit[40] & reg_we & !reg_error;

  assign data_in_38_wd = reg_wdata[31:0];
  assign data_in_39_we = addr_hit[41] & reg_we & !reg_error;

  assign data_in_39_wd = reg_wdata[31:0];
  assign data_in_40_we = addr_hit[42] & reg_we & !reg_error;

  assign data_in_40_wd = reg_wdata[31:0];
  assign data_in_41_we = addr_hit[43] & reg_we & !reg_error;

  assign data_in_41_wd = reg_wdata[31:0];

  // Assign write-enables to checker logic vector.
  always_comb begin
    reg_we_check = '0;
    reg_we_check[0] = ctrl_signals_we;
    reg_we_check[1] = 1'b0;
    reg_we_check[2] = data_in_0_we;
    reg_we_check[3] = data_in_1_we;
    reg_we_check[4] = data_in_2_we;
    reg_we_check[5] = data_in_3_we;
    reg_we_check[6] = data_in_4_we;
    reg_we_check[7] = data_in_5_we;
    reg_we_check[8] = data_in_6_we;
    reg_we_check[9] = data_in_7_we;
    reg_we_check[10] = data_in_8_we;
    reg_we_check[11] = data_in_9_we;
    reg_we_check[12] = data_in_10_we;
    reg_we_check[13] = data_in_11_we;
    reg_we_check[14] = data_in_12_we;
    reg_we_check[15] = data_in_13_we;
    reg_we_check[16] = data_in_14_we;
    reg_we_check[17] = data_in_15_we;
    reg_we_check[18] = data_in_16_we;
    reg_we_check[19] = data_in_17_we;
    reg_we_check[20] = data_in_18_we;
    reg_we_check[21] = data_in_19_we;
    reg_we_check[22] = data_in_20_we;
    reg_we_check[23] = data_in_21_we;
    reg_we_check[24] = data_in_22_we;
    reg_we_check[25] = data_in_23_we;
    reg_we_check[26] = data_in_24_we;
    reg_we_check[27] = data_in_25_we;
    reg_we_check[28] = data_in_26_we;
    reg_we_check[29] = data_in_27_we;
    reg_we_check[30] = data_in_28_we;
    reg_we_check[31] = data_in_29_we;
    reg_we_check[32] = data_in_30_we;
    reg_we_check[33] = data_in_31_we;
    reg_we_check[34] = data_in_32_we;
    reg_we_check[35] = data_in_33_we;
    reg_we_check[36] = data_in_34_we;
    reg_we_check[37] = data_in_35_we;
    reg_we_check[38] = data_in_36_we;
    reg_we_check[39] = data_in_37_we;
    reg_we_check[40] = data_in_38_we;
    reg_we_check[41] = data_in_39_we;
    reg_we_check[42] = data_in_40_we;
    reg_we_check[43] = data_in_41_we;
    reg_we_check[44] = 1'b0;
    reg_we_check[45] = 1'b0;
    reg_we_check[46] = 1'b0;
    reg_we_check[47] = 1'b0;
    reg_we_check[48] = 1'b0;
    reg_we_check[49] = 1'b0;
    reg_we_check[50] = 1'b0;
    reg_we_check[51] = 1'b0;
    reg_we_check[52] = 1'b0;
    reg_we_check[53] = 1'b0;
    reg_we_check[54] = 1'b0;
    reg_we_check[55] = 1'b0;
    reg_we_check[56] = 1'b0;
    reg_we_check[57] = 1'b0;
    reg_we_check[58] = 1'b0;
    reg_we_check[59] = 1'b0;
    reg_we_check[60] = 1'b0;
    reg_we_check[61] = 1'b0;
    reg_we_check[62] = 1'b0;
    reg_we_check[63] = 1'b0;
    reg_we_check[64] = 1'b0;
    reg_we_check[65] = 1'b0;
    reg_we_check[66] = 1'b0;
    reg_we_check[67] = 1'b0;
    reg_we_check[68] = 1'b0;
    reg_we_check[69] = 1'b0;
    reg_we_check[70] = 1'b0;
    reg_we_check[71] = 1'b0;
    reg_we_check[72] = 1'b0;
    reg_we_check[73] = 1'b0;
    reg_we_check[74] = 1'b0;
    reg_we_check[75] = 1'b0;
    reg_we_check[76] = 1'b0;
    reg_we_check[77] = 1'b0;
    reg_we_check[78] = 1'b0;
    reg_we_check[79] = 1'b0;
    reg_we_check[80] = 1'b0;
    reg_we_check[81] = 1'b0;
    reg_we_check[82] = 1'b0;
    reg_we_check[83] = 1'b0;
    reg_we_check[84] = 1'b0;
    reg_we_check[85] = 1'b0;
    reg_we_check[86] = 1'b0;
    reg_we_check[87] = 1'b0;
    reg_we_check[88] = 1'b0;
    reg_we_check[89] = 1'b0;
    reg_we_check[90] = 1'b0;
    reg_we_check[91] = 1'b0;
    reg_we_check[92] = 1'b0;
    reg_we_check[93] = 1'b0;
  end

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[0] = ctrl_signals_encode_en_qs;
        reg_rdata_next[1] = ctrl_signals_clrn_qs;
      end

      addr_hit[1]: begin
        reg_rdata_next[0] = state_signals_valid_bit_qs;
        reg_rdata_next[1] = state_signals_ready_bit_qs;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = data_in_0_qs;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = data_in_1_qs;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = data_in_2_qs;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = data_in_3_qs;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = data_in_4_qs;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = data_in_5_qs;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = data_in_6_qs;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = data_in_7_qs;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = data_in_8_qs;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = data_in_9_qs;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = data_in_10_qs;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = data_in_11_qs;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = data_in_12_qs;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = data_in_13_qs;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = data_in_14_qs;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = data_in_15_qs;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = data_in_16_qs;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = data_in_17_qs;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = data_in_18_qs;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = data_in_19_qs;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = data_in_20_qs;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = data_in_21_qs;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = data_in_22_qs;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = data_in_23_qs;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = data_in_24_qs;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = data_in_25_qs;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = data_in_26_qs;
      end

      addr_hit[29]: begin
        reg_rdata_next[31:0] = data_in_27_qs;
      end

      addr_hit[30]: begin
        reg_rdata_next[31:0] = data_in_28_qs;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = data_in_29_qs;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = data_in_30_qs;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = data_in_31_qs;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = data_in_32_qs;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = data_in_33_qs;
      end

      addr_hit[36]: begin
        reg_rdata_next[31:0] = data_in_34_qs;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = data_in_35_qs;
      end

      addr_hit[38]: begin
        reg_rdata_next[31:0] = data_in_36_qs;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = data_in_37_qs;
      end

      addr_hit[40]: begin
        reg_rdata_next[31:0] = data_in_38_qs;
      end

      addr_hit[41]: begin
        reg_rdata_next[31:0] = data_in_39_qs;
      end

      addr_hit[42]: begin
        reg_rdata_next[31:0] = data_in_40_qs;
      end

      addr_hit[43]: begin
        reg_rdata_next[31:0] = data_in_41_qs;
      end

      addr_hit[44]: begin
        reg_rdata_next[31:0] = encoded_data_out_0_qs;
      end

      addr_hit[45]: begin
        reg_rdata_next[31:0] = encoded_data_out_1_qs;
      end

      addr_hit[46]: begin
        reg_rdata_next[31:0] = encoded_data_out_2_qs;
      end

      addr_hit[47]: begin
        reg_rdata_next[31:0] = encoded_data_out_3_qs;
      end

      addr_hit[48]: begin
        reg_rdata_next[31:0] = encoded_data_out_4_qs;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = encoded_data_out_5_qs;
      end

      addr_hit[50]: begin
        reg_rdata_next[31:0] = encoded_data_out_6_qs;
      end

      addr_hit[51]: begin
        reg_rdata_next[31:0] = encoded_data_out_7_qs;
      end

      addr_hit[52]: begin
        reg_rdata_next[31:0] = encoded_data_out_8_qs;
      end

      addr_hit[53]: begin
        reg_rdata_next[31:0] = encoded_data_out_9_qs;
      end

      addr_hit[54]: begin
        reg_rdata_next[31:0] = encoded_data_out_10_qs;
      end

      addr_hit[55]: begin
        reg_rdata_next[31:0] = encoded_data_out_11_qs;
      end

      addr_hit[56]: begin
        reg_rdata_next[31:0] = encoded_data_out_12_qs;
      end

      addr_hit[57]: begin
        reg_rdata_next[31:0] = encoded_data_out_13_qs;
      end

      addr_hit[58]: begin
        reg_rdata_next[31:0] = encoded_data_out_14_qs;
      end

      addr_hit[59]: begin
        reg_rdata_next[31:0] = encoded_data_out_15_qs;
      end

      addr_hit[60]: begin
        reg_rdata_next[31:0] = encoded_data_out_16_qs;
      end

      addr_hit[61]: begin
        reg_rdata_next[31:0] = encoded_data_out_17_qs;
      end

      addr_hit[62]: begin
        reg_rdata_next[31:0] = encoded_data_out_18_qs;
      end

      addr_hit[63]: begin
        reg_rdata_next[31:0] = encoded_data_out_19_qs;
      end

      addr_hit[64]: begin
        reg_rdata_next[31:0] = encoded_data_out_20_qs;
      end

      addr_hit[65]: begin
        reg_rdata_next[31:0] = encoded_data_out_21_qs;
      end

      addr_hit[66]: begin
        reg_rdata_next[31:0] = encoded_data_out_22_qs;
      end

      addr_hit[67]: begin
        reg_rdata_next[31:0] = encoded_data_out_23_qs;
      end

      addr_hit[68]: begin
        reg_rdata_next[31:0] = encoded_data_out_24_qs;
      end

      addr_hit[69]: begin
        reg_rdata_next[31:0] = encoded_data_out_25_qs;
      end

      addr_hit[70]: begin
        reg_rdata_next[31:0] = encoded_data_out_26_qs;
      end

      addr_hit[71]: begin
        reg_rdata_next[31:0] = encoded_data_out_27_qs;
      end

      addr_hit[72]: begin
        reg_rdata_next[31:0] = encoded_data_out_28_qs;
      end

      addr_hit[73]: begin
        reg_rdata_next[31:0] = encoded_data_out_29_qs;
      end

      addr_hit[74]: begin
        reg_rdata_next[31:0] = encoded_data_out_30_qs;
      end

      addr_hit[75]: begin
        reg_rdata_next[31:0] = encoded_data_out_31_qs;
      end

      addr_hit[76]: begin
        reg_rdata_next[31:0] = encoded_data_out_32_qs;
      end

      addr_hit[77]: begin
        reg_rdata_next[31:0] = encoded_data_out_33_qs;
      end

      addr_hit[78]: begin
        reg_rdata_next[31:0] = encoded_data_out_34_qs;
      end

      addr_hit[79]: begin
        reg_rdata_next[31:0] = encoded_data_out_35_qs;
      end

      addr_hit[80]: begin
        reg_rdata_next[31:0] = encoded_data_out_36_qs;
      end

      addr_hit[81]: begin
        reg_rdata_next[31:0] = encoded_data_out_37_qs;
      end

      addr_hit[82]: begin
        reg_rdata_next[31:0] = encoded_data_out_38_qs;
      end

      addr_hit[83]: begin
        reg_rdata_next[31:0] = encoded_data_out_39_qs;
      end

      addr_hit[84]: begin
        reg_rdata_next[31:0] = encoded_data_out_40_qs;
      end

      addr_hit[85]: begin
        reg_rdata_next[31:0] = encoded_data_out_41_qs;
      end

      addr_hit[86]: begin
        reg_rdata_next[31:0] = encoded_data_out_42_qs;
      end

      addr_hit[87]: begin
        reg_rdata_next[31:0] = encoded_data_out_43_qs;
      end

      addr_hit[88]: begin
        reg_rdata_next[31:0] = encoded_data_out_44_qs;
      end

      addr_hit[89]: begin
        reg_rdata_next[31:0] = encoded_data_out_45_qs;
      end

      addr_hit[90]: begin
        reg_rdata_next[31:0] = encoded_data_out_46_qs;
      end

      addr_hit[91]: begin
        reg_rdata_next[31:0] = encoded_data_out_47_qs;
      end

      addr_hit[92]: begin
        reg_rdata_next[31:0] = encoded_data_out_48_qs;
      end

      addr_hit[93]: begin
        reg_rdata_next[31:0] = encoded_data_out_49_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // shadow busy
  logic shadow_busy;
  assign shadow_busy = 1'b0;

  // register busy
  assign reg_busy = shadow_busy;

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT_PULSE(wePulse, reg_we, clk_i, !rst_ni)
  `ASSERT_PULSE(rePulse, reg_re, clk_i, !rst_ni)

  `ASSERT(reAfterRv, $rose(reg_re || reg_we) |=> tl_o_pre.d_valid, clk_i, !rst_ni)

  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit), clk_i, !rst_ni)

  // this is formulated as an assumption such that the FPV testbenches do disprove this
  // property by mistake
  //`ASSUME(reqParity, tl_reg_h2d.a_valid |-> tl_reg_h2d.a_user.chk_en == tlul_pkg::CheckDis)

endmodule


`include "prim_assert.sv"

module rs_encode
  import rs_encode_reg_pkg::*;
(
  input  logic                                      clk_i,
  input  logic                                      rst_ni,
  input  logic                                      scan_mode,
  // Bus interface
  input  tlul_pkg::tl_h2d_t                         tl_i,
  output tlul_pkg::tl_d2h_t                         tl_o
);

  rs_encode_reg2hw_t               reg2hw;
  rs_encode_hw2reg_t               hw2reg;
  //wire                       ready_out;

  rs_encode_reg_top  u_rs_encode_reg_top (
    .clk_i                             ( clk_i           ),
    .rst_ni                            ( rst_ni          ),
    .tl_i                              ( tl_i            ),
    .hw2reg                            ( hw2reg          ),
    .devmode_i                         ( 1'b1            ),

    .tl_o                              ( tl_o            ),
    .reg2hw                            ( reg2hw          ),
    .intg_err_o                        (                 )
);

assign hw2reg.ctrl_signals.clrn.de = 1'd0;
assign hw2reg.ctrl_signals.encode_en.de = 1'd0;
always_comb begin
  for (int i = 0; i < 42; i++) begin
    hw2reg.data_in[i].de = 1'd0;
  end
end

rs_encode_wrapper  u_rs_encode_wrapper (
    .clk                     ( clk_i                         ),
    .rst_n                   ( rst_ni                        ),
    .clrn                    ( reg2hw.ctrl_signals.clrn.q ),
    .scan_mode                (scan_mode),
    .encode_en               ( reg2hw.ctrl_signals.encode_en.q ),
    .datain                  ( {reg2hw.data_in[41].q,reg2hw.data_in[40].q,reg2hw.data_in[39].q,reg2hw.data_in[38].q,reg2hw.data_in[37].q,reg2hw.data_in[36].q,reg2hw.data_in[35].q,reg2hw.data_in[34].q,reg2hw.data_in[33].q,reg2hw.data_in[32].q,reg2hw.data_in[31].q,reg2hw.data_in[30].q,reg2hw.data_in[29].q,reg2hw.data_in[28].q,reg2hw.data_in[27].q,reg2hw.data_in[26].q,reg2hw.data_in[25].q,reg2hw.data_in[24].q,reg2hw.data_in[23].q,reg2hw.data_in[22].q,reg2hw.data_in[21].q,reg2hw.data_in[20].q,reg2hw.data_in[19].q,reg2hw.data_in[18].q,reg2hw.data_in[17].q,reg2hw.data_in[16].q,reg2hw.data_in[15].q,reg2hw.data_in[14].q,reg2hw.data_in[13].q,reg2hw.data_in[12].q,reg2hw.data_in[11].q,reg2hw.data_in[10].q,reg2hw.data_in[9].q,reg2hw.data_in[8].q,reg2hw.data_in[7].q,reg2hw.data_in[6].q,reg2hw.data_in[5].q,reg2hw.data_in[4].q,reg2hw.data_in[3].q,reg2hw.data_in[2].q,reg2hw.data_in[1].q,reg2hw.data_in[0].q}),

    .encoded_data            ( {hw2reg.encoded_data_out[49].d,hw2reg.encoded_data_out[48].d,hw2reg.encoded_data_out[47].d,hw2reg.encoded_data_out[46].d,hw2reg.encoded_data_out[45].d,hw2reg.encoded_data_out[44].d,hw2reg.encoded_data_out[43].d,hw2reg.encoded_data_out[42].d,hw2reg.encoded_data_out[41].d,hw2reg.encoded_data_out[40].d,hw2reg.encoded_data_out[39].d,hw2reg.encoded_data_out[38].d,hw2reg.encoded_data_out[37].d,hw2reg.encoded_data_out[36].d,hw2reg.encoded_data_out[35].d,hw2reg.encoded_data_out[34].d,hw2reg.encoded_data_out[33].d,hw2reg.encoded_data_out[32].d,hw2reg.encoded_data_out[31].d,hw2reg.encoded_data_out[30].d,hw2reg.encoded_data_out[29].d,hw2reg.encoded_data_out[28].d,hw2reg.encoded_data_out[27].d,hw2reg.encoded_data_out[26].d,hw2reg.encoded_data_out[25].d,hw2reg.encoded_data_out[24].d,hw2reg.encoded_data_out[23].d,hw2reg.encoded_data_out[22].d,hw2reg.encoded_data_out[21].d,hw2reg.encoded_data_out[20].d,hw2reg.encoded_data_out[19].d,hw2reg.encoded_data_out[18].d,hw2reg.encoded_data_out[17].d,hw2reg.encoded_data_out[16].d,hw2reg.encoded_data_out[15].d,hw2reg.encoded_data_out[14].d,hw2reg.encoded_data_out[13].d,hw2reg.encoded_data_out[12].d,hw2reg.encoded_data_out[11].d,hw2reg.encoded_data_out[10].d,hw2reg.encoded_data_out[9].d,hw2reg.encoded_data_out[8].d,hw2reg.encoded_data_out[7].d,hw2reg.encoded_data_out[6].d,hw2reg.encoded_data_out[5].d,hw2reg.encoded_data_out[4].d,hw2reg.encoded_data_out[3].d,hw2reg.encoded_data_out[2].d,hw2reg.encoded_data_out[1].d,hw2reg.encoded_data_out[0].d} ),
    .valid                   ( hw2reg.state_signals.valid_bit.d ),
    .ready                   ( hw2reg.state_signals.ready_bit.d ),
    .ready_re                ( hw2reg.state_signals.ready_bit.de ),
    .valid_re                ( hw2reg.state_signals.valid_bit.de ),
    .encoded_data_re         ( {hw2reg.encoded_data_out[49].de,hw2reg.encoded_data_out[48].de,hw2reg.encoded_data_out[47].de,hw2reg.encoded_data_out[46].de,hw2reg.encoded_data_out[45].de,hw2reg.encoded_data_out[44].de,hw2reg.encoded_data_out[43].de,hw2reg.encoded_data_out[42].de,hw2reg.encoded_data_out[41].de,hw2reg.encoded_data_out[40].de,hw2reg.encoded_data_out[39].de,hw2reg.encoded_data_out[38].de,hw2reg.encoded_data_out[37].de,hw2reg.encoded_data_out[36].de,hw2reg.encoded_data_out[35].de,hw2reg.encoded_data_out[34].de,hw2reg.encoded_data_out[33].de,hw2reg.encoded_data_out[32].de,hw2reg.encoded_data_out[31].de,hw2reg.encoded_data_out[30].de,hw2reg.encoded_data_out[29].de,hw2reg.encoded_data_out[28].de,hw2reg.encoded_data_out[27].de,hw2reg.encoded_data_out[26].de,hw2reg.encoded_data_out[25].de,hw2reg.encoded_data_out[24].de,hw2reg.encoded_data_out[23].de,hw2reg.encoded_data_out[22].de,hw2reg.encoded_data_out[21].de,hw2reg.encoded_data_out[20].de,hw2reg.encoded_data_out[19].de,hw2reg.encoded_data_out[18].de,hw2reg.encoded_data_out[17].de,hw2reg.encoded_data_out[16].de,hw2reg.encoded_data_out[15].de,hw2reg.encoded_data_out[14].de,hw2reg.encoded_data_out[13].de,hw2reg.encoded_data_out[12].de,hw2reg.encoded_data_out[11].de,hw2reg.encoded_data_out[10].de,hw2reg.encoded_data_out[9].de,hw2reg.encoded_data_out[8].de,hw2reg.encoded_data_out[7].de,hw2reg.encoded_data_out[6].de,hw2reg.encoded_data_out[5].de,hw2reg.encoded_data_out[4].de,hw2reg.encoded_data_out[3].de,hw2reg.encoded_data_out[2].de,hw2reg.encoded_data_out[1].de,hw2reg.encoded_data_out[0].de} )
);

endmodule



