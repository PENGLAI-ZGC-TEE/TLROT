// -------------------------------------------------------------------------
//The inverse lookup table for Galois field
//Copyright (C) Tue Apr  2 17:07:28 2002
//by Ming-Han Lei(hendrik@humanistic.org)
//
//This program is free software; you can redistribute it and/or
//modify it under the terms of the GNU Lesser General Public License
//as published by the Free Software Foundation; either version 2
//of the License, or (at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU Lesser General Public License for more details.
//
//You should have received a copy of the GNU Lesser General Public License
//along with this program; if not, write to the Free Software
//Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
// --------------------------------------------------------------------------

module inverse(y, x);
	input [7:0] x;
	output [7:0] y;
	reg [7:0] y;

	always @ (x)
	case (x) // synopsys full_case parallel_case
		1: y = 1; // 0 -> 255
		2: y = 195; // 1 -> 254
		4: y = 162; // 2 -> 253
		8: y = 81; // 3 -> 252
		16: y = 235; // 4 -> 251
		32: y = 182; // 5 -> 250
		64: y = 91; // 6 -> 249
		128: y = 238; // 7 -> 248
		135: y = 119; // 8 -> 247
		137: y = 248; // 9 -> 246
		149: y = 124; // 10 -> 245
		173: y = 62; // 11 -> 244
		221: y = 31; // 12 -> 243
		61: y = 204; // 13 -> 242
		122: y = 102; // 14 -> 241
		244: y = 51; // 15 -> 240
		111: y = 218; // 16 -> 239
		222: y = 109; // 17 -> 238
		59: y = 245; // 18 -> 237
		118: y = 185; // 19 -> 236
		236: y = 159; // 20 -> 235
		95: y = 140; // 21 -> 234
		190: y = 70; // 22 -> 233
		251: y = 35; // 23 -> 232
		113: y = 210; // 24 -> 231
		226: y = 105; // 25 -> 230
		67: y = 247; // 26 -> 229
		134: y = 184; // 27 -> 228
		139: y = 92; // 28 -> 227
		145: y = 46; // 29 -> 226
		165: y = 23; // 30 -> 225
		205: y = 200; // 31 -> 224
		29: y = 100; // 32 -> 223
		58: y = 50; // 33 -> 222
		116: y = 25; // 34 -> 221
		232: y = 207; // 35 -> 220
		87: y = 164; // 36 -> 219
		174: y = 82; // 37 -> 218
		219: y = 41; // 38 -> 217
		49: y = 215; // 39 -> 216
		98: y = 168; // 40 -> 215
		196: y = 84; // 41 -> 214
		15: y = 42; // 42 -> 213
		30: y = 21; // 43 -> 212
		60: y = 201; // 44 -> 211
		120: y = 167; // 45 -> 210
		240: y = 144; // 46 -> 209
		103: y = 72; // 47 -> 208
		206: y = 36; // 48 -> 207
		27: y = 18; // 49 -> 206
		54: y = 9; // 50 -> 205
		108: y = 199; // 51 -> 204
		216: y = 160; // 52 -> 203
		55: y = 80; // 53 -> 202
		110: y = 40; // 54 -> 201
		220: y = 20; // 55 -> 200
		63: y = 10; // 56 -> 199
		126: y = 5; // 57 -> 198
		252: y = 193; // 58 -> 197
		127: y = 163; // 59 -> 196
		254: y = 146; // 60 -> 195
		123: y = 73; // 61 -> 194
		246: y = 231; // 62 -> 193
		107: y = 176; // 63 -> 192
		214: y = 88; // 64 -> 191
		43: y = 44; // 65 -> 190
		86: y = 22; // 66 -> 189
		172: y = 11; // 67 -> 188
		223: y = 198; // 68 -> 187
		57: y = 99; // 69 -> 186
		114: y = 242; // 70 -> 185
		228: y = 121; // 71 -> 184
		79: y = 255; // 72 -> 183
		158: y = 188; // 73 -> 182
		187: y = 94; // 74 -> 181
		241: y = 47; // 75 -> 180
		101: y = 212; // 76 -> 179
		202: y = 106; // 77 -> 178
		19: y = 53; // 78 -> 177
		38: y = 217; // 79 -> 176
		76: y = 175; // 80 -> 175
		152: y = 148; // 81 -> 174
		183: y = 74; // 82 -> 173
		233: y = 37; // 83 -> 172
		85: y = 209; // 84 -> 171
		170: y = 171; // 85 -> 170
		211: y = 150; // 86 -> 169
		33: y = 75; // 87 -> 168
		66: y = 230; // 88 -> 167
		132: y = 115; // 89 -> 166
		143: y = 250; // 90 -> 165
		153: y = 125; // 91 -> 164
		181: y = 253; // 92 -> 163
		237: y = 189; // 93 -> 162
		93: y = 157; // 94 -> 161
		186: y = 141; // 95 -> 160
		243: y = 133; // 96 -> 159
		97: y = 129; // 97 -> 158
		194: y = 131; // 98 -> 157
		3: y = 130; // 99 -> 156
		6: y = 65; // 100 -> 155
		12: y = 227; // 101 -> 154
		24: y = 178; // 102 -> 153
		48: y = 89; // 103 -> 152
		96: y = 239; // 104 -> 151
		192: y = 180; // 105 -> 150
		7: y = 90; // 106 -> 149
		14: y = 45; // 107 -> 148
		28: y = 213; // 108 -> 147
		56: y = 169; // 109 -> 146
		112: y = 151; // 110 -> 145
		224: y = 136; // 111 -> 144
		71: y = 68; // 112 -> 143
		142: y = 34; // 113 -> 142
		155: y = 17; // 114 -> 141
		177: y = 203; // 115 -> 140
		229: y = 166; // 116 -> 139
		77: y = 83; // 117 -> 138
		154: y = 234; // 118 -> 137
		179: y = 117; // 119 -> 136
		225: y = 249; // 120 -> 135
		69: y = 191; // 121 -> 134
		138: y = 156; // 122 -> 133
		147: y = 78; // 123 -> 132
		161: y = 39; // 124 -> 131
		197: y = 208; // 125 -> 130
		13: y = 104; // 126 -> 129
		26: y = 52; // 127 -> 128
		52: y = 26; // 128 -> 127
		104: y = 13; // 129 -> 126
		208: y = 197; // 130 -> 125
		39: y = 161; // 131 -> 124
		78: y = 147; // 132 -> 123
		156: y = 138; // 133 -> 122
		191: y = 69; // 134 -> 121
		249: y = 225; // 135 -> 120
		117: y = 179; // 136 -> 119
		234: y = 154; // 137 -> 118
		83: y = 77; // 138 -> 117
		166: y = 229; // 139 -> 116
		203: y = 177; // 140 -> 115
		17: y = 155; // 141 -> 114
		34: y = 142; // 142 -> 113
		68: y = 71; // 143 -> 112
		136: y = 224; // 144 -> 111
		151: y = 112; // 145 -> 110
		169: y = 56; // 146 -> 109
		213: y = 28; // 147 -> 108
		45: y = 14; // 148 -> 107
		90: y = 7; // 149 -> 106
		180: y = 192; // 150 -> 105
		239: y = 96; // 151 -> 104
		89: y = 48; // 152 -> 103
		178: y = 24; // 153 -> 102
		227: y = 12; // 154 -> 101
		65: y = 6; // 155 -> 100
		130: y = 3; // 156 -> 99
		131: y = 194; // 157 -> 98
		129: y = 97; // 158 -> 97
		133: y = 243; // 159 -> 96
		141: y = 186; // 160 -> 95
		157: y = 93; // 161 -> 94
		189: y = 237; // 162 -> 93
		253: y = 181; // 163 -> 92
		125: y = 153; // 164 -> 91
		250: y = 143; // 165 -> 90
		115: y = 132; // 166 -> 89
		230: y = 66; // 167 -> 88
		75: y = 33; // 168 -> 87
		150: y = 211; // 169 -> 86
		171: y = 170; // 170 -> 85
		209: y = 85; // 171 -> 84
		37: y = 233; // 172 -> 83
		74: y = 183; // 173 -> 82
		148: y = 152; // 174 -> 81
		175: y = 76; // 175 -> 80
		217: y = 38; // 176 -> 79
		53: y = 19; // 177 -> 78
		106: y = 202; // 178 -> 77
		212: y = 101; // 179 -> 76
		47: y = 241; // 180 -> 75
		94: y = 187; // 181 -> 74
		188: y = 158; // 182 -> 73
		255: y = 79; // 183 -> 72
		121: y = 228; // 184 -> 71
		242: y = 114; // 185 -> 70
		99: y = 57; // 186 -> 69
		198: y = 223; // 187 -> 68
		11: y = 172; // 188 -> 67
		22: y = 86; // 189 -> 66
		44: y = 43; // 190 -> 65
		88: y = 214; // 191 -> 64
		176: y = 107; // 192 -> 63
		231: y = 246; // 193 -> 62
		73: y = 123; // 194 -> 61
		146: y = 254; // 195 -> 60
		163: y = 127; // 196 -> 59
		193: y = 252; // 197 -> 58
		5: y = 126; // 198 -> 57
		10: y = 63; // 199 -> 56
		20: y = 220; // 200 -> 55
		40: y = 110; // 201 -> 54
		80: y = 55; // 202 -> 53
		160: y = 216; // 203 -> 52
		199: y = 108; // 204 -> 51
		9: y = 54; // 205 -> 50
		18: y = 27; // 206 -> 49
		36: y = 206; // 207 -> 48
		72: y = 103; // 208 -> 47
		144: y = 240; // 209 -> 46
		167: y = 120; // 210 -> 45
		201: y = 60; // 211 -> 44
		21: y = 30; // 212 -> 43
		42: y = 15; // 213 -> 42
		84: y = 196; // 214 -> 41
		168: y = 98; // 215 -> 40
		215: y = 49; // 216 -> 39
		41: y = 219; // 217 -> 38
		82: y = 174; // 218 -> 37
		164: y = 87; // 219 -> 36
		207: y = 232; // 220 -> 35
		25: y = 116; // 221 -> 34
		50: y = 58; // 222 -> 33
		100: y = 29; // 223 -> 32
		200: y = 205; // 224 -> 31
		23: y = 165; // 225 -> 30
		46: y = 145; // 226 -> 29
		92: y = 139; // 227 -> 28
		184: y = 134; // 228 -> 27
		247: y = 67; // 229 -> 26
		105: y = 226; // 230 -> 25
		210: y = 113; // 231 -> 24
		35: y = 251; // 232 -> 23
		70: y = 190; // 233 -> 22
		140: y = 95; // 234 -> 21
		159: y = 236; // 235 -> 20
		185: y = 118; // 236 -> 19
		245: y = 59; // 237 -> 18
		109: y = 222; // 238 -> 17
		218: y = 111; // 239 -> 16
		51: y = 244; // 240 -> 15
		102: y = 122; // 241 -> 14
		204: y = 61; // 242 -> 13
		31: y = 221; // 243 -> 12
		62: y = 173; // 244 -> 11
		124: y = 149; // 245 -> 10
		248: y = 137; // 246 -> 9
		119: y = 135; // 247 -> 8
		238: y = 128; // 248 -> 7
		91: y = 64; // 249 -> 6
		182: y = 32; // 250 -> 5
		235: y = 16; // 251 -> 4
		81: y = 8; // 252 -> 3
		162: y = 4; // 253 -> 2
		195: y = 2; // 254 -> 1
		default: y = 0;
	endcase
endmodule
